magic
tech sky130A
magscale 1 2
timestamp 1759434611
<< obsli1 >>
rect 1104 2159 68816 67473
<< obsm1 >>
rect 198 1368 69998 69284
<< metal2 >>
rect 3330 69200 3386 70000
rect 3606 69200 3662 70000
rect 3882 69200 3938 70000
rect 4158 69200 4214 70000
rect 4434 69200 4490 70000
rect 4710 69200 4766 70000
rect 4986 69200 5042 70000
rect 5262 69200 5318 70000
rect 5538 69200 5594 70000
rect 5814 69200 5870 70000
rect 6090 69200 6146 70000
rect 6366 69200 6422 70000
rect 6642 69200 6698 70000
rect 6918 69200 6974 70000
rect 7194 69200 7250 70000
rect 7470 69200 7526 70000
rect 7746 69200 7802 70000
rect 8022 69200 8078 70000
rect 8298 69200 8354 70000
rect 8574 69200 8630 70000
rect 8850 69200 8906 70000
rect 9126 69200 9182 70000
rect 9402 69200 9458 70000
rect 9678 69200 9734 70000
rect 9954 69200 10010 70000
rect 10230 69200 10286 70000
rect 10506 69200 10562 70000
rect 10782 69200 10838 70000
rect 11058 69200 11114 70000
rect 11334 69200 11390 70000
rect 11610 69200 11666 70000
rect 11886 69200 11942 70000
rect 12162 69200 12218 70000
rect 12438 69200 12494 70000
rect 12714 69200 12770 70000
rect 12990 69200 13046 70000
rect 13266 69200 13322 70000
rect 13542 69200 13598 70000
rect 13818 69200 13874 70000
rect 14094 69200 14150 70000
rect 14370 69200 14426 70000
rect 14646 69200 14702 70000
rect 14922 69200 14978 70000
rect 15198 69200 15254 70000
rect 15474 69200 15530 70000
rect 15750 69200 15806 70000
rect 16026 69200 16082 70000
rect 16302 69200 16358 70000
rect 16578 69200 16634 70000
rect 16854 69200 16910 70000
rect 17130 69200 17186 70000
rect 17406 69200 17462 70000
rect 17682 69200 17738 70000
rect 17958 69200 18014 70000
rect 18234 69200 18290 70000
rect 18510 69200 18566 70000
rect 18786 69200 18842 70000
rect 19062 69200 19118 70000
rect 19338 69200 19394 70000
rect 19614 69200 19670 70000
rect 19890 69200 19946 70000
rect 20166 69200 20222 70000
rect 20442 69200 20498 70000
rect 20718 69200 20774 70000
rect 20994 69200 21050 70000
rect 21270 69200 21326 70000
rect 21546 69200 21602 70000
rect 21822 69200 21878 70000
rect 22098 69200 22154 70000
rect 22374 69200 22430 70000
rect 22650 69200 22706 70000
rect 22926 69200 22982 70000
rect 23202 69200 23258 70000
rect 23478 69200 23534 70000
rect 23754 69200 23810 70000
rect 24030 69200 24086 70000
rect 24306 69200 24362 70000
rect 24582 69200 24638 70000
rect 24858 69200 24914 70000
rect 25134 69200 25190 70000
rect 25410 69200 25466 70000
rect 25686 69200 25742 70000
rect 25962 69200 26018 70000
rect 26238 69200 26294 70000
rect 26514 69200 26570 70000
rect 26790 69200 26846 70000
rect 27066 69200 27122 70000
rect 27342 69200 27398 70000
rect 27618 69200 27674 70000
rect 27894 69200 27950 70000
rect 28170 69200 28226 70000
rect 28446 69200 28502 70000
rect 28722 69200 28778 70000
rect 28998 69200 29054 70000
rect 29274 69200 29330 70000
rect 29550 69200 29606 70000
rect 29826 69200 29882 70000
rect 30102 69200 30158 70000
rect 30378 69200 30434 70000
rect 30654 69200 30710 70000
rect 30930 69200 30986 70000
rect 31206 69200 31262 70000
rect 31482 69200 31538 70000
rect 31758 69200 31814 70000
rect 32034 69200 32090 70000
rect 32310 69200 32366 70000
rect 32586 69200 32642 70000
rect 32862 69200 32918 70000
rect 33138 69200 33194 70000
rect 33414 69200 33470 70000
rect 33690 69200 33746 70000
rect 33966 69200 34022 70000
rect 34242 69200 34298 70000
rect 34518 69200 34574 70000
rect 34794 69200 34850 70000
rect 35070 69200 35126 70000
rect 35346 69200 35402 70000
rect 35622 69200 35678 70000
rect 35898 69200 35954 70000
rect 36174 69200 36230 70000
rect 36450 69200 36506 70000
rect 36726 69200 36782 70000
rect 37002 69200 37058 70000
rect 37278 69200 37334 70000
rect 37554 69200 37610 70000
rect 37830 69200 37886 70000
rect 38106 69200 38162 70000
rect 38382 69200 38438 70000
rect 38658 69200 38714 70000
rect 38934 69200 38990 70000
rect 39210 69200 39266 70000
rect 39486 69200 39542 70000
rect 39762 69200 39818 70000
rect 40038 69200 40094 70000
rect 40314 69200 40370 70000
rect 40590 69200 40646 70000
rect 40866 69200 40922 70000
rect 41142 69200 41198 70000
rect 41418 69200 41474 70000
rect 41694 69200 41750 70000
rect 41970 69200 42026 70000
rect 42246 69200 42302 70000
rect 42522 69200 42578 70000
rect 42798 69200 42854 70000
rect 43074 69200 43130 70000
rect 43350 69200 43406 70000
rect 43626 69200 43682 70000
rect 43902 69200 43958 70000
rect 44178 69200 44234 70000
rect 44454 69200 44510 70000
rect 44730 69200 44786 70000
rect 45006 69200 45062 70000
rect 45282 69200 45338 70000
rect 45558 69200 45614 70000
rect 45834 69200 45890 70000
rect 46110 69200 46166 70000
rect 46386 69200 46442 70000
rect 46662 69200 46718 70000
rect 46938 69200 46994 70000
rect 47214 69200 47270 70000
rect 47490 69200 47546 70000
rect 47766 69200 47822 70000
rect 48042 69200 48098 70000
rect 48318 69200 48374 70000
rect 48594 69200 48650 70000
rect 48870 69200 48926 70000
rect 49146 69200 49202 70000
rect 49422 69200 49478 70000
rect 49698 69200 49754 70000
rect 49974 69200 50030 70000
rect 50250 69200 50306 70000
rect 50526 69200 50582 70000
rect 50802 69200 50858 70000
rect 51078 69200 51134 70000
rect 51354 69200 51410 70000
rect 51630 69200 51686 70000
rect 51906 69200 51962 70000
rect 52182 69200 52238 70000
rect 52458 69200 52514 70000
rect 52734 69200 52790 70000
rect 53010 69200 53066 70000
rect 53286 69200 53342 70000
rect 53562 69200 53618 70000
rect 53838 69200 53894 70000
rect 54114 69200 54170 70000
rect 54390 69200 54446 70000
rect 54666 69200 54722 70000
rect 54942 69200 54998 70000
rect 55218 69200 55274 70000
rect 55494 69200 55550 70000
rect 55770 69200 55826 70000
rect 56046 69200 56102 70000
rect 56322 69200 56378 70000
rect 56598 69200 56654 70000
rect 56874 69200 56930 70000
rect 57150 69200 57206 70000
rect 57426 69200 57482 70000
rect 57702 69200 57758 70000
rect 57978 69200 58034 70000
rect 58254 69200 58310 70000
rect 58530 69200 58586 70000
rect 58806 69200 58862 70000
rect 59082 69200 59138 70000
rect 59358 69200 59414 70000
rect 59634 69200 59690 70000
rect 59910 69200 59966 70000
rect 60186 69200 60242 70000
rect 60462 69200 60518 70000
rect 60738 69200 60794 70000
rect 61014 69200 61070 70000
rect 61290 69200 61346 70000
rect 61566 69200 61622 70000
rect 61842 69200 61898 70000
rect 62118 69200 62174 70000
rect 62394 69200 62450 70000
rect 62670 69200 62726 70000
rect 62946 69200 63002 70000
rect 63222 69200 63278 70000
rect 63498 69200 63554 70000
rect 63774 69200 63830 70000
rect 64050 69200 64106 70000
rect 64326 69200 64382 70000
rect 64602 69200 64658 70000
rect 64878 69200 64934 70000
rect 65154 69200 65210 70000
rect 65430 69200 65486 70000
rect 65706 69200 65762 70000
rect 65982 69200 66038 70000
rect 66258 69200 66314 70000
rect 66534 69200 66590 70000
rect 3882 0 3938 800
rect 4342 0 4398 800
rect 4802 0 4858 800
rect 5262 0 5318 800
rect 5722 0 5778 800
rect 6182 0 6238 800
rect 6642 0 6698 800
rect 7102 0 7158 800
rect 7562 0 7618 800
rect 8022 0 8078 800
rect 8482 0 8538 800
rect 8942 0 8998 800
rect 9402 0 9458 800
rect 9862 0 9918 800
rect 10322 0 10378 800
rect 10782 0 10838 800
rect 11242 0 11298 800
rect 11702 0 11758 800
rect 12162 0 12218 800
rect 12622 0 12678 800
rect 13082 0 13138 800
rect 13542 0 13598 800
rect 14002 0 14058 800
rect 14462 0 14518 800
rect 14922 0 14978 800
rect 15382 0 15438 800
rect 15842 0 15898 800
rect 16302 0 16358 800
rect 16762 0 16818 800
rect 17222 0 17278 800
rect 17682 0 17738 800
rect 18142 0 18198 800
rect 18602 0 18658 800
rect 19062 0 19118 800
rect 19522 0 19578 800
rect 19982 0 20038 800
rect 20442 0 20498 800
rect 20902 0 20958 800
rect 21362 0 21418 800
rect 21822 0 21878 800
rect 22282 0 22338 800
rect 22742 0 22798 800
rect 23202 0 23258 800
rect 23662 0 23718 800
rect 24122 0 24178 800
rect 24582 0 24638 800
rect 25042 0 25098 800
rect 25502 0 25558 800
rect 25962 0 26018 800
rect 26422 0 26478 800
rect 26882 0 26938 800
rect 27342 0 27398 800
rect 27802 0 27858 800
rect 28262 0 28318 800
rect 28722 0 28778 800
rect 29182 0 29238 800
rect 29642 0 29698 800
rect 30102 0 30158 800
rect 30562 0 30618 800
rect 31022 0 31078 800
rect 31482 0 31538 800
rect 31942 0 31998 800
rect 32402 0 32458 800
rect 32862 0 32918 800
rect 33322 0 33378 800
rect 33782 0 33838 800
rect 34242 0 34298 800
rect 34702 0 34758 800
rect 35162 0 35218 800
rect 35622 0 35678 800
rect 36082 0 36138 800
rect 36542 0 36598 800
rect 37002 0 37058 800
rect 37462 0 37518 800
rect 37922 0 37978 800
rect 38382 0 38438 800
rect 38842 0 38898 800
rect 39302 0 39358 800
rect 39762 0 39818 800
rect 40222 0 40278 800
rect 40682 0 40738 800
rect 41142 0 41198 800
rect 41602 0 41658 800
rect 42062 0 42118 800
rect 42522 0 42578 800
rect 42982 0 43038 800
rect 43442 0 43498 800
rect 43902 0 43958 800
rect 44362 0 44418 800
rect 44822 0 44878 800
rect 45282 0 45338 800
rect 45742 0 45798 800
rect 46202 0 46258 800
rect 46662 0 46718 800
rect 47122 0 47178 800
rect 47582 0 47638 800
rect 48042 0 48098 800
rect 48502 0 48558 800
rect 48962 0 49018 800
rect 49422 0 49478 800
rect 49882 0 49938 800
rect 50342 0 50398 800
rect 50802 0 50858 800
rect 51262 0 51318 800
rect 51722 0 51778 800
rect 52182 0 52238 800
rect 52642 0 52698 800
rect 53102 0 53158 800
rect 53562 0 53618 800
rect 54022 0 54078 800
rect 54482 0 54538 800
rect 54942 0 54998 800
rect 55402 0 55458 800
rect 55862 0 55918 800
rect 56322 0 56378 800
rect 56782 0 56838 800
rect 57242 0 57298 800
rect 57702 0 57758 800
rect 58162 0 58218 800
rect 58622 0 58678 800
rect 59082 0 59138 800
rect 59542 0 59598 800
rect 60002 0 60058 800
rect 60462 0 60518 800
rect 60922 0 60978 800
rect 61382 0 61438 800
rect 61842 0 61898 800
rect 62302 0 62358 800
rect 62762 0 62818 800
rect 63222 0 63278 800
rect 63682 0 63738 800
rect 64142 0 64198 800
rect 64602 0 64658 800
rect 65062 0 65118 800
rect 65522 0 65578 800
rect 65982 0 66038 800
<< obsm2 >>
rect 204 69144 3274 69306
rect 3442 69144 3550 69306
rect 3718 69144 3826 69306
rect 3994 69144 4102 69306
rect 4270 69144 4378 69306
rect 4546 69144 4654 69306
rect 4822 69144 4930 69306
rect 5098 69144 5206 69306
rect 5374 69144 5482 69306
rect 5650 69144 5758 69306
rect 5926 69144 6034 69306
rect 6202 69144 6310 69306
rect 6478 69144 6586 69306
rect 6754 69144 6862 69306
rect 7030 69144 7138 69306
rect 7306 69144 7414 69306
rect 7582 69144 7690 69306
rect 7858 69144 7966 69306
rect 8134 69144 8242 69306
rect 8410 69144 8518 69306
rect 8686 69144 8794 69306
rect 8962 69144 9070 69306
rect 9238 69144 9346 69306
rect 9514 69144 9622 69306
rect 9790 69144 9898 69306
rect 10066 69144 10174 69306
rect 10342 69144 10450 69306
rect 10618 69144 10726 69306
rect 10894 69144 11002 69306
rect 11170 69144 11278 69306
rect 11446 69144 11554 69306
rect 11722 69144 11830 69306
rect 11998 69144 12106 69306
rect 12274 69144 12382 69306
rect 12550 69144 12658 69306
rect 12826 69144 12934 69306
rect 13102 69144 13210 69306
rect 13378 69144 13486 69306
rect 13654 69144 13762 69306
rect 13930 69144 14038 69306
rect 14206 69144 14314 69306
rect 14482 69144 14590 69306
rect 14758 69144 14866 69306
rect 15034 69144 15142 69306
rect 15310 69144 15418 69306
rect 15586 69144 15694 69306
rect 15862 69144 15970 69306
rect 16138 69144 16246 69306
rect 16414 69144 16522 69306
rect 16690 69144 16798 69306
rect 16966 69144 17074 69306
rect 17242 69144 17350 69306
rect 17518 69144 17626 69306
rect 17794 69144 17902 69306
rect 18070 69144 18178 69306
rect 18346 69144 18454 69306
rect 18622 69144 18730 69306
rect 18898 69144 19006 69306
rect 19174 69144 19282 69306
rect 19450 69144 19558 69306
rect 19726 69144 19834 69306
rect 20002 69144 20110 69306
rect 20278 69144 20386 69306
rect 20554 69144 20662 69306
rect 20830 69144 20938 69306
rect 21106 69144 21214 69306
rect 21382 69144 21490 69306
rect 21658 69144 21766 69306
rect 21934 69144 22042 69306
rect 22210 69144 22318 69306
rect 22486 69144 22594 69306
rect 22762 69144 22870 69306
rect 23038 69144 23146 69306
rect 23314 69144 23422 69306
rect 23590 69144 23698 69306
rect 23866 69144 23974 69306
rect 24142 69144 24250 69306
rect 24418 69144 24526 69306
rect 24694 69144 24802 69306
rect 24970 69144 25078 69306
rect 25246 69144 25354 69306
rect 25522 69144 25630 69306
rect 25798 69144 25906 69306
rect 26074 69144 26182 69306
rect 26350 69144 26458 69306
rect 26626 69144 26734 69306
rect 26902 69144 27010 69306
rect 27178 69144 27286 69306
rect 27454 69144 27562 69306
rect 27730 69144 27838 69306
rect 28006 69144 28114 69306
rect 28282 69144 28390 69306
rect 28558 69144 28666 69306
rect 28834 69144 28942 69306
rect 29110 69144 29218 69306
rect 29386 69144 29494 69306
rect 29662 69144 29770 69306
rect 29938 69144 30046 69306
rect 30214 69144 30322 69306
rect 30490 69144 30598 69306
rect 30766 69144 30874 69306
rect 31042 69144 31150 69306
rect 31318 69144 31426 69306
rect 31594 69144 31702 69306
rect 31870 69144 31978 69306
rect 32146 69144 32254 69306
rect 32422 69144 32530 69306
rect 32698 69144 32806 69306
rect 32974 69144 33082 69306
rect 33250 69144 33358 69306
rect 33526 69144 33634 69306
rect 33802 69144 33910 69306
rect 34078 69144 34186 69306
rect 34354 69144 34462 69306
rect 34630 69144 34738 69306
rect 34906 69144 35014 69306
rect 35182 69144 35290 69306
rect 35458 69144 35566 69306
rect 35734 69144 35842 69306
rect 36010 69144 36118 69306
rect 36286 69144 36394 69306
rect 36562 69144 36670 69306
rect 36838 69144 36946 69306
rect 37114 69144 37222 69306
rect 37390 69144 37498 69306
rect 37666 69144 37774 69306
rect 37942 69144 38050 69306
rect 38218 69144 38326 69306
rect 38494 69144 38602 69306
rect 38770 69144 38878 69306
rect 39046 69144 39154 69306
rect 39322 69144 39430 69306
rect 39598 69144 39706 69306
rect 39874 69144 39982 69306
rect 40150 69144 40258 69306
rect 40426 69144 40534 69306
rect 40702 69144 40810 69306
rect 40978 69144 41086 69306
rect 41254 69144 41362 69306
rect 41530 69144 41638 69306
rect 41806 69144 41914 69306
rect 42082 69144 42190 69306
rect 42358 69144 42466 69306
rect 42634 69144 42742 69306
rect 42910 69144 43018 69306
rect 43186 69144 43294 69306
rect 43462 69144 43570 69306
rect 43738 69144 43846 69306
rect 44014 69144 44122 69306
rect 44290 69144 44398 69306
rect 44566 69144 44674 69306
rect 44842 69144 44950 69306
rect 45118 69144 45226 69306
rect 45394 69144 45502 69306
rect 45670 69144 45778 69306
rect 45946 69144 46054 69306
rect 46222 69144 46330 69306
rect 46498 69144 46606 69306
rect 46774 69144 46882 69306
rect 47050 69144 47158 69306
rect 47326 69144 47434 69306
rect 47602 69144 47710 69306
rect 47878 69144 47986 69306
rect 48154 69144 48262 69306
rect 48430 69144 48538 69306
rect 48706 69144 48814 69306
rect 48982 69144 49090 69306
rect 49258 69144 49366 69306
rect 49534 69144 49642 69306
rect 49810 69144 49918 69306
rect 50086 69144 50194 69306
rect 50362 69144 50470 69306
rect 50638 69144 50746 69306
rect 50914 69144 51022 69306
rect 51190 69144 51298 69306
rect 51466 69144 51574 69306
rect 51742 69144 51850 69306
rect 52018 69144 52126 69306
rect 52294 69144 52402 69306
rect 52570 69144 52678 69306
rect 52846 69144 52954 69306
rect 53122 69144 53230 69306
rect 53398 69144 53506 69306
rect 53674 69144 53782 69306
rect 53950 69144 54058 69306
rect 54226 69144 54334 69306
rect 54502 69144 54610 69306
rect 54778 69144 54886 69306
rect 55054 69144 55162 69306
rect 55330 69144 55438 69306
rect 55606 69144 55714 69306
rect 55882 69144 55990 69306
rect 56158 69144 56266 69306
rect 56434 69144 56542 69306
rect 56710 69144 56818 69306
rect 56986 69144 57094 69306
rect 57262 69144 57370 69306
rect 57538 69144 57646 69306
rect 57814 69144 57922 69306
rect 58090 69144 58198 69306
rect 58366 69144 58474 69306
rect 58642 69144 58750 69306
rect 58918 69144 59026 69306
rect 59194 69144 59302 69306
rect 59470 69144 59578 69306
rect 59746 69144 59854 69306
rect 60022 69144 60130 69306
rect 60298 69144 60406 69306
rect 60574 69144 60682 69306
rect 60850 69144 60958 69306
rect 61126 69144 61234 69306
rect 61402 69144 61510 69306
rect 61678 69144 61786 69306
rect 61954 69144 62062 69306
rect 62230 69144 62338 69306
rect 62506 69144 62614 69306
rect 62782 69144 62890 69306
rect 63058 69144 63166 69306
rect 63334 69144 63442 69306
rect 63610 69144 63718 69306
rect 63886 69144 63994 69306
rect 64162 69144 64270 69306
rect 64438 69144 64546 69306
rect 64714 69144 64822 69306
rect 64990 69144 65098 69306
rect 65266 69144 65374 69306
rect 65542 69144 65650 69306
rect 65818 69144 65926 69306
rect 66094 69144 66202 69306
rect 66370 69144 66478 69306
rect 66646 69144 69992 69306
rect 204 856 69992 69144
rect 204 734 3826 856
rect 3994 734 4286 856
rect 4454 734 4746 856
rect 4914 734 5206 856
rect 5374 734 5666 856
rect 5834 734 6126 856
rect 6294 734 6586 856
rect 6754 734 7046 856
rect 7214 734 7506 856
rect 7674 734 7966 856
rect 8134 734 8426 856
rect 8594 734 8886 856
rect 9054 734 9346 856
rect 9514 734 9806 856
rect 9974 734 10266 856
rect 10434 734 10726 856
rect 10894 734 11186 856
rect 11354 734 11646 856
rect 11814 734 12106 856
rect 12274 734 12566 856
rect 12734 734 13026 856
rect 13194 734 13486 856
rect 13654 734 13946 856
rect 14114 734 14406 856
rect 14574 734 14866 856
rect 15034 734 15326 856
rect 15494 734 15786 856
rect 15954 734 16246 856
rect 16414 734 16706 856
rect 16874 734 17166 856
rect 17334 734 17626 856
rect 17794 734 18086 856
rect 18254 734 18546 856
rect 18714 734 19006 856
rect 19174 734 19466 856
rect 19634 734 19926 856
rect 20094 734 20386 856
rect 20554 734 20846 856
rect 21014 734 21306 856
rect 21474 734 21766 856
rect 21934 734 22226 856
rect 22394 734 22686 856
rect 22854 734 23146 856
rect 23314 734 23606 856
rect 23774 734 24066 856
rect 24234 734 24526 856
rect 24694 734 24986 856
rect 25154 734 25446 856
rect 25614 734 25906 856
rect 26074 734 26366 856
rect 26534 734 26826 856
rect 26994 734 27286 856
rect 27454 734 27746 856
rect 27914 734 28206 856
rect 28374 734 28666 856
rect 28834 734 29126 856
rect 29294 734 29586 856
rect 29754 734 30046 856
rect 30214 734 30506 856
rect 30674 734 30966 856
rect 31134 734 31426 856
rect 31594 734 31886 856
rect 32054 734 32346 856
rect 32514 734 32806 856
rect 32974 734 33266 856
rect 33434 734 33726 856
rect 33894 734 34186 856
rect 34354 734 34646 856
rect 34814 734 35106 856
rect 35274 734 35566 856
rect 35734 734 36026 856
rect 36194 734 36486 856
rect 36654 734 36946 856
rect 37114 734 37406 856
rect 37574 734 37866 856
rect 38034 734 38326 856
rect 38494 734 38786 856
rect 38954 734 39246 856
rect 39414 734 39706 856
rect 39874 734 40166 856
rect 40334 734 40626 856
rect 40794 734 41086 856
rect 41254 734 41546 856
rect 41714 734 42006 856
rect 42174 734 42466 856
rect 42634 734 42926 856
rect 43094 734 43386 856
rect 43554 734 43846 856
rect 44014 734 44306 856
rect 44474 734 44766 856
rect 44934 734 45226 856
rect 45394 734 45686 856
rect 45854 734 46146 856
rect 46314 734 46606 856
rect 46774 734 47066 856
rect 47234 734 47526 856
rect 47694 734 47986 856
rect 48154 734 48446 856
rect 48614 734 48906 856
rect 49074 734 49366 856
rect 49534 734 49826 856
rect 49994 734 50286 856
rect 50454 734 50746 856
rect 50914 734 51206 856
rect 51374 734 51666 856
rect 51834 734 52126 856
rect 52294 734 52586 856
rect 52754 734 53046 856
rect 53214 734 53506 856
rect 53674 734 53966 856
rect 54134 734 54426 856
rect 54594 734 54886 856
rect 55054 734 55346 856
rect 55514 734 55806 856
rect 55974 734 56266 856
rect 56434 734 56726 856
rect 56894 734 57186 856
rect 57354 734 57646 856
rect 57814 734 58106 856
rect 58274 734 58566 856
rect 58734 734 59026 856
rect 59194 734 59486 856
rect 59654 734 59946 856
rect 60114 734 60406 856
rect 60574 734 60866 856
rect 61034 734 61326 856
rect 61494 734 61786 856
rect 61954 734 62246 856
rect 62414 734 62706 856
rect 62874 734 63166 856
rect 63334 734 63626 856
rect 63794 734 64086 856
rect 64254 734 64546 856
rect 64714 734 65006 856
rect 65174 734 65466 856
rect 65634 734 65926 856
rect 66094 734 69992 856
<< metal3 >>
rect 0 65560 800 65680
rect 0 65288 800 65408
rect 0 65016 800 65136
rect 0 64744 800 64864
rect 0 64472 800 64592
rect 0 64200 800 64320
rect 0 63928 800 64048
rect 0 63656 800 63776
rect 0 63384 800 63504
rect 0 63112 800 63232
rect 0 62840 800 62960
rect 0 62568 800 62688
rect 0 62296 800 62416
rect 0 62024 800 62144
rect 0 61752 800 61872
rect 0 61480 800 61600
rect 0 61208 800 61328
rect 0 60936 800 61056
rect 0 60664 800 60784
rect 0 60392 800 60512
rect 0 60120 800 60240
rect 0 59848 800 59968
rect 0 59576 800 59696
rect 0 59304 800 59424
rect 0 59032 800 59152
rect 0 58760 800 58880
rect 0 58488 800 58608
rect 0 58216 800 58336
rect 0 57944 800 58064
rect 0 57672 800 57792
rect 0 57400 800 57520
rect 0 57128 800 57248
rect 0 56856 800 56976
rect 0 56584 800 56704
rect 0 56312 800 56432
rect 0 56040 800 56160
rect 0 55768 800 55888
rect 0 55496 800 55616
rect 0 55224 800 55344
rect 0 54952 800 55072
rect 0 54680 800 54800
rect 0 54408 800 54528
rect 0 54136 800 54256
rect 0 53864 800 53984
rect 0 53592 800 53712
rect 0 53320 800 53440
rect 0 53048 800 53168
rect 0 52776 800 52896
rect 0 52504 800 52624
rect 0 52232 800 52352
rect 0 51960 800 52080
rect 0 51688 800 51808
rect 0 51416 800 51536
rect 0 51144 800 51264
rect 0 50872 800 50992
rect 0 50600 800 50720
rect 0 50328 800 50448
rect 0 50056 800 50176
rect 0 49784 800 49904
rect 0 49512 800 49632
rect 0 49240 800 49360
rect 0 48968 800 49088
rect 0 48696 800 48816
rect 0 48424 800 48544
rect 0 48152 800 48272
rect 0 47880 800 48000
rect 0 47608 800 47728
rect 0 47336 800 47456
rect 0 47064 800 47184
rect 0 46792 800 46912
rect 0 46520 800 46640
rect 0 46248 800 46368
rect 0 45976 800 46096
rect 0 45704 800 45824
rect 0 45432 800 45552
rect 0 45160 800 45280
rect 0 44888 800 45008
rect 0 44616 800 44736
rect 0 44344 800 44464
rect 0 44072 800 44192
rect 0 43800 800 43920
rect 0 43528 800 43648
rect 0 43256 800 43376
rect 0 42984 800 43104
rect 0 42712 800 42832
rect 0 42440 800 42560
rect 0 42168 800 42288
rect 0 41896 800 42016
rect 0 41624 800 41744
rect 0 41352 800 41472
rect 0 41080 800 41200
rect 0 40808 800 40928
rect 0 40536 800 40656
rect 0 40264 800 40384
rect 0 39992 800 40112
rect 0 39720 800 39840
rect 0 39448 800 39568
rect 0 39176 800 39296
rect 0 38904 800 39024
rect 0 38632 800 38752
rect 0 38360 800 38480
rect 0 38088 800 38208
rect 0 37816 800 37936
rect 0 37544 800 37664
rect 0 37272 800 37392
rect 0 37000 800 37120
rect 0 36728 800 36848
rect 0 36456 800 36576
rect 0 36184 800 36304
rect 0 35912 800 36032
rect 0 35640 800 35760
rect 0 35368 800 35488
rect 0 35096 800 35216
rect 0 34824 800 34944
rect 0 34552 800 34672
rect 0 34280 800 34400
rect 0 34008 800 34128
rect 0 33736 800 33856
rect 0 33464 800 33584
rect 0 33192 800 33312
rect 0 32920 800 33040
rect 0 32648 800 32768
rect 0 32376 800 32496
rect 0 32104 800 32224
rect 0 31832 800 31952
rect 0 31560 800 31680
rect 0 31288 800 31408
rect 0 31016 800 31136
rect 0 30744 800 30864
rect 0 30472 800 30592
rect 0 30200 800 30320
rect 0 29928 800 30048
rect 0 29656 800 29776
rect 0 29384 800 29504
rect 0 29112 800 29232
rect 0 28840 800 28960
rect 0 28568 800 28688
rect 0 28296 800 28416
rect 0 28024 800 28144
rect 0 27752 800 27872
rect 0 27480 800 27600
rect 0 27208 800 27328
rect 0 26936 800 27056
rect 0 26664 800 26784
rect 0 26392 800 26512
rect 0 26120 800 26240
rect 0 25848 800 25968
rect 0 25576 800 25696
rect 0 25304 800 25424
rect 0 25032 800 25152
rect 0 24760 800 24880
rect 0 24488 800 24608
rect 0 24216 800 24336
rect 0 23944 800 24064
rect 0 23672 800 23792
rect 0 23400 800 23520
rect 0 23128 800 23248
rect 0 22856 800 22976
rect 0 22584 800 22704
rect 0 22312 800 22432
rect 0 22040 800 22160
rect 0 21768 800 21888
rect 0 21496 800 21616
rect 0 21224 800 21344
rect 0 20952 800 21072
rect 0 20680 800 20800
rect 0 20408 800 20528
rect 0 20136 800 20256
rect 0 19864 800 19984
rect 0 19592 800 19712
rect 0 19320 800 19440
rect 0 19048 800 19168
rect 0 18776 800 18896
rect 0 18504 800 18624
rect 0 18232 800 18352
rect 0 17960 800 18080
rect 0 17688 800 17808
rect 0 17416 800 17536
rect 0 17144 800 17264
rect 0 16872 800 16992
rect 0 16600 800 16720
rect 0 16328 800 16448
rect 69200 53048 70000 53168
rect 69200 52776 70000 52896
rect 69200 52504 70000 52624
rect 69200 52232 70000 52352
rect 69200 51960 70000 52080
rect 69200 51688 70000 51808
rect 69200 51416 70000 51536
rect 69200 51144 70000 51264
rect 69200 50872 70000 50992
rect 69200 50600 70000 50720
rect 69200 50328 70000 50448
rect 69200 50056 70000 50176
rect 69200 49784 70000 49904
rect 69200 49512 70000 49632
rect 69200 49240 70000 49360
rect 69200 48968 70000 49088
rect 69200 48696 70000 48816
rect 69200 48424 70000 48544
rect 69200 48152 70000 48272
rect 69200 47880 70000 48000
rect 69200 47608 70000 47728
rect 69200 47336 70000 47456
rect 69200 47064 70000 47184
rect 69200 46792 70000 46912
rect 69200 46520 70000 46640
rect 69200 46248 70000 46368
rect 69200 45976 70000 46096
rect 69200 45704 70000 45824
rect 69200 45432 70000 45552
rect 69200 45160 70000 45280
rect 69200 44888 70000 45008
rect 69200 44616 70000 44736
rect 69200 44344 70000 44464
rect 69200 44072 70000 44192
rect 69200 43800 70000 43920
rect 69200 43528 70000 43648
rect 69200 43256 70000 43376
rect 69200 42984 70000 43104
rect 69200 42712 70000 42832
rect 69200 42440 70000 42560
rect 69200 42168 70000 42288
rect 69200 41896 70000 42016
rect 69200 41624 70000 41744
rect 69200 41352 70000 41472
rect 69200 41080 70000 41200
rect 69200 40808 70000 40928
rect 69200 40536 70000 40656
rect 69200 40264 70000 40384
rect 69200 39992 70000 40112
rect 69200 39720 70000 39840
rect 69200 39448 70000 39568
rect 69200 39176 70000 39296
rect 69200 38904 70000 39024
rect 69200 38632 70000 38752
rect 69200 38360 70000 38480
rect 69200 38088 70000 38208
rect 69200 37816 70000 37936
rect 69200 37544 70000 37664
rect 69200 37272 70000 37392
rect 69200 37000 70000 37120
rect 69200 36728 70000 36848
rect 69200 36456 70000 36576
rect 69200 36184 70000 36304
rect 69200 35912 70000 36032
rect 69200 35640 70000 35760
rect 69200 35368 70000 35488
rect 69200 35096 70000 35216
rect 69200 34824 70000 34944
rect 69200 34552 70000 34672
rect 69200 34280 70000 34400
rect 69200 34008 70000 34128
rect 69200 33736 70000 33856
rect 69200 33464 70000 33584
rect 69200 33192 70000 33312
rect 69200 32920 70000 33040
rect 69200 32648 70000 32768
rect 69200 32376 70000 32496
rect 69200 32104 70000 32224
rect 69200 31832 70000 31952
rect 69200 31560 70000 31680
rect 69200 31288 70000 31408
rect 69200 31016 70000 31136
rect 69200 30744 70000 30864
rect 69200 30472 70000 30592
rect 69200 30200 70000 30320
rect 69200 29928 70000 30048
rect 69200 29656 70000 29776
rect 69200 29384 70000 29504
rect 69200 29112 70000 29232
rect 69200 28840 70000 28960
rect 69200 28568 70000 28688
rect 69200 28296 70000 28416
rect 69200 28024 70000 28144
rect 69200 27752 70000 27872
rect 69200 27480 70000 27600
rect 69200 27208 70000 27328
rect 69200 26936 70000 27056
rect 69200 26664 70000 26784
rect 69200 26392 70000 26512
rect 69200 26120 70000 26240
rect 69200 25848 70000 25968
rect 69200 25576 70000 25696
rect 69200 25304 70000 25424
rect 69200 25032 70000 25152
rect 69200 24760 70000 24880
rect 69200 24488 70000 24608
rect 69200 24216 70000 24336
rect 69200 23944 70000 24064
rect 69200 23672 70000 23792
rect 69200 23400 70000 23520
rect 69200 23128 70000 23248
rect 69200 22856 70000 22976
rect 69200 22584 70000 22704
rect 69200 22312 70000 22432
rect 69200 22040 70000 22160
rect 69200 21768 70000 21888
rect 69200 21496 70000 21616
rect 69200 21224 70000 21344
rect 69200 20952 70000 21072
rect 69200 20680 70000 20800
rect 69200 20408 70000 20528
rect 69200 20136 70000 20256
rect 69200 19864 70000 19984
rect 69200 19592 70000 19712
rect 69200 19320 70000 19440
rect 69200 19048 70000 19168
rect 69200 18776 70000 18896
rect 69200 18504 70000 18624
rect 69200 18232 70000 18352
rect 69200 17960 70000 18080
rect 69200 17688 70000 17808
rect 69200 17416 70000 17536
rect 69200 17144 70000 17264
rect 69200 16872 70000 16992
rect 69200 16600 70000 16720
rect 69200 16328 70000 16448
rect 0 16056 800 16176
rect 0 15784 800 15904
rect 0 15512 800 15632
rect 0 15240 800 15360
rect 0 14968 800 15088
rect 0 14696 800 14816
rect 0 14424 800 14544
rect 0 14152 800 14272
rect 0 13880 800 14000
rect 0 13608 800 13728
rect 0 13336 800 13456
rect 0 13064 800 13184
rect 0 12792 800 12912
rect 0 12520 800 12640
rect 0 12248 800 12368
rect 0 11976 800 12096
rect 0 11704 800 11824
rect 0 11432 800 11552
rect 0 11160 800 11280
rect 0 10888 800 11008
rect 0 10616 800 10736
rect 0 10344 800 10464
rect 0 10072 800 10192
rect 0 9800 800 9920
rect 0 9528 800 9648
rect 0 9256 800 9376
rect 0 8984 800 9104
rect 0 8712 800 8832
rect 0 8440 800 8560
rect 0 8168 800 8288
rect 0 7896 800 8016
rect 0 7624 800 7744
rect 0 7352 800 7472
rect 0 7080 800 7200
rect 0 6808 800 6928
rect 0 6536 800 6656
rect 0 6264 800 6384
rect 0 5992 800 6112
rect 0 5720 800 5840
rect 0 5448 800 5568
rect 0 5176 800 5296
rect 0 4904 800 5024
rect 0 4632 800 4752
rect 0 4360 800 4480
rect 0 4088 800 4208
rect 0 3816 800 3936
<< obsm3 >>
rect 800 65760 69200 69053
rect 880 53248 69200 65760
rect 880 16248 69120 53248
rect 880 3736 69200 16248
rect 800 2143 69200 3736
<< metal4 >>
rect 4208 2128 4528 67504
rect 19568 2128 19888 67504
rect 34928 2128 35248 67504
rect 50288 2128 50608 67504
rect 65648 2128 65968 67504
<< obsm4 >>
rect 614 67584 68941 68917
rect 614 4659 4128 67584
rect 4608 4659 19488 67584
rect 19968 4659 34848 67584
rect 35328 4659 50208 67584
rect 50688 4659 65568 67584
rect 66048 4659 68941 67584
<< labels >>
rlabel metal2 s 3330 69200 3386 70000 6 clk_i
port 1 nsew signal input
rlabel metal2 s 3882 69200 3938 70000 6 mports_i[0]
port 2 nsew signal input
rlabel metal2 s 31482 69200 31538 70000 6 mports_i[100]
port 3 nsew signal input
rlabel metal2 s 31758 69200 31814 70000 6 mports_i[101]
port 4 nsew signal input
rlabel metal2 s 32034 69200 32090 70000 6 mports_i[102]
port 5 nsew signal input
rlabel metal2 s 32310 69200 32366 70000 6 mports_i[103]
port 6 nsew signal input
rlabel metal2 s 32586 69200 32642 70000 6 mports_i[104]
port 7 nsew signal input
rlabel metal2 s 32862 69200 32918 70000 6 mports_i[105]
port 8 nsew signal input
rlabel metal2 s 33138 69200 33194 70000 6 mports_i[106]
port 9 nsew signal input
rlabel metal2 s 33414 69200 33470 70000 6 mports_i[107]
port 10 nsew signal input
rlabel metal2 s 33690 69200 33746 70000 6 mports_i[108]
port 11 nsew signal input
rlabel metal2 s 33966 69200 34022 70000 6 mports_i[109]
port 12 nsew signal input
rlabel metal2 s 6642 69200 6698 70000 6 mports_i[10]
port 13 nsew signal input
rlabel metal2 s 34242 69200 34298 70000 6 mports_i[110]
port 14 nsew signal input
rlabel metal2 s 34518 69200 34574 70000 6 mports_i[111]
port 15 nsew signal input
rlabel metal2 s 34794 69200 34850 70000 6 mports_i[112]
port 16 nsew signal input
rlabel metal2 s 35070 69200 35126 70000 6 mports_i[113]
port 17 nsew signal input
rlabel metal2 s 35346 69200 35402 70000 6 mports_i[114]
port 18 nsew signal input
rlabel metal2 s 35622 69200 35678 70000 6 mports_i[115]
port 19 nsew signal input
rlabel metal2 s 35898 69200 35954 70000 6 mports_i[116]
port 20 nsew signal input
rlabel metal2 s 36174 69200 36230 70000 6 mports_i[117]
port 21 nsew signal input
rlabel metal2 s 36450 69200 36506 70000 6 mports_i[118]
port 22 nsew signal input
rlabel metal2 s 36726 69200 36782 70000 6 mports_i[119]
port 23 nsew signal input
rlabel metal2 s 6918 69200 6974 70000 6 mports_i[11]
port 24 nsew signal input
rlabel metal2 s 37002 69200 37058 70000 6 mports_i[120]
port 25 nsew signal input
rlabel metal2 s 37278 69200 37334 70000 6 mports_i[121]
port 26 nsew signal input
rlabel metal2 s 37554 69200 37610 70000 6 mports_i[122]
port 27 nsew signal input
rlabel metal2 s 37830 69200 37886 70000 6 mports_i[123]
port 28 nsew signal input
rlabel metal2 s 38106 69200 38162 70000 6 mports_i[124]
port 29 nsew signal input
rlabel metal2 s 38382 69200 38438 70000 6 mports_i[125]
port 30 nsew signal input
rlabel metal2 s 38658 69200 38714 70000 6 mports_i[126]
port 31 nsew signal input
rlabel metal2 s 38934 69200 38990 70000 6 mports_i[127]
port 32 nsew signal input
rlabel metal2 s 39210 69200 39266 70000 6 mports_i[128]
port 33 nsew signal input
rlabel metal2 s 39486 69200 39542 70000 6 mports_i[129]
port 34 nsew signal input
rlabel metal2 s 7194 69200 7250 70000 6 mports_i[12]
port 35 nsew signal input
rlabel metal2 s 39762 69200 39818 70000 6 mports_i[130]
port 36 nsew signal input
rlabel metal2 s 40038 69200 40094 70000 6 mports_i[131]
port 37 nsew signal input
rlabel metal2 s 40314 69200 40370 70000 6 mports_i[132]
port 38 nsew signal input
rlabel metal2 s 40590 69200 40646 70000 6 mports_i[133]
port 39 nsew signal input
rlabel metal2 s 40866 69200 40922 70000 6 mports_i[134]
port 40 nsew signal input
rlabel metal2 s 41142 69200 41198 70000 6 mports_i[135]
port 41 nsew signal input
rlabel metal2 s 41418 69200 41474 70000 6 mports_i[136]
port 42 nsew signal input
rlabel metal2 s 41694 69200 41750 70000 6 mports_i[137]
port 43 nsew signal input
rlabel metal2 s 41970 69200 42026 70000 6 mports_i[138]
port 44 nsew signal input
rlabel metal2 s 42246 69200 42302 70000 6 mports_i[139]
port 45 nsew signal input
rlabel metal2 s 7470 69200 7526 70000 6 mports_i[13]
port 46 nsew signal input
rlabel metal2 s 42522 69200 42578 70000 6 mports_i[140]
port 47 nsew signal input
rlabel metal2 s 42798 69200 42854 70000 6 mports_i[141]
port 48 nsew signal input
rlabel metal2 s 43074 69200 43130 70000 6 mports_i[142]
port 49 nsew signal input
rlabel metal2 s 43350 69200 43406 70000 6 mports_i[143]
port 50 nsew signal input
rlabel metal2 s 43626 69200 43682 70000 6 mports_i[144]
port 51 nsew signal input
rlabel metal2 s 43902 69200 43958 70000 6 mports_i[145]
port 52 nsew signal input
rlabel metal2 s 44178 69200 44234 70000 6 mports_i[146]
port 53 nsew signal input
rlabel metal2 s 44454 69200 44510 70000 6 mports_i[147]
port 54 nsew signal input
rlabel metal2 s 44730 69200 44786 70000 6 mports_i[148]
port 55 nsew signal input
rlabel metal2 s 45006 69200 45062 70000 6 mports_i[149]
port 56 nsew signal input
rlabel metal2 s 7746 69200 7802 70000 6 mports_i[14]
port 57 nsew signal input
rlabel metal2 s 45282 69200 45338 70000 6 mports_i[150]
port 58 nsew signal input
rlabel metal2 s 45558 69200 45614 70000 6 mports_i[151]
port 59 nsew signal input
rlabel metal2 s 45834 69200 45890 70000 6 mports_i[152]
port 60 nsew signal input
rlabel metal2 s 46110 69200 46166 70000 6 mports_i[153]
port 61 nsew signal input
rlabel metal2 s 46386 69200 46442 70000 6 mports_i[154]
port 62 nsew signal input
rlabel metal2 s 46662 69200 46718 70000 6 mports_i[155]
port 63 nsew signal input
rlabel metal2 s 46938 69200 46994 70000 6 mports_i[156]
port 64 nsew signal input
rlabel metal2 s 47214 69200 47270 70000 6 mports_i[157]
port 65 nsew signal input
rlabel metal2 s 47490 69200 47546 70000 6 mports_i[158]
port 66 nsew signal input
rlabel metal2 s 47766 69200 47822 70000 6 mports_i[159]
port 67 nsew signal input
rlabel metal2 s 8022 69200 8078 70000 6 mports_i[15]
port 68 nsew signal input
rlabel metal2 s 48042 69200 48098 70000 6 mports_i[160]
port 69 nsew signal input
rlabel metal2 s 48318 69200 48374 70000 6 mports_i[161]
port 70 nsew signal input
rlabel metal2 s 48594 69200 48650 70000 6 mports_i[162]
port 71 nsew signal input
rlabel metal2 s 48870 69200 48926 70000 6 mports_i[163]
port 72 nsew signal input
rlabel metal2 s 49146 69200 49202 70000 6 mports_i[164]
port 73 nsew signal input
rlabel metal2 s 49422 69200 49478 70000 6 mports_i[165]
port 74 nsew signal input
rlabel metal2 s 49698 69200 49754 70000 6 mports_i[166]
port 75 nsew signal input
rlabel metal2 s 49974 69200 50030 70000 6 mports_i[167]
port 76 nsew signal input
rlabel metal2 s 50250 69200 50306 70000 6 mports_i[168]
port 77 nsew signal input
rlabel metal2 s 50526 69200 50582 70000 6 mports_i[169]
port 78 nsew signal input
rlabel metal2 s 8298 69200 8354 70000 6 mports_i[16]
port 79 nsew signal input
rlabel metal2 s 50802 69200 50858 70000 6 mports_i[170]
port 80 nsew signal input
rlabel metal2 s 51078 69200 51134 70000 6 mports_i[171]
port 81 nsew signal input
rlabel metal2 s 51354 69200 51410 70000 6 mports_i[172]
port 82 nsew signal input
rlabel metal2 s 51630 69200 51686 70000 6 mports_i[173]
port 83 nsew signal input
rlabel metal2 s 51906 69200 51962 70000 6 mports_i[174]
port 84 nsew signal input
rlabel metal2 s 52182 69200 52238 70000 6 mports_i[175]
port 85 nsew signal input
rlabel metal2 s 52458 69200 52514 70000 6 mports_i[176]
port 86 nsew signal input
rlabel metal2 s 52734 69200 52790 70000 6 mports_i[177]
port 87 nsew signal input
rlabel metal2 s 53010 69200 53066 70000 6 mports_i[178]
port 88 nsew signal input
rlabel metal2 s 53286 69200 53342 70000 6 mports_i[179]
port 89 nsew signal input
rlabel metal2 s 8574 69200 8630 70000 6 mports_i[17]
port 90 nsew signal input
rlabel metal2 s 53562 69200 53618 70000 6 mports_i[180]
port 91 nsew signal input
rlabel metal2 s 53838 69200 53894 70000 6 mports_i[181]
port 92 nsew signal input
rlabel metal2 s 54114 69200 54170 70000 6 mports_i[182]
port 93 nsew signal input
rlabel metal2 s 54390 69200 54446 70000 6 mports_i[183]
port 94 nsew signal input
rlabel metal2 s 54666 69200 54722 70000 6 mports_i[184]
port 95 nsew signal input
rlabel metal2 s 54942 69200 54998 70000 6 mports_i[185]
port 96 nsew signal input
rlabel metal2 s 55218 69200 55274 70000 6 mports_i[186]
port 97 nsew signal input
rlabel metal2 s 55494 69200 55550 70000 6 mports_i[187]
port 98 nsew signal input
rlabel metal2 s 55770 69200 55826 70000 6 mports_i[188]
port 99 nsew signal input
rlabel metal2 s 56046 69200 56102 70000 6 mports_i[189]
port 100 nsew signal input
rlabel metal2 s 8850 69200 8906 70000 6 mports_i[18]
port 101 nsew signal input
rlabel metal2 s 56322 69200 56378 70000 6 mports_i[190]
port 102 nsew signal input
rlabel metal2 s 56598 69200 56654 70000 6 mports_i[191]
port 103 nsew signal input
rlabel metal2 s 56874 69200 56930 70000 6 mports_i[192]
port 104 nsew signal input
rlabel metal2 s 57150 69200 57206 70000 6 mports_i[193]
port 105 nsew signal input
rlabel metal2 s 57426 69200 57482 70000 6 mports_i[194]
port 106 nsew signal input
rlabel metal2 s 57702 69200 57758 70000 6 mports_i[195]
port 107 nsew signal input
rlabel metal2 s 57978 69200 58034 70000 6 mports_i[196]
port 108 nsew signal input
rlabel metal2 s 58254 69200 58310 70000 6 mports_i[197]
port 109 nsew signal input
rlabel metal2 s 58530 69200 58586 70000 6 mports_i[198]
port 110 nsew signal input
rlabel metal2 s 58806 69200 58862 70000 6 mports_i[199]
port 111 nsew signal input
rlabel metal2 s 9126 69200 9182 70000 6 mports_i[19]
port 112 nsew signal input
rlabel metal2 s 4158 69200 4214 70000 6 mports_i[1]
port 113 nsew signal input
rlabel metal2 s 59082 69200 59138 70000 6 mports_i[200]
port 114 nsew signal input
rlabel metal2 s 59358 69200 59414 70000 6 mports_i[201]
port 115 nsew signal input
rlabel metal2 s 59634 69200 59690 70000 6 mports_i[202]
port 116 nsew signal input
rlabel metal2 s 59910 69200 59966 70000 6 mports_i[203]
port 117 nsew signal input
rlabel metal2 s 60186 69200 60242 70000 6 mports_i[204]
port 118 nsew signal input
rlabel metal2 s 60462 69200 60518 70000 6 mports_i[205]
port 119 nsew signal input
rlabel metal2 s 60738 69200 60794 70000 6 mports_i[206]
port 120 nsew signal input
rlabel metal2 s 61014 69200 61070 70000 6 mports_i[207]
port 121 nsew signal input
rlabel metal2 s 61290 69200 61346 70000 6 mports_i[208]
port 122 nsew signal input
rlabel metal2 s 61566 69200 61622 70000 6 mports_i[209]
port 123 nsew signal input
rlabel metal2 s 9402 69200 9458 70000 6 mports_i[20]
port 124 nsew signal input
rlabel metal2 s 61842 69200 61898 70000 6 mports_i[210]
port 125 nsew signal input
rlabel metal2 s 62118 69200 62174 70000 6 mports_i[211]
port 126 nsew signal input
rlabel metal2 s 62394 69200 62450 70000 6 mports_i[212]
port 127 nsew signal input
rlabel metal2 s 62670 69200 62726 70000 6 mports_i[213]
port 128 nsew signal input
rlabel metal2 s 62946 69200 63002 70000 6 mports_i[214]
port 129 nsew signal input
rlabel metal2 s 63222 69200 63278 70000 6 mports_i[215]
port 130 nsew signal input
rlabel metal2 s 63498 69200 63554 70000 6 mports_i[216]
port 131 nsew signal input
rlabel metal2 s 63774 69200 63830 70000 6 mports_i[217]
port 132 nsew signal input
rlabel metal2 s 64050 69200 64106 70000 6 mports_i[218]
port 133 nsew signal input
rlabel metal2 s 64326 69200 64382 70000 6 mports_i[219]
port 134 nsew signal input
rlabel metal2 s 9678 69200 9734 70000 6 mports_i[21]
port 135 nsew signal input
rlabel metal2 s 64602 69200 64658 70000 6 mports_i[220]
port 136 nsew signal input
rlabel metal2 s 64878 69200 64934 70000 6 mports_i[221]
port 137 nsew signal input
rlabel metal2 s 65154 69200 65210 70000 6 mports_i[222]
port 138 nsew signal input
rlabel metal2 s 65430 69200 65486 70000 6 mports_i[223]
port 139 nsew signal input
rlabel metal2 s 65706 69200 65762 70000 6 mports_i[224]
port 140 nsew signal input
rlabel metal2 s 65982 69200 66038 70000 6 mports_i[225]
port 141 nsew signal input
rlabel metal2 s 66258 69200 66314 70000 6 mports_i[226]
port 142 nsew signal input
rlabel metal2 s 66534 69200 66590 70000 6 mports_i[227]
port 143 nsew signal input
rlabel metal2 s 9954 69200 10010 70000 6 mports_i[22]
port 144 nsew signal input
rlabel metal2 s 10230 69200 10286 70000 6 mports_i[23]
port 145 nsew signal input
rlabel metal2 s 10506 69200 10562 70000 6 mports_i[24]
port 146 nsew signal input
rlabel metal2 s 10782 69200 10838 70000 6 mports_i[25]
port 147 nsew signal input
rlabel metal2 s 11058 69200 11114 70000 6 mports_i[26]
port 148 nsew signal input
rlabel metal2 s 11334 69200 11390 70000 6 mports_i[27]
port 149 nsew signal input
rlabel metal2 s 11610 69200 11666 70000 6 mports_i[28]
port 150 nsew signal input
rlabel metal2 s 11886 69200 11942 70000 6 mports_i[29]
port 151 nsew signal input
rlabel metal2 s 4434 69200 4490 70000 6 mports_i[2]
port 152 nsew signal input
rlabel metal2 s 12162 69200 12218 70000 6 mports_i[30]
port 153 nsew signal input
rlabel metal2 s 12438 69200 12494 70000 6 mports_i[31]
port 154 nsew signal input
rlabel metal2 s 12714 69200 12770 70000 6 mports_i[32]
port 155 nsew signal input
rlabel metal2 s 12990 69200 13046 70000 6 mports_i[33]
port 156 nsew signal input
rlabel metal2 s 13266 69200 13322 70000 6 mports_i[34]
port 157 nsew signal input
rlabel metal2 s 13542 69200 13598 70000 6 mports_i[35]
port 158 nsew signal input
rlabel metal2 s 13818 69200 13874 70000 6 mports_i[36]
port 159 nsew signal input
rlabel metal2 s 14094 69200 14150 70000 6 mports_i[37]
port 160 nsew signal input
rlabel metal2 s 14370 69200 14426 70000 6 mports_i[38]
port 161 nsew signal input
rlabel metal2 s 14646 69200 14702 70000 6 mports_i[39]
port 162 nsew signal input
rlabel metal2 s 4710 69200 4766 70000 6 mports_i[3]
port 163 nsew signal input
rlabel metal2 s 14922 69200 14978 70000 6 mports_i[40]
port 164 nsew signal input
rlabel metal2 s 15198 69200 15254 70000 6 mports_i[41]
port 165 nsew signal input
rlabel metal2 s 15474 69200 15530 70000 6 mports_i[42]
port 166 nsew signal input
rlabel metal2 s 15750 69200 15806 70000 6 mports_i[43]
port 167 nsew signal input
rlabel metal2 s 16026 69200 16082 70000 6 mports_i[44]
port 168 nsew signal input
rlabel metal2 s 16302 69200 16358 70000 6 mports_i[45]
port 169 nsew signal input
rlabel metal2 s 16578 69200 16634 70000 6 mports_i[46]
port 170 nsew signal input
rlabel metal2 s 16854 69200 16910 70000 6 mports_i[47]
port 171 nsew signal input
rlabel metal2 s 17130 69200 17186 70000 6 mports_i[48]
port 172 nsew signal input
rlabel metal2 s 17406 69200 17462 70000 6 mports_i[49]
port 173 nsew signal input
rlabel metal2 s 4986 69200 5042 70000 6 mports_i[4]
port 174 nsew signal input
rlabel metal2 s 17682 69200 17738 70000 6 mports_i[50]
port 175 nsew signal input
rlabel metal2 s 17958 69200 18014 70000 6 mports_i[51]
port 176 nsew signal input
rlabel metal2 s 18234 69200 18290 70000 6 mports_i[52]
port 177 nsew signal input
rlabel metal2 s 18510 69200 18566 70000 6 mports_i[53]
port 178 nsew signal input
rlabel metal2 s 18786 69200 18842 70000 6 mports_i[54]
port 179 nsew signal input
rlabel metal2 s 19062 69200 19118 70000 6 mports_i[55]
port 180 nsew signal input
rlabel metal2 s 19338 69200 19394 70000 6 mports_i[56]
port 181 nsew signal input
rlabel metal2 s 19614 69200 19670 70000 6 mports_i[57]
port 182 nsew signal input
rlabel metal2 s 19890 69200 19946 70000 6 mports_i[58]
port 183 nsew signal input
rlabel metal2 s 20166 69200 20222 70000 6 mports_i[59]
port 184 nsew signal input
rlabel metal2 s 5262 69200 5318 70000 6 mports_i[5]
port 185 nsew signal input
rlabel metal2 s 20442 69200 20498 70000 6 mports_i[60]
port 186 nsew signal input
rlabel metal2 s 20718 69200 20774 70000 6 mports_i[61]
port 187 nsew signal input
rlabel metal2 s 20994 69200 21050 70000 6 mports_i[62]
port 188 nsew signal input
rlabel metal2 s 21270 69200 21326 70000 6 mports_i[63]
port 189 nsew signal input
rlabel metal2 s 21546 69200 21602 70000 6 mports_i[64]
port 190 nsew signal input
rlabel metal2 s 21822 69200 21878 70000 6 mports_i[65]
port 191 nsew signal input
rlabel metal2 s 22098 69200 22154 70000 6 mports_i[66]
port 192 nsew signal input
rlabel metal2 s 22374 69200 22430 70000 6 mports_i[67]
port 193 nsew signal input
rlabel metal2 s 22650 69200 22706 70000 6 mports_i[68]
port 194 nsew signal input
rlabel metal2 s 22926 69200 22982 70000 6 mports_i[69]
port 195 nsew signal input
rlabel metal2 s 5538 69200 5594 70000 6 mports_i[6]
port 196 nsew signal input
rlabel metal2 s 23202 69200 23258 70000 6 mports_i[70]
port 197 nsew signal input
rlabel metal2 s 23478 69200 23534 70000 6 mports_i[71]
port 198 nsew signal input
rlabel metal2 s 23754 69200 23810 70000 6 mports_i[72]
port 199 nsew signal input
rlabel metal2 s 24030 69200 24086 70000 6 mports_i[73]
port 200 nsew signal input
rlabel metal2 s 24306 69200 24362 70000 6 mports_i[74]
port 201 nsew signal input
rlabel metal2 s 24582 69200 24638 70000 6 mports_i[75]
port 202 nsew signal input
rlabel metal2 s 24858 69200 24914 70000 6 mports_i[76]
port 203 nsew signal input
rlabel metal2 s 25134 69200 25190 70000 6 mports_i[77]
port 204 nsew signal input
rlabel metal2 s 25410 69200 25466 70000 6 mports_i[78]
port 205 nsew signal input
rlabel metal2 s 25686 69200 25742 70000 6 mports_i[79]
port 206 nsew signal input
rlabel metal2 s 5814 69200 5870 70000 6 mports_i[7]
port 207 nsew signal input
rlabel metal2 s 25962 69200 26018 70000 6 mports_i[80]
port 208 nsew signal input
rlabel metal2 s 26238 69200 26294 70000 6 mports_i[81]
port 209 nsew signal input
rlabel metal2 s 26514 69200 26570 70000 6 mports_i[82]
port 210 nsew signal input
rlabel metal2 s 26790 69200 26846 70000 6 mports_i[83]
port 211 nsew signal input
rlabel metal2 s 27066 69200 27122 70000 6 mports_i[84]
port 212 nsew signal input
rlabel metal2 s 27342 69200 27398 70000 6 mports_i[85]
port 213 nsew signal input
rlabel metal2 s 27618 69200 27674 70000 6 mports_i[86]
port 214 nsew signal input
rlabel metal2 s 27894 69200 27950 70000 6 mports_i[87]
port 215 nsew signal input
rlabel metal2 s 28170 69200 28226 70000 6 mports_i[88]
port 216 nsew signal input
rlabel metal2 s 28446 69200 28502 70000 6 mports_i[89]
port 217 nsew signal input
rlabel metal2 s 6090 69200 6146 70000 6 mports_i[8]
port 218 nsew signal input
rlabel metal2 s 28722 69200 28778 70000 6 mports_i[90]
port 219 nsew signal input
rlabel metal2 s 28998 69200 29054 70000 6 mports_i[91]
port 220 nsew signal input
rlabel metal2 s 29274 69200 29330 70000 6 mports_i[92]
port 221 nsew signal input
rlabel metal2 s 29550 69200 29606 70000 6 mports_i[93]
port 222 nsew signal input
rlabel metal2 s 29826 69200 29882 70000 6 mports_i[94]
port 223 nsew signal input
rlabel metal2 s 30102 69200 30158 70000 6 mports_i[95]
port 224 nsew signal input
rlabel metal2 s 30378 69200 30434 70000 6 mports_i[96]
port 225 nsew signal input
rlabel metal2 s 30654 69200 30710 70000 6 mports_i[97]
port 226 nsew signal input
rlabel metal2 s 30930 69200 30986 70000 6 mports_i[98]
port 227 nsew signal input
rlabel metal2 s 31206 69200 31262 70000 6 mports_i[99]
port 228 nsew signal input
rlabel metal2 s 6366 69200 6422 70000 6 mports_i[9]
port 229 nsew signal input
rlabel metal2 s 3882 0 3938 800 6 mports_o[0]
port 230 nsew signal output
rlabel metal2 s 49882 0 49938 800 6 mports_o[100]
port 231 nsew signal output
rlabel metal2 s 50342 0 50398 800 6 mports_o[101]
port 232 nsew signal output
rlabel metal2 s 50802 0 50858 800 6 mports_o[102]
port 233 nsew signal output
rlabel metal2 s 51262 0 51318 800 6 mports_o[103]
port 234 nsew signal output
rlabel metal2 s 51722 0 51778 800 6 mports_o[104]
port 235 nsew signal output
rlabel metal2 s 52182 0 52238 800 6 mports_o[105]
port 236 nsew signal output
rlabel metal2 s 52642 0 52698 800 6 mports_o[106]
port 237 nsew signal output
rlabel metal2 s 53102 0 53158 800 6 mports_o[107]
port 238 nsew signal output
rlabel metal2 s 53562 0 53618 800 6 mports_o[108]
port 239 nsew signal output
rlabel metal2 s 54022 0 54078 800 6 mports_o[109]
port 240 nsew signal output
rlabel metal2 s 8482 0 8538 800 6 mports_o[10]
port 241 nsew signal output
rlabel metal2 s 54482 0 54538 800 6 mports_o[110]
port 242 nsew signal output
rlabel metal2 s 54942 0 54998 800 6 mports_o[111]
port 243 nsew signal output
rlabel metal2 s 55402 0 55458 800 6 mports_o[112]
port 244 nsew signal output
rlabel metal2 s 55862 0 55918 800 6 mports_o[113]
port 245 nsew signal output
rlabel metal2 s 56322 0 56378 800 6 mports_o[114]
port 246 nsew signal output
rlabel metal2 s 56782 0 56838 800 6 mports_o[115]
port 247 nsew signal output
rlabel metal2 s 57242 0 57298 800 6 mports_o[116]
port 248 nsew signal output
rlabel metal2 s 57702 0 57758 800 6 mports_o[117]
port 249 nsew signal output
rlabel metal2 s 58162 0 58218 800 6 mports_o[118]
port 250 nsew signal output
rlabel metal2 s 58622 0 58678 800 6 mports_o[119]
port 251 nsew signal output
rlabel metal2 s 8942 0 8998 800 6 mports_o[11]
port 252 nsew signal output
rlabel metal2 s 59082 0 59138 800 6 mports_o[120]
port 253 nsew signal output
rlabel metal2 s 59542 0 59598 800 6 mports_o[121]
port 254 nsew signal output
rlabel metal2 s 60002 0 60058 800 6 mports_o[122]
port 255 nsew signal output
rlabel metal2 s 60462 0 60518 800 6 mports_o[123]
port 256 nsew signal output
rlabel metal2 s 60922 0 60978 800 6 mports_o[124]
port 257 nsew signal output
rlabel metal2 s 61382 0 61438 800 6 mports_o[125]
port 258 nsew signal output
rlabel metal2 s 61842 0 61898 800 6 mports_o[126]
port 259 nsew signal output
rlabel metal2 s 62302 0 62358 800 6 mports_o[127]
port 260 nsew signal output
rlabel metal2 s 62762 0 62818 800 6 mports_o[128]
port 261 nsew signal output
rlabel metal2 s 63222 0 63278 800 6 mports_o[129]
port 262 nsew signal output
rlabel metal2 s 9402 0 9458 800 6 mports_o[12]
port 263 nsew signal output
rlabel metal2 s 63682 0 63738 800 6 mports_o[130]
port 264 nsew signal output
rlabel metal2 s 64142 0 64198 800 6 mports_o[131]
port 265 nsew signal output
rlabel metal2 s 64602 0 64658 800 6 mports_o[132]
port 266 nsew signal output
rlabel metal2 s 65062 0 65118 800 6 mports_o[133]
port 267 nsew signal output
rlabel metal2 s 65522 0 65578 800 6 mports_o[134]
port 268 nsew signal output
rlabel metal2 s 65982 0 66038 800 6 mports_o[135]
port 269 nsew signal output
rlabel metal2 s 9862 0 9918 800 6 mports_o[13]
port 270 nsew signal output
rlabel metal2 s 10322 0 10378 800 6 mports_o[14]
port 271 nsew signal output
rlabel metal2 s 10782 0 10838 800 6 mports_o[15]
port 272 nsew signal output
rlabel metal2 s 11242 0 11298 800 6 mports_o[16]
port 273 nsew signal output
rlabel metal2 s 11702 0 11758 800 6 mports_o[17]
port 274 nsew signal output
rlabel metal2 s 12162 0 12218 800 6 mports_o[18]
port 275 nsew signal output
rlabel metal2 s 12622 0 12678 800 6 mports_o[19]
port 276 nsew signal output
rlabel metal2 s 4342 0 4398 800 6 mports_o[1]
port 277 nsew signal output
rlabel metal2 s 13082 0 13138 800 6 mports_o[20]
port 278 nsew signal output
rlabel metal2 s 13542 0 13598 800 6 mports_o[21]
port 279 nsew signal output
rlabel metal2 s 14002 0 14058 800 6 mports_o[22]
port 280 nsew signal output
rlabel metal2 s 14462 0 14518 800 6 mports_o[23]
port 281 nsew signal output
rlabel metal2 s 14922 0 14978 800 6 mports_o[24]
port 282 nsew signal output
rlabel metal2 s 15382 0 15438 800 6 mports_o[25]
port 283 nsew signal output
rlabel metal2 s 15842 0 15898 800 6 mports_o[26]
port 284 nsew signal output
rlabel metal2 s 16302 0 16358 800 6 mports_o[27]
port 285 nsew signal output
rlabel metal2 s 16762 0 16818 800 6 mports_o[28]
port 286 nsew signal output
rlabel metal2 s 17222 0 17278 800 6 mports_o[29]
port 287 nsew signal output
rlabel metal2 s 4802 0 4858 800 6 mports_o[2]
port 288 nsew signal output
rlabel metal2 s 17682 0 17738 800 6 mports_o[30]
port 289 nsew signal output
rlabel metal2 s 18142 0 18198 800 6 mports_o[31]
port 290 nsew signal output
rlabel metal2 s 18602 0 18658 800 6 mports_o[32]
port 291 nsew signal output
rlabel metal2 s 19062 0 19118 800 6 mports_o[33]
port 292 nsew signal output
rlabel metal2 s 19522 0 19578 800 6 mports_o[34]
port 293 nsew signal output
rlabel metal2 s 19982 0 20038 800 6 mports_o[35]
port 294 nsew signal output
rlabel metal2 s 20442 0 20498 800 6 mports_o[36]
port 295 nsew signal output
rlabel metal2 s 20902 0 20958 800 6 mports_o[37]
port 296 nsew signal output
rlabel metal2 s 21362 0 21418 800 6 mports_o[38]
port 297 nsew signal output
rlabel metal2 s 21822 0 21878 800 6 mports_o[39]
port 298 nsew signal output
rlabel metal2 s 5262 0 5318 800 6 mports_o[3]
port 299 nsew signal output
rlabel metal2 s 22282 0 22338 800 6 mports_o[40]
port 300 nsew signal output
rlabel metal2 s 22742 0 22798 800 6 mports_o[41]
port 301 nsew signal output
rlabel metal2 s 23202 0 23258 800 6 mports_o[42]
port 302 nsew signal output
rlabel metal2 s 23662 0 23718 800 6 mports_o[43]
port 303 nsew signal output
rlabel metal2 s 24122 0 24178 800 6 mports_o[44]
port 304 nsew signal output
rlabel metal2 s 24582 0 24638 800 6 mports_o[45]
port 305 nsew signal output
rlabel metal2 s 25042 0 25098 800 6 mports_o[46]
port 306 nsew signal output
rlabel metal2 s 25502 0 25558 800 6 mports_o[47]
port 307 nsew signal output
rlabel metal2 s 25962 0 26018 800 6 mports_o[48]
port 308 nsew signal output
rlabel metal2 s 26422 0 26478 800 6 mports_o[49]
port 309 nsew signal output
rlabel metal2 s 5722 0 5778 800 6 mports_o[4]
port 310 nsew signal output
rlabel metal2 s 26882 0 26938 800 6 mports_o[50]
port 311 nsew signal output
rlabel metal2 s 27342 0 27398 800 6 mports_o[51]
port 312 nsew signal output
rlabel metal2 s 27802 0 27858 800 6 mports_o[52]
port 313 nsew signal output
rlabel metal2 s 28262 0 28318 800 6 mports_o[53]
port 314 nsew signal output
rlabel metal2 s 28722 0 28778 800 6 mports_o[54]
port 315 nsew signal output
rlabel metal2 s 29182 0 29238 800 6 mports_o[55]
port 316 nsew signal output
rlabel metal2 s 29642 0 29698 800 6 mports_o[56]
port 317 nsew signal output
rlabel metal2 s 30102 0 30158 800 6 mports_o[57]
port 318 nsew signal output
rlabel metal2 s 30562 0 30618 800 6 mports_o[58]
port 319 nsew signal output
rlabel metal2 s 31022 0 31078 800 6 mports_o[59]
port 320 nsew signal output
rlabel metal2 s 6182 0 6238 800 6 mports_o[5]
port 321 nsew signal output
rlabel metal2 s 31482 0 31538 800 6 mports_o[60]
port 322 nsew signal output
rlabel metal2 s 31942 0 31998 800 6 mports_o[61]
port 323 nsew signal output
rlabel metal2 s 32402 0 32458 800 6 mports_o[62]
port 324 nsew signal output
rlabel metal2 s 32862 0 32918 800 6 mports_o[63]
port 325 nsew signal output
rlabel metal2 s 33322 0 33378 800 6 mports_o[64]
port 326 nsew signal output
rlabel metal2 s 33782 0 33838 800 6 mports_o[65]
port 327 nsew signal output
rlabel metal2 s 34242 0 34298 800 6 mports_o[66]
port 328 nsew signal output
rlabel metal2 s 34702 0 34758 800 6 mports_o[67]
port 329 nsew signal output
rlabel metal2 s 35162 0 35218 800 6 mports_o[68]
port 330 nsew signal output
rlabel metal2 s 35622 0 35678 800 6 mports_o[69]
port 331 nsew signal output
rlabel metal2 s 6642 0 6698 800 6 mports_o[6]
port 332 nsew signal output
rlabel metal2 s 36082 0 36138 800 6 mports_o[70]
port 333 nsew signal output
rlabel metal2 s 36542 0 36598 800 6 mports_o[71]
port 334 nsew signal output
rlabel metal2 s 37002 0 37058 800 6 mports_o[72]
port 335 nsew signal output
rlabel metal2 s 37462 0 37518 800 6 mports_o[73]
port 336 nsew signal output
rlabel metal2 s 37922 0 37978 800 6 mports_o[74]
port 337 nsew signal output
rlabel metal2 s 38382 0 38438 800 6 mports_o[75]
port 338 nsew signal output
rlabel metal2 s 38842 0 38898 800 6 mports_o[76]
port 339 nsew signal output
rlabel metal2 s 39302 0 39358 800 6 mports_o[77]
port 340 nsew signal output
rlabel metal2 s 39762 0 39818 800 6 mports_o[78]
port 341 nsew signal output
rlabel metal2 s 40222 0 40278 800 6 mports_o[79]
port 342 nsew signal output
rlabel metal2 s 7102 0 7158 800 6 mports_o[7]
port 343 nsew signal output
rlabel metal2 s 40682 0 40738 800 6 mports_o[80]
port 344 nsew signal output
rlabel metal2 s 41142 0 41198 800 6 mports_o[81]
port 345 nsew signal output
rlabel metal2 s 41602 0 41658 800 6 mports_o[82]
port 346 nsew signal output
rlabel metal2 s 42062 0 42118 800 6 mports_o[83]
port 347 nsew signal output
rlabel metal2 s 42522 0 42578 800 6 mports_o[84]
port 348 nsew signal output
rlabel metal2 s 42982 0 43038 800 6 mports_o[85]
port 349 nsew signal output
rlabel metal2 s 43442 0 43498 800 6 mports_o[86]
port 350 nsew signal output
rlabel metal2 s 43902 0 43958 800 6 mports_o[87]
port 351 nsew signal output
rlabel metal2 s 44362 0 44418 800 6 mports_o[88]
port 352 nsew signal output
rlabel metal2 s 44822 0 44878 800 6 mports_o[89]
port 353 nsew signal output
rlabel metal2 s 7562 0 7618 800 6 mports_o[8]
port 354 nsew signal output
rlabel metal2 s 45282 0 45338 800 6 mports_o[90]
port 355 nsew signal output
rlabel metal2 s 45742 0 45798 800 6 mports_o[91]
port 356 nsew signal output
rlabel metal2 s 46202 0 46258 800 6 mports_o[92]
port 357 nsew signal output
rlabel metal2 s 46662 0 46718 800 6 mports_o[93]
port 358 nsew signal output
rlabel metal2 s 47122 0 47178 800 6 mports_o[94]
port 359 nsew signal output
rlabel metal2 s 47582 0 47638 800 6 mports_o[95]
port 360 nsew signal output
rlabel metal2 s 48042 0 48098 800 6 mports_o[96]
port 361 nsew signal output
rlabel metal2 s 48502 0 48558 800 6 mports_o[97]
port 362 nsew signal output
rlabel metal2 s 48962 0 49018 800 6 mports_o[98]
port 363 nsew signal output
rlabel metal2 s 49422 0 49478 800 6 mports_o[99]
port 364 nsew signal output
rlabel metal2 s 8022 0 8078 800 6 mports_o[9]
port 365 nsew signal output
rlabel metal2 s 3606 69200 3662 70000 6 nrst_i
port 366 nsew signal input
rlabel metal3 s 69200 16328 70000 16448 6 sports_i[0]
port 367 nsew signal input
rlabel metal3 s 69200 43528 70000 43648 6 sports_i[100]
port 368 nsew signal input
rlabel metal3 s 69200 43800 70000 43920 6 sports_i[101]
port 369 nsew signal input
rlabel metal3 s 69200 44072 70000 44192 6 sports_i[102]
port 370 nsew signal input
rlabel metal3 s 69200 44344 70000 44464 6 sports_i[103]
port 371 nsew signal input
rlabel metal3 s 69200 44616 70000 44736 6 sports_i[104]
port 372 nsew signal input
rlabel metal3 s 69200 44888 70000 45008 6 sports_i[105]
port 373 nsew signal input
rlabel metal3 s 69200 45160 70000 45280 6 sports_i[106]
port 374 nsew signal input
rlabel metal3 s 69200 45432 70000 45552 6 sports_i[107]
port 375 nsew signal input
rlabel metal3 s 69200 45704 70000 45824 6 sports_i[108]
port 376 nsew signal input
rlabel metal3 s 69200 45976 70000 46096 6 sports_i[109]
port 377 nsew signal input
rlabel metal3 s 69200 19048 70000 19168 6 sports_i[10]
port 378 nsew signal input
rlabel metal3 s 69200 46248 70000 46368 6 sports_i[110]
port 379 nsew signal input
rlabel metal3 s 69200 46520 70000 46640 6 sports_i[111]
port 380 nsew signal input
rlabel metal3 s 69200 46792 70000 46912 6 sports_i[112]
port 381 nsew signal input
rlabel metal3 s 69200 47064 70000 47184 6 sports_i[113]
port 382 nsew signal input
rlabel metal3 s 69200 47336 70000 47456 6 sports_i[114]
port 383 nsew signal input
rlabel metal3 s 69200 47608 70000 47728 6 sports_i[115]
port 384 nsew signal input
rlabel metal3 s 69200 47880 70000 48000 6 sports_i[116]
port 385 nsew signal input
rlabel metal3 s 69200 48152 70000 48272 6 sports_i[117]
port 386 nsew signal input
rlabel metal3 s 69200 48424 70000 48544 6 sports_i[118]
port 387 nsew signal input
rlabel metal3 s 69200 48696 70000 48816 6 sports_i[119]
port 388 nsew signal input
rlabel metal3 s 69200 19320 70000 19440 6 sports_i[11]
port 389 nsew signal input
rlabel metal3 s 69200 48968 70000 49088 6 sports_i[120]
port 390 nsew signal input
rlabel metal3 s 69200 49240 70000 49360 6 sports_i[121]
port 391 nsew signal input
rlabel metal3 s 69200 49512 70000 49632 6 sports_i[122]
port 392 nsew signal input
rlabel metal3 s 69200 49784 70000 49904 6 sports_i[123]
port 393 nsew signal input
rlabel metal3 s 69200 50056 70000 50176 6 sports_i[124]
port 394 nsew signal input
rlabel metal3 s 69200 50328 70000 50448 6 sports_i[125]
port 395 nsew signal input
rlabel metal3 s 69200 50600 70000 50720 6 sports_i[126]
port 396 nsew signal input
rlabel metal3 s 69200 50872 70000 50992 6 sports_i[127]
port 397 nsew signal input
rlabel metal3 s 69200 51144 70000 51264 6 sports_i[128]
port 398 nsew signal input
rlabel metal3 s 69200 51416 70000 51536 6 sports_i[129]
port 399 nsew signal input
rlabel metal3 s 69200 19592 70000 19712 6 sports_i[12]
port 400 nsew signal input
rlabel metal3 s 69200 51688 70000 51808 6 sports_i[130]
port 401 nsew signal input
rlabel metal3 s 69200 51960 70000 52080 6 sports_i[131]
port 402 nsew signal input
rlabel metal3 s 69200 52232 70000 52352 6 sports_i[132]
port 403 nsew signal input
rlabel metal3 s 69200 52504 70000 52624 6 sports_i[133]
port 404 nsew signal input
rlabel metal3 s 69200 52776 70000 52896 6 sports_i[134]
port 405 nsew signal input
rlabel metal3 s 69200 53048 70000 53168 6 sports_i[135]
port 406 nsew signal input
rlabel metal3 s 69200 19864 70000 19984 6 sports_i[13]
port 407 nsew signal input
rlabel metal3 s 69200 20136 70000 20256 6 sports_i[14]
port 408 nsew signal input
rlabel metal3 s 69200 20408 70000 20528 6 sports_i[15]
port 409 nsew signal input
rlabel metal3 s 69200 20680 70000 20800 6 sports_i[16]
port 410 nsew signal input
rlabel metal3 s 69200 20952 70000 21072 6 sports_i[17]
port 411 nsew signal input
rlabel metal3 s 69200 21224 70000 21344 6 sports_i[18]
port 412 nsew signal input
rlabel metal3 s 69200 21496 70000 21616 6 sports_i[19]
port 413 nsew signal input
rlabel metal3 s 69200 16600 70000 16720 6 sports_i[1]
port 414 nsew signal input
rlabel metal3 s 69200 21768 70000 21888 6 sports_i[20]
port 415 nsew signal input
rlabel metal3 s 69200 22040 70000 22160 6 sports_i[21]
port 416 nsew signal input
rlabel metal3 s 69200 22312 70000 22432 6 sports_i[22]
port 417 nsew signal input
rlabel metal3 s 69200 22584 70000 22704 6 sports_i[23]
port 418 nsew signal input
rlabel metal3 s 69200 22856 70000 22976 6 sports_i[24]
port 419 nsew signal input
rlabel metal3 s 69200 23128 70000 23248 6 sports_i[25]
port 420 nsew signal input
rlabel metal3 s 69200 23400 70000 23520 6 sports_i[26]
port 421 nsew signal input
rlabel metal3 s 69200 23672 70000 23792 6 sports_i[27]
port 422 nsew signal input
rlabel metal3 s 69200 23944 70000 24064 6 sports_i[28]
port 423 nsew signal input
rlabel metal3 s 69200 24216 70000 24336 6 sports_i[29]
port 424 nsew signal input
rlabel metal3 s 69200 16872 70000 16992 6 sports_i[2]
port 425 nsew signal input
rlabel metal3 s 69200 24488 70000 24608 6 sports_i[30]
port 426 nsew signal input
rlabel metal3 s 69200 24760 70000 24880 6 sports_i[31]
port 427 nsew signal input
rlabel metal3 s 69200 25032 70000 25152 6 sports_i[32]
port 428 nsew signal input
rlabel metal3 s 69200 25304 70000 25424 6 sports_i[33]
port 429 nsew signal input
rlabel metal3 s 69200 25576 70000 25696 6 sports_i[34]
port 430 nsew signal input
rlabel metal3 s 69200 25848 70000 25968 6 sports_i[35]
port 431 nsew signal input
rlabel metal3 s 69200 26120 70000 26240 6 sports_i[36]
port 432 nsew signal input
rlabel metal3 s 69200 26392 70000 26512 6 sports_i[37]
port 433 nsew signal input
rlabel metal3 s 69200 26664 70000 26784 6 sports_i[38]
port 434 nsew signal input
rlabel metal3 s 69200 26936 70000 27056 6 sports_i[39]
port 435 nsew signal input
rlabel metal3 s 69200 17144 70000 17264 6 sports_i[3]
port 436 nsew signal input
rlabel metal3 s 69200 27208 70000 27328 6 sports_i[40]
port 437 nsew signal input
rlabel metal3 s 69200 27480 70000 27600 6 sports_i[41]
port 438 nsew signal input
rlabel metal3 s 69200 27752 70000 27872 6 sports_i[42]
port 439 nsew signal input
rlabel metal3 s 69200 28024 70000 28144 6 sports_i[43]
port 440 nsew signal input
rlabel metal3 s 69200 28296 70000 28416 6 sports_i[44]
port 441 nsew signal input
rlabel metal3 s 69200 28568 70000 28688 6 sports_i[45]
port 442 nsew signal input
rlabel metal3 s 69200 28840 70000 28960 6 sports_i[46]
port 443 nsew signal input
rlabel metal3 s 69200 29112 70000 29232 6 sports_i[47]
port 444 nsew signal input
rlabel metal3 s 69200 29384 70000 29504 6 sports_i[48]
port 445 nsew signal input
rlabel metal3 s 69200 29656 70000 29776 6 sports_i[49]
port 446 nsew signal input
rlabel metal3 s 69200 17416 70000 17536 6 sports_i[4]
port 447 nsew signal input
rlabel metal3 s 69200 29928 70000 30048 6 sports_i[50]
port 448 nsew signal input
rlabel metal3 s 69200 30200 70000 30320 6 sports_i[51]
port 449 nsew signal input
rlabel metal3 s 69200 30472 70000 30592 6 sports_i[52]
port 450 nsew signal input
rlabel metal3 s 69200 30744 70000 30864 6 sports_i[53]
port 451 nsew signal input
rlabel metal3 s 69200 31016 70000 31136 6 sports_i[54]
port 452 nsew signal input
rlabel metal3 s 69200 31288 70000 31408 6 sports_i[55]
port 453 nsew signal input
rlabel metal3 s 69200 31560 70000 31680 6 sports_i[56]
port 454 nsew signal input
rlabel metal3 s 69200 31832 70000 31952 6 sports_i[57]
port 455 nsew signal input
rlabel metal3 s 69200 32104 70000 32224 6 sports_i[58]
port 456 nsew signal input
rlabel metal3 s 69200 32376 70000 32496 6 sports_i[59]
port 457 nsew signal input
rlabel metal3 s 69200 17688 70000 17808 6 sports_i[5]
port 458 nsew signal input
rlabel metal3 s 69200 32648 70000 32768 6 sports_i[60]
port 459 nsew signal input
rlabel metal3 s 69200 32920 70000 33040 6 sports_i[61]
port 460 nsew signal input
rlabel metal3 s 69200 33192 70000 33312 6 sports_i[62]
port 461 nsew signal input
rlabel metal3 s 69200 33464 70000 33584 6 sports_i[63]
port 462 nsew signal input
rlabel metal3 s 69200 33736 70000 33856 6 sports_i[64]
port 463 nsew signal input
rlabel metal3 s 69200 34008 70000 34128 6 sports_i[65]
port 464 nsew signal input
rlabel metal3 s 69200 34280 70000 34400 6 sports_i[66]
port 465 nsew signal input
rlabel metal3 s 69200 34552 70000 34672 6 sports_i[67]
port 466 nsew signal input
rlabel metal3 s 69200 34824 70000 34944 6 sports_i[68]
port 467 nsew signal input
rlabel metal3 s 69200 35096 70000 35216 6 sports_i[69]
port 468 nsew signal input
rlabel metal3 s 69200 17960 70000 18080 6 sports_i[6]
port 469 nsew signal input
rlabel metal3 s 69200 35368 70000 35488 6 sports_i[70]
port 470 nsew signal input
rlabel metal3 s 69200 35640 70000 35760 6 sports_i[71]
port 471 nsew signal input
rlabel metal3 s 69200 35912 70000 36032 6 sports_i[72]
port 472 nsew signal input
rlabel metal3 s 69200 36184 70000 36304 6 sports_i[73]
port 473 nsew signal input
rlabel metal3 s 69200 36456 70000 36576 6 sports_i[74]
port 474 nsew signal input
rlabel metal3 s 69200 36728 70000 36848 6 sports_i[75]
port 475 nsew signal input
rlabel metal3 s 69200 37000 70000 37120 6 sports_i[76]
port 476 nsew signal input
rlabel metal3 s 69200 37272 70000 37392 6 sports_i[77]
port 477 nsew signal input
rlabel metal3 s 69200 37544 70000 37664 6 sports_i[78]
port 478 nsew signal input
rlabel metal3 s 69200 37816 70000 37936 6 sports_i[79]
port 479 nsew signal input
rlabel metal3 s 69200 18232 70000 18352 6 sports_i[7]
port 480 nsew signal input
rlabel metal3 s 69200 38088 70000 38208 6 sports_i[80]
port 481 nsew signal input
rlabel metal3 s 69200 38360 70000 38480 6 sports_i[81]
port 482 nsew signal input
rlabel metal3 s 69200 38632 70000 38752 6 sports_i[82]
port 483 nsew signal input
rlabel metal3 s 69200 38904 70000 39024 6 sports_i[83]
port 484 nsew signal input
rlabel metal3 s 69200 39176 70000 39296 6 sports_i[84]
port 485 nsew signal input
rlabel metal3 s 69200 39448 70000 39568 6 sports_i[85]
port 486 nsew signal input
rlabel metal3 s 69200 39720 70000 39840 6 sports_i[86]
port 487 nsew signal input
rlabel metal3 s 69200 39992 70000 40112 6 sports_i[87]
port 488 nsew signal input
rlabel metal3 s 69200 40264 70000 40384 6 sports_i[88]
port 489 nsew signal input
rlabel metal3 s 69200 40536 70000 40656 6 sports_i[89]
port 490 nsew signal input
rlabel metal3 s 69200 18504 70000 18624 6 sports_i[8]
port 491 nsew signal input
rlabel metal3 s 69200 40808 70000 40928 6 sports_i[90]
port 492 nsew signal input
rlabel metal3 s 69200 41080 70000 41200 6 sports_i[91]
port 493 nsew signal input
rlabel metal3 s 69200 41352 70000 41472 6 sports_i[92]
port 494 nsew signal input
rlabel metal3 s 69200 41624 70000 41744 6 sports_i[93]
port 495 nsew signal input
rlabel metal3 s 69200 41896 70000 42016 6 sports_i[94]
port 496 nsew signal input
rlabel metal3 s 69200 42168 70000 42288 6 sports_i[95]
port 497 nsew signal input
rlabel metal3 s 69200 42440 70000 42560 6 sports_i[96]
port 498 nsew signal input
rlabel metal3 s 69200 42712 70000 42832 6 sports_i[97]
port 499 nsew signal input
rlabel metal3 s 69200 42984 70000 43104 6 sports_i[98]
port 500 nsew signal input
rlabel metal3 s 69200 43256 70000 43376 6 sports_i[99]
port 501 nsew signal input
rlabel metal3 s 69200 18776 70000 18896 6 sports_i[9]
port 502 nsew signal input
rlabel metal3 s 0 3816 800 3936 6 sports_o[0]
port 503 nsew signal output
rlabel metal3 s 0 31016 800 31136 6 sports_o[100]
port 504 nsew signal output
rlabel metal3 s 0 31288 800 31408 6 sports_o[101]
port 505 nsew signal output
rlabel metal3 s 0 31560 800 31680 6 sports_o[102]
port 506 nsew signal output
rlabel metal3 s 0 31832 800 31952 6 sports_o[103]
port 507 nsew signal output
rlabel metal3 s 0 32104 800 32224 6 sports_o[104]
port 508 nsew signal output
rlabel metal3 s 0 32376 800 32496 6 sports_o[105]
port 509 nsew signal output
rlabel metal3 s 0 32648 800 32768 6 sports_o[106]
port 510 nsew signal output
rlabel metal3 s 0 32920 800 33040 6 sports_o[107]
port 511 nsew signal output
rlabel metal3 s 0 33192 800 33312 6 sports_o[108]
port 512 nsew signal output
rlabel metal3 s 0 33464 800 33584 6 sports_o[109]
port 513 nsew signal output
rlabel metal3 s 0 6536 800 6656 6 sports_o[10]
port 514 nsew signal output
rlabel metal3 s 0 33736 800 33856 6 sports_o[110]
port 515 nsew signal output
rlabel metal3 s 0 34008 800 34128 6 sports_o[111]
port 516 nsew signal output
rlabel metal3 s 0 34280 800 34400 6 sports_o[112]
port 517 nsew signal output
rlabel metal3 s 0 34552 800 34672 6 sports_o[113]
port 518 nsew signal output
rlabel metal3 s 0 34824 800 34944 6 sports_o[114]
port 519 nsew signal output
rlabel metal3 s 0 35096 800 35216 6 sports_o[115]
port 520 nsew signal output
rlabel metal3 s 0 35368 800 35488 6 sports_o[116]
port 521 nsew signal output
rlabel metal3 s 0 35640 800 35760 6 sports_o[117]
port 522 nsew signal output
rlabel metal3 s 0 35912 800 36032 6 sports_o[118]
port 523 nsew signal output
rlabel metal3 s 0 36184 800 36304 6 sports_o[119]
port 524 nsew signal output
rlabel metal3 s 0 6808 800 6928 6 sports_o[11]
port 525 nsew signal output
rlabel metal3 s 0 36456 800 36576 6 sports_o[120]
port 526 nsew signal output
rlabel metal3 s 0 36728 800 36848 6 sports_o[121]
port 527 nsew signal output
rlabel metal3 s 0 37000 800 37120 6 sports_o[122]
port 528 nsew signal output
rlabel metal3 s 0 37272 800 37392 6 sports_o[123]
port 529 nsew signal output
rlabel metal3 s 0 37544 800 37664 6 sports_o[124]
port 530 nsew signal output
rlabel metal3 s 0 37816 800 37936 6 sports_o[125]
port 531 nsew signal output
rlabel metal3 s 0 38088 800 38208 6 sports_o[126]
port 532 nsew signal output
rlabel metal3 s 0 38360 800 38480 6 sports_o[127]
port 533 nsew signal output
rlabel metal3 s 0 38632 800 38752 6 sports_o[128]
port 534 nsew signal output
rlabel metal3 s 0 38904 800 39024 6 sports_o[129]
port 535 nsew signal output
rlabel metal3 s 0 7080 800 7200 6 sports_o[12]
port 536 nsew signal output
rlabel metal3 s 0 39176 800 39296 6 sports_o[130]
port 537 nsew signal output
rlabel metal3 s 0 39448 800 39568 6 sports_o[131]
port 538 nsew signal output
rlabel metal3 s 0 39720 800 39840 6 sports_o[132]
port 539 nsew signal output
rlabel metal3 s 0 39992 800 40112 6 sports_o[133]
port 540 nsew signal output
rlabel metal3 s 0 40264 800 40384 6 sports_o[134]
port 541 nsew signal output
rlabel metal3 s 0 40536 800 40656 6 sports_o[135]
port 542 nsew signal output
rlabel metal3 s 0 40808 800 40928 6 sports_o[136]
port 543 nsew signal output
rlabel metal3 s 0 41080 800 41200 6 sports_o[137]
port 544 nsew signal output
rlabel metal3 s 0 41352 800 41472 6 sports_o[138]
port 545 nsew signal output
rlabel metal3 s 0 41624 800 41744 6 sports_o[139]
port 546 nsew signal output
rlabel metal3 s 0 7352 800 7472 6 sports_o[13]
port 547 nsew signal output
rlabel metal3 s 0 41896 800 42016 6 sports_o[140]
port 548 nsew signal output
rlabel metal3 s 0 42168 800 42288 6 sports_o[141]
port 549 nsew signal output
rlabel metal3 s 0 42440 800 42560 6 sports_o[142]
port 550 nsew signal output
rlabel metal3 s 0 42712 800 42832 6 sports_o[143]
port 551 nsew signal output
rlabel metal3 s 0 42984 800 43104 6 sports_o[144]
port 552 nsew signal output
rlabel metal3 s 0 43256 800 43376 6 sports_o[145]
port 553 nsew signal output
rlabel metal3 s 0 43528 800 43648 6 sports_o[146]
port 554 nsew signal output
rlabel metal3 s 0 43800 800 43920 6 sports_o[147]
port 555 nsew signal output
rlabel metal3 s 0 44072 800 44192 6 sports_o[148]
port 556 nsew signal output
rlabel metal3 s 0 44344 800 44464 6 sports_o[149]
port 557 nsew signal output
rlabel metal3 s 0 7624 800 7744 6 sports_o[14]
port 558 nsew signal output
rlabel metal3 s 0 44616 800 44736 6 sports_o[150]
port 559 nsew signal output
rlabel metal3 s 0 44888 800 45008 6 sports_o[151]
port 560 nsew signal output
rlabel metal3 s 0 45160 800 45280 6 sports_o[152]
port 561 nsew signal output
rlabel metal3 s 0 45432 800 45552 6 sports_o[153]
port 562 nsew signal output
rlabel metal3 s 0 45704 800 45824 6 sports_o[154]
port 563 nsew signal output
rlabel metal3 s 0 45976 800 46096 6 sports_o[155]
port 564 nsew signal output
rlabel metal3 s 0 46248 800 46368 6 sports_o[156]
port 565 nsew signal output
rlabel metal3 s 0 46520 800 46640 6 sports_o[157]
port 566 nsew signal output
rlabel metal3 s 0 46792 800 46912 6 sports_o[158]
port 567 nsew signal output
rlabel metal3 s 0 47064 800 47184 6 sports_o[159]
port 568 nsew signal output
rlabel metal3 s 0 7896 800 8016 6 sports_o[15]
port 569 nsew signal output
rlabel metal3 s 0 47336 800 47456 6 sports_o[160]
port 570 nsew signal output
rlabel metal3 s 0 47608 800 47728 6 sports_o[161]
port 571 nsew signal output
rlabel metal3 s 0 47880 800 48000 6 sports_o[162]
port 572 nsew signal output
rlabel metal3 s 0 48152 800 48272 6 sports_o[163]
port 573 nsew signal output
rlabel metal3 s 0 48424 800 48544 6 sports_o[164]
port 574 nsew signal output
rlabel metal3 s 0 48696 800 48816 6 sports_o[165]
port 575 nsew signal output
rlabel metal3 s 0 48968 800 49088 6 sports_o[166]
port 576 nsew signal output
rlabel metal3 s 0 49240 800 49360 6 sports_o[167]
port 577 nsew signal output
rlabel metal3 s 0 49512 800 49632 6 sports_o[168]
port 578 nsew signal output
rlabel metal3 s 0 49784 800 49904 6 sports_o[169]
port 579 nsew signal output
rlabel metal3 s 0 8168 800 8288 6 sports_o[16]
port 580 nsew signal output
rlabel metal3 s 0 50056 800 50176 6 sports_o[170]
port 581 nsew signal output
rlabel metal3 s 0 50328 800 50448 6 sports_o[171]
port 582 nsew signal output
rlabel metal3 s 0 50600 800 50720 6 sports_o[172]
port 583 nsew signal output
rlabel metal3 s 0 50872 800 50992 6 sports_o[173]
port 584 nsew signal output
rlabel metal3 s 0 51144 800 51264 6 sports_o[174]
port 585 nsew signal output
rlabel metal3 s 0 51416 800 51536 6 sports_o[175]
port 586 nsew signal output
rlabel metal3 s 0 51688 800 51808 6 sports_o[176]
port 587 nsew signal output
rlabel metal3 s 0 51960 800 52080 6 sports_o[177]
port 588 nsew signal output
rlabel metal3 s 0 52232 800 52352 6 sports_o[178]
port 589 nsew signal output
rlabel metal3 s 0 52504 800 52624 6 sports_o[179]
port 590 nsew signal output
rlabel metal3 s 0 8440 800 8560 6 sports_o[17]
port 591 nsew signal output
rlabel metal3 s 0 52776 800 52896 6 sports_o[180]
port 592 nsew signal output
rlabel metal3 s 0 53048 800 53168 6 sports_o[181]
port 593 nsew signal output
rlabel metal3 s 0 53320 800 53440 6 sports_o[182]
port 594 nsew signal output
rlabel metal3 s 0 53592 800 53712 6 sports_o[183]
port 595 nsew signal output
rlabel metal3 s 0 53864 800 53984 6 sports_o[184]
port 596 nsew signal output
rlabel metal3 s 0 54136 800 54256 6 sports_o[185]
port 597 nsew signal output
rlabel metal3 s 0 54408 800 54528 6 sports_o[186]
port 598 nsew signal output
rlabel metal3 s 0 54680 800 54800 6 sports_o[187]
port 599 nsew signal output
rlabel metal3 s 0 54952 800 55072 6 sports_o[188]
port 600 nsew signal output
rlabel metal3 s 0 55224 800 55344 6 sports_o[189]
port 601 nsew signal output
rlabel metal3 s 0 8712 800 8832 6 sports_o[18]
port 602 nsew signal output
rlabel metal3 s 0 55496 800 55616 6 sports_o[190]
port 603 nsew signal output
rlabel metal3 s 0 55768 800 55888 6 sports_o[191]
port 604 nsew signal output
rlabel metal3 s 0 56040 800 56160 6 sports_o[192]
port 605 nsew signal output
rlabel metal3 s 0 56312 800 56432 6 sports_o[193]
port 606 nsew signal output
rlabel metal3 s 0 56584 800 56704 6 sports_o[194]
port 607 nsew signal output
rlabel metal3 s 0 56856 800 56976 6 sports_o[195]
port 608 nsew signal output
rlabel metal3 s 0 57128 800 57248 6 sports_o[196]
port 609 nsew signal output
rlabel metal3 s 0 57400 800 57520 6 sports_o[197]
port 610 nsew signal output
rlabel metal3 s 0 57672 800 57792 6 sports_o[198]
port 611 nsew signal output
rlabel metal3 s 0 57944 800 58064 6 sports_o[199]
port 612 nsew signal output
rlabel metal3 s 0 8984 800 9104 6 sports_o[19]
port 613 nsew signal output
rlabel metal3 s 0 4088 800 4208 6 sports_o[1]
port 614 nsew signal output
rlabel metal3 s 0 58216 800 58336 6 sports_o[200]
port 615 nsew signal output
rlabel metal3 s 0 58488 800 58608 6 sports_o[201]
port 616 nsew signal output
rlabel metal3 s 0 58760 800 58880 6 sports_o[202]
port 617 nsew signal output
rlabel metal3 s 0 59032 800 59152 6 sports_o[203]
port 618 nsew signal output
rlabel metal3 s 0 59304 800 59424 6 sports_o[204]
port 619 nsew signal output
rlabel metal3 s 0 59576 800 59696 6 sports_o[205]
port 620 nsew signal output
rlabel metal3 s 0 59848 800 59968 6 sports_o[206]
port 621 nsew signal output
rlabel metal3 s 0 60120 800 60240 6 sports_o[207]
port 622 nsew signal output
rlabel metal3 s 0 60392 800 60512 6 sports_o[208]
port 623 nsew signal output
rlabel metal3 s 0 60664 800 60784 6 sports_o[209]
port 624 nsew signal output
rlabel metal3 s 0 9256 800 9376 6 sports_o[20]
port 625 nsew signal output
rlabel metal3 s 0 60936 800 61056 6 sports_o[210]
port 626 nsew signal output
rlabel metal3 s 0 61208 800 61328 6 sports_o[211]
port 627 nsew signal output
rlabel metal3 s 0 61480 800 61600 6 sports_o[212]
port 628 nsew signal output
rlabel metal3 s 0 61752 800 61872 6 sports_o[213]
port 629 nsew signal output
rlabel metal3 s 0 62024 800 62144 6 sports_o[214]
port 630 nsew signal output
rlabel metal3 s 0 62296 800 62416 6 sports_o[215]
port 631 nsew signal output
rlabel metal3 s 0 62568 800 62688 6 sports_o[216]
port 632 nsew signal output
rlabel metal3 s 0 62840 800 62960 6 sports_o[217]
port 633 nsew signal output
rlabel metal3 s 0 63112 800 63232 6 sports_o[218]
port 634 nsew signal output
rlabel metal3 s 0 63384 800 63504 6 sports_o[219]
port 635 nsew signal output
rlabel metal3 s 0 9528 800 9648 6 sports_o[21]
port 636 nsew signal output
rlabel metal3 s 0 63656 800 63776 6 sports_o[220]
port 637 nsew signal output
rlabel metal3 s 0 63928 800 64048 6 sports_o[221]
port 638 nsew signal output
rlabel metal3 s 0 64200 800 64320 6 sports_o[222]
port 639 nsew signal output
rlabel metal3 s 0 64472 800 64592 6 sports_o[223]
port 640 nsew signal output
rlabel metal3 s 0 64744 800 64864 6 sports_o[224]
port 641 nsew signal output
rlabel metal3 s 0 65016 800 65136 6 sports_o[225]
port 642 nsew signal output
rlabel metal3 s 0 65288 800 65408 6 sports_o[226]
port 643 nsew signal output
rlabel metal3 s 0 65560 800 65680 6 sports_o[227]
port 644 nsew signal output
rlabel metal3 s 0 9800 800 9920 6 sports_o[22]
port 645 nsew signal output
rlabel metal3 s 0 10072 800 10192 6 sports_o[23]
port 646 nsew signal output
rlabel metal3 s 0 10344 800 10464 6 sports_o[24]
port 647 nsew signal output
rlabel metal3 s 0 10616 800 10736 6 sports_o[25]
port 648 nsew signal output
rlabel metal3 s 0 10888 800 11008 6 sports_o[26]
port 649 nsew signal output
rlabel metal3 s 0 11160 800 11280 6 sports_o[27]
port 650 nsew signal output
rlabel metal3 s 0 11432 800 11552 6 sports_o[28]
port 651 nsew signal output
rlabel metal3 s 0 11704 800 11824 6 sports_o[29]
port 652 nsew signal output
rlabel metal3 s 0 4360 800 4480 6 sports_o[2]
port 653 nsew signal output
rlabel metal3 s 0 11976 800 12096 6 sports_o[30]
port 654 nsew signal output
rlabel metal3 s 0 12248 800 12368 6 sports_o[31]
port 655 nsew signal output
rlabel metal3 s 0 12520 800 12640 6 sports_o[32]
port 656 nsew signal output
rlabel metal3 s 0 12792 800 12912 6 sports_o[33]
port 657 nsew signal output
rlabel metal3 s 0 13064 800 13184 6 sports_o[34]
port 658 nsew signal output
rlabel metal3 s 0 13336 800 13456 6 sports_o[35]
port 659 nsew signal output
rlabel metal3 s 0 13608 800 13728 6 sports_o[36]
port 660 nsew signal output
rlabel metal3 s 0 13880 800 14000 6 sports_o[37]
port 661 nsew signal output
rlabel metal3 s 0 14152 800 14272 6 sports_o[38]
port 662 nsew signal output
rlabel metal3 s 0 14424 800 14544 6 sports_o[39]
port 663 nsew signal output
rlabel metal3 s 0 4632 800 4752 6 sports_o[3]
port 664 nsew signal output
rlabel metal3 s 0 14696 800 14816 6 sports_o[40]
port 665 nsew signal output
rlabel metal3 s 0 14968 800 15088 6 sports_o[41]
port 666 nsew signal output
rlabel metal3 s 0 15240 800 15360 6 sports_o[42]
port 667 nsew signal output
rlabel metal3 s 0 15512 800 15632 6 sports_o[43]
port 668 nsew signal output
rlabel metal3 s 0 15784 800 15904 6 sports_o[44]
port 669 nsew signal output
rlabel metal3 s 0 16056 800 16176 6 sports_o[45]
port 670 nsew signal output
rlabel metal3 s 0 16328 800 16448 6 sports_o[46]
port 671 nsew signal output
rlabel metal3 s 0 16600 800 16720 6 sports_o[47]
port 672 nsew signal output
rlabel metal3 s 0 16872 800 16992 6 sports_o[48]
port 673 nsew signal output
rlabel metal3 s 0 17144 800 17264 6 sports_o[49]
port 674 nsew signal output
rlabel metal3 s 0 4904 800 5024 6 sports_o[4]
port 675 nsew signal output
rlabel metal3 s 0 17416 800 17536 6 sports_o[50]
port 676 nsew signal output
rlabel metal3 s 0 17688 800 17808 6 sports_o[51]
port 677 nsew signal output
rlabel metal3 s 0 17960 800 18080 6 sports_o[52]
port 678 nsew signal output
rlabel metal3 s 0 18232 800 18352 6 sports_o[53]
port 679 nsew signal output
rlabel metal3 s 0 18504 800 18624 6 sports_o[54]
port 680 nsew signal output
rlabel metal3 s 0 18776 800 18896 6 sports_o[55]
port 681 nsew signal output
rlabel metal3 s 0 19048 800 19168 6 sports_o[56]
port 682 nsew signal output
rlabel metal3 s 0 19320 800 19440 6 sports_o[57]
port 683 nsew signal output
rlabel metal3 s 0 19592 800 19712 6 sports_o[58]
port 684 nsew signal output
rlabel metal3 s 0 19864 800 19984 6 sports_o[59]
port 685 nsew signal output
rlabel metal3 s 0 5176 800 5296 6 sports_o[5]
port 686 nsew signal output
rlabel metal3 s 0 20136 800 20256 6 sports_o[60]
port 687 nsew signal output
rlabel metal3 s 0 20408 800 20528 6 sports_o[61]
port 688 nsew signal output
rlabel metal3 s 0 20680 800 20800 6 sports_o[62]
port 689 nsew signal output
rlabel metal3 s 0 20952 800 21072 6 sports_o[63]
port 690 nsew signal output
rlabel metal3 s 0 21224 800 21344 6 sports_o[64]
port 691 nsew signal output
rlabel metal3 s 0 21496 800 21616 6 sports_o[65]
port 692 nsew signal output
rlabel metal3 s 0 21768 800 21888 6 sports_o[66]
port 693 nsew signal output
rlabel metal3 s 0 22040 800 22160 6 sports_o[67]
port 694 nsew signal output
rlabel metal3 s 0 22312 800 22432 6 sports_o[68]
port 695 nsew signal output
rlabel metal3 s 0 22584 800 22704 6 sports_o[69]
port 696 nsew signal output
rlabel metal3 s 0 5448 800 5568 6 sports_o[6]
port 697 nsew signal output
rlabel metal3 s 0 22856 800 22976 6 sports_o[70]
port 698 nsew signal output
rlabel metal3 s 0 23128 800 23248 6 sports_o[71]
port 699 nsew signal output
rlabel metal3 s 0 23400 800 23520 6 sports_o[72]
port 700 nsew signal output
rlabel metal3 s 0 23672 800 23792 6 sports_o[73]
port 701 nsew signal output
rlabel metal3 s 0 23944 800 24064 6 sports_o[74]
port 702 nsew signal output
rlabel metal3 s 0 24216 800 24336 6 sports_o[75]
port 703 nsew signal output
rlabel metal3 s 0 24488 800 24608 6 sports_o[76]
port 704 nsew signal output
rlabel metal3 s 0 24760 800 24880 6 sports_o[77]
port 705 nsew signal output
rlabel metal3 s 0 25032 800 25152 6 sports_o[78]
port 706 nsew signal output
rlabel metal3 s 0 25304 800 25424 6 sports_o[79]
port 707 nsew signal output
rlabel metal3 s 0 5720 800 5840 6 sports_o[7]
port 708 nsew signal output
rlabel metal3 s 0 25576 800 25696 6 sports_o[80]
port 709 nsew signal output
rlabel metal3 s 0 25848 800 25968 6 sports_o[81]
port 710 nsew signal output
rlabel metal3 s 0 26120 800 26240 6 sports_o[82]
port 711 nsew signal output
rlabel metal3 s 0 26392 800 26512 6 sports_o[83]
port 712 nsew signal output
rlabel metal3 s 0 26664 800 26784 6 sports_o[84]
port 713 nsew signal output
rlabel metal3 s 0 26936 800 27056 6 sports_o[85]
port 714 nsew signal output
rlabel metal3 s 0 27208 800 27328 6 sports_o[86]
port 715 nsew signal output
rlabel metal3 s 0 27480 800 27600 6 sports_o[87]
port 716 nsew signal output
rlabel metal3 s 0 27752 800 27872 6 sports_o[88]
port 717 nsew signal output
rlabel metal3 s 0 28024 800 28144 6 sports_o[89]
port 718 nsew signal output
rlabel metal3 s 0 5992 800 6112 6 sports_o[8]
port 719 nsew signal output
rlabel metal3 s 0 28296 800 28416 6 sports_o[90]
port 720 nsew signal output
rlabel metal3 s 0 28568 800 28688 6 sports_o[91]
port 721 nsew signal output
rlabel metal3 s 0 28840 800 28960 6 sports_o[92]
port 722 nsew signal output
rlabel metal3 s 0 29112 800 29232 6 sports_o[93]
port 723 nsew signal output
rlabel metal3 s 0 29384 800 29504 6 sports_o[94]
port 724 nsew signal output
rlabel metal3 s 0 29656 800 29776 6 sports_o[95]
port 725 nsew signal output
rlabel metal3 s 0 29928 800 30048 6 sports_o[96]
port 726 nsew signal output
rlabel metal3 s 0 30200 800 30320 6 sports_o[97]
port 727 nsew signal output
rlabel metal3 s 0 30472 800 30592 6 sports_o[98]
port 728 nsew signal output
rlabel metal3 s 0 30744 800 30864 6 sports_o[99]
port 729 nsew signal output
rlabel metal3 s 0 6264 800 6384 6 sports_o[9]
port 730 nsew signal output
rlabel metal4 s 4208 2128 4528 67504 6 vccd1
port 731 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 67504 6 vccd1
port 731 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 67504 6 vccd1
port 731 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 67504 6 vssd1
port 732 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 67504 6 vssd1
port 732 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 70000 70000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 8067562
string GDS_FILE /local/colinm22/sdmay26-24/openlane/busarb_2_2/runs/25_10_02_14_45/results/signoff/busarb_2_2.magic.gds
string GDS_START 543220
<< end >>

