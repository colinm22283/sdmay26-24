// This is the unpowered netlist.
module mac_piped (clk,
    nrst,
    a_i,
    b_i,
    y_o);
 input clk;
 input nrst;
 input [31:0] a_i;
 input [31:0] b_i;
 output [31:0] y_o;

 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire \ab[0] ;
 wire \ab[10] ;
 wire \ab[11] ;
 wire \ab[12] ;
 wire \ab[13] ;
 wire \ab[14] ;
 wire \ab[15] ;
 wire \ab[16] ;
 wire \ab[17] ;
 wire \ab[18] ;
 wire \ab[19] ;
 wire \ab[1] ;
 wire \ab[20] ;
 wire \ab[21] ;
 wire \ab[2] ;
 wire \ab[3] ;
 wire \ab[4] ;
 wire \ab[5] ;
 wire \ab[6] ;
 wire \ab[7] ;
 wire \ab[8] ;
 wire \ab[9] ;
 wire \abprod[0] ;
 wire \abprod[10] ;
 wire \abprod[11] ;
 wire \abprod[12] ;
 wire \abprod[13] ;
 wire \abprod[14] ;
 wire \abprod[15] ;
 wire \abprod[16] ;
 wire \abprod[17] ;
 wire \abprod[18] ;
 wire \abprod[19] ;
 wire \abprod[1] ;
 wire \abprod[20] ;
 wire \abprod[21] ;
 wire \abprod[2] ;
 wire \abprod[3] ;
 wire \abprod[4] ;
 wire \abprod[5] ;
 wire \abprod[6] ;
 wire \abprod[7] ;
 wire \abprod[8] ;
 wire \abprod[9] ;
 wire \absum[0] ;
 wire \absum[10] ;
 wire \absum[11] ;
 wire \absum[12] ;
 wire \absum[13] ;
 wire \absum[14] ;
 wire \absum[15] ;
 wire \absum[16] ;
 wire \absum[17] ;
 wire \absum[18] ;
 wire \absum[19] ;
 wire \absum[1] ;
 wire \absum[20] ;
 wire \absum[21] ;
 wire \absum[22] ;
 wire \absum[23] ;
 wire \absum[24] ;
 wire \absum[25] ;
 wire \absum[26] ;
 wire \absum[27] ;
 wire \absum[28] ;
 wire \absum[29] ;
 wire \absum[2] ;
 wire \absum[30] ;
 wire \absum[31] ;
 wire \absum[3] ;
 wire \absum[4] ;
 wire \absum[5] ;
 wire \absum[6] ;
 wire \absum[7] ;
 wire \absum[8] ;
 wire \absum[9] ;
 wire clknet_0_clk;
 wire clknet_2_0__leaf_clk;
 wire clknet_2_1__leaf_clk;
 wire clknet_2_2__leaf_clk;
 wire clknet_2_3__leaf_clk;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net15;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net16;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net17;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net18;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net19;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net2;
 wire net20;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net21;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net22;
 wire net220;
 wire net221;
 wire net222;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net3;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net4;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net5;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net6;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net7;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net8;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;

 sky130_fd_sc_hd__diode_2 ANTENNA__05203__A (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA__05204__A (.DIODE(_00740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05204__B (.DIODE(_00751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05207__A (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA__05208__A (.DIODE(_00784_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05208__B (.DIODE(_00795_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05213__A (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__05214__A (.DIODE(_00850_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05214__B (.DIODE(_00861_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05221__A (.DIODE(_00850_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05221__B (.DIODE(_00751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05222__A (.DIODE(_00740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05222__B (.DIODE(_00795_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05224__A (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__05224__B (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__05231__A (.DIODE(_01037_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05231__B (.DIODE(_01048_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05233__A (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__05235__A (.DIODE(_01081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05235__B (.DIODE(_01092_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05239__A (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__05241__A (.DIODE(_01147_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05241__B (.DIODE(_01158_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05253__A (.DIODE(_00784_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05253__B (.DIODE(_00751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05256__A (.DIODE(_01323_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05256__B (.DIODE(_00795_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05259__A (.DIODE(_00740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05259__B (.DIODE(_00861_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05270__A (.DIODE(_01081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05270__B (.DIODE(_01048_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05272__A (.DIODE(_00850_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05272__B (.DIODE(_01092_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05277__A (.DIODE(_01158_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05278__A (.DIODE(_01037_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05278__B (.DIODE(_01565_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05297__A (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__05297__B (.DIODE(_01774_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05300__A (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__05300__B (.DIODE(_01807_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05305__A (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__05307__A (.DIODE(_01873_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05307__B (.DIODE(_01884_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05316__A (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__05316__B (.DIODE(_01807_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05318__A (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__05318__B (.DIODE(_01774_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05321__A (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA__05322__A (.DIODE(_02049_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05322__B (.DIODE(_01884_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05349__A (.DIODE(_00751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05350__A (.DIODE(_01081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05350__B (.DIODE(_02357_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05351__A (.DIODE(_00795_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05352__A (.DIODE(_00850_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05352__B (.DIODE(_02379_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05354__A (.DIODE(_01037_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05354__B (.DIODE(_00861_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05359__A (.DIODE(_01147_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05359__B (.DIODE(_01048_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05361__B (.DIODE(_01092_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05366__A (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__05367__A (.DIODE(_02544_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05367__B (.DIODE(_01158_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05386__A (.DIODE(_02753_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05386__B (.DIODE(_01884_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05387__A (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA__05387__B (.DIODE(_01774_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05389__A (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__05389__B (.DIODE(_01807_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05408__A (.DIODE(_02753_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05408__B (.DIODE(_02995_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05411__A (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA__05411__B (.DIODE(_03028_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05417__A (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__05417__B (.DIODE(_03094_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05422__A (.DIODE(_02753_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05423__A (.DIODE(_03160_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05423__B (.DIODE(_03028_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05424__A (.DIODE(_03094_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05425__A (.DIODE(_03182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05425__B (.DIODE(_02995_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05427__A (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__05429__A (.DIODE(_03215_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05429__B (.DIODE(_03226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05437__A (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__05437__B (.DIODE(_03314_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05439__A (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__05439__B (.DIODE(_03226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05445__A (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__05445__B (.DIODE(_03402_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05466__A (.DIODE(_03226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05466__B (.DIODE(_02995_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05467__A (.DIODE(_03094_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05467__B (.DIODE(_03028_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05469__A (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__05469__B (.DIODE(_03314_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05476__A (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__05476__B (.DIODE(_03402_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05477__A (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__05477__B (.DIODE(_03314_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05481__A (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__05483__A (.DIODE(_03809_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05483__B (.DIODE(_03820_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05507__A (.DIODE(_02379_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05507__B (.DIODE(_04084_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05509__A (.DIODE(_01323_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05509__B (.DIODE(_00751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05512__A (.DIODE(_00784_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05512__B (.DIODE(_00861_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05522__A (.DIODE(_01048_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05523__A (.DIODE(_00850_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05523__B (.DIODE(_04260_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05525__A (.DIODE(_01092_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05526__A (.DIODE(_00740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05526__B (.DIODE(_04293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05531__A (.DIODE(_01081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05531__B (.DIODE(_01158_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05542__A (.DIODE(_01147_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05542__B (.DIODE(_01774_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05544__B (.DIODE(_01807_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05549__A (.DIODE(_02544_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05549__B (.DIODE(_01884_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05578__A (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA__05578__B (.DIODE(_02995_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05580__A (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__05580__B (.DIODE(_03028_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05585__A (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__05585__B (.DIODE(_02753_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05595__A (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__05595__B (.DIODE(_03226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05597__A (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__05597__B (.DIODE(_03094_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05602__A (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__05602__B (.DIODE(_03314_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05635__A (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__05637__A (.DIODE(_04808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05637__B (.DIODE(_04809_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05639__A (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__05640__A (.DIODE(_04812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05640__B (.DIODE(_03820_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05647__A (.DIODE(_04818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05647__B (.DIODE(_04819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05654__A (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__05655__A (.DIODE(_04827_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05656__A (.DIODE(_04818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05656__B (.DIODE(_04828_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05657__A (.DIODE(_04812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05657__B (.DIODE(_04809_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05659__A (.DIODE(_04808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05659__B (.DIODE(_04819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05667__A (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__05667__B (.DIODE(_03820_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05669__A (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__05669__B (.DIODE(_03402_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05674__A (.DIODE(_04818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05674__B (.DIODE(_04809_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05698__A (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__05699__A (.DIODE(_04871_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05699__B (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__05701__A (.DIODE(_04873_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05701__B (.DIODE(_04827_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05704__A (.DIODE(_04876_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05704__B (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05708__A (.DIODE(_04871_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05708__B (.DIODE(_04827_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05709__A (.DIODE(_04873_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05709__B (.DIODE(_04819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05714__A (.DIODE(_04876_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05714__B (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__05722__A (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05723__A (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__05723__B (.DIODE(_04895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05738__A (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__05739__A (.DIODE(_04873_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05739__B (.DIODE(_04871_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05739__C (.DIODE(_04911_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05739__D (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__05754__A (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__05754__B (.DIODE(_03820_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05755__A (.DIODE(_03402_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05756__A (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__05756__B (.DIODE(_04928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05758__A (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__05758__B (.DIODE(_04809_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05763__A (.DIODE(_04808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05763__B (.DIODE(_04827_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05764__A (.DIODE(_04812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05764__B (.DIODE(_04819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05768__A (.DIODE(_04818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05768__B (.DIODE(_04911_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05789__A (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__05790__A (.DIODE(_04962_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05790__B (.DIODE(_04809_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05791__A (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__05792__A (.DIODE(_04964_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05792__B (.DIODE(_03820_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05794__A (.DIODE(_03809_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05794__B (.DIODE(_04819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05799__A (.DIODE(_04818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05799__B (.DIODE(_04895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05800__A (.DIODE(_04808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05800__B (.DIODE(_04911_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05802__A (.DIODE(_04812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05802__B (.DIODE(_04827_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05818__A (.DIODE(_04911_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05819__A (.DIODE(_04895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05820__A1 (.DIODE(_04873_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05820__A2 (.DIODE(_04991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05820__B1 (.DIODE(_04871_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05820__B2 (.DIODE(_04992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05832__A (.DIODE(_01873_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05832__B (.DIODE(_01565_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05834__A (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__05834__B (.DIODE(_01048_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05835__A (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__05835__B (.DIODE(_01092_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05842__A (.DIODE(_02753_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05842__B (.DIODE(_01774_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05844__A (.DIODE(_02049_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05844__B (.DIODE(_01807_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05847__A (.DIODE(_03182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05847__B (.DIODE(_01884_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05855__A (.DIODE(_03314_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05856__A (.DIODE(_02995_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05857__A (.DIODE(_05028_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05857__B (.DIODE(_05029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05858__A (.DIODE(_03226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05859__A (.DIODE(_03028_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05860__A (.DIODE(_05031_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05860__B (.DIODE(_05032_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05862__A (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__05862__B (.DIODE(_04928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05939__A (.DIODE(_01037_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05939__B (.DIODE(_02357_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05940__A (.DIODE(_01081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05940__B (.DIODE(_02379_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05942__A (.DIODE(_01147_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05942__B (.DIODE(_00861_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05985__A (.DIODE(_00751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05985__B (.DIODE(_04084_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05988__A (.DIODE(_00795_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05988__B (.DIODE(_05160_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05993__A (.DIODE(_01323_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05993__B (.DIODE(_00861_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06003__A (.DIODE(_00740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06003__B (.DIODE(_01048_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06005__A (.DIODE(_00784_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06005__B (.DIODE(_01092_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06010__A (.DIODE(_00850_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06010__B (.DIODE(_01158_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06025__A (.DIODE(_01037_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06025__B (.DIODE(_01774_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06027__A (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__06027__B (.DIODE(_01807_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06032__A (.DIODE(_01884_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06033__A (.DIODE(_01147_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06033__B (.DIODE(_00003_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06054__A (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__06054__B (.DIODE(_03094_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06055__A (.DIODE(_04964_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06055__B (.DIODE(_03160_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06060__A (.DIODE(_03809_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06060__B (.DIODE(_03226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06068__A (.DIODE(_01873_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06068__B (.DIODE(_02995_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06070__A (.DIODE(_02544_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06070__B (.DIODE(_03028_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06073__A (.DIODE(_03215_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06073__B (.DIODE(_02049_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06109__A (.DIODE(_04808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06109__B (.DIODE(_03402_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06111__A (.DIODE(_04812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06111__B (.DIODE(_03314_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06116__A (.DIODE(_04818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06116__B (.DIODE(_03820_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06137__A (.DIODE(_04871_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06137__B (.DIODE(_04819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06138__B (.DIODE(_04873_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06138__C (.DIODE(_04809_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06139__A (.DIODE(_04873_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06140__A (.DIODE(_04809_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06143__A (.DIODE(_04876_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06143__B (.DIODE(_04827_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06154__A (.DIODE(_00124_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06154__B (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06155__A (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__06155__B (.DIODE(_04911_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06171__A (.DIODE(_00141_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06173__A (.DIODE(_00141_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06225__A (.DIODE(_01873_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06225__B (.DIODE(_04260_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06226__A (.DIODE(_02544_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06226__B (.DIODE(_04293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06228__A (.DIODE(_02049_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06228__B (.DIODE(_01158_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06233__A (.DIODE(_01807_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06234__A (.DIODE(_03160_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06234__B (.DIODE(_00204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06236__A (.DIODE(_03182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06236__B (.DIODE(_01774_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06239__A (.DIODE(_05031_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06239__B (.DIODE(_01884_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06247__A (.DIODE(_04928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06247__B (.DIODE(_05029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06248__A (.DIODE(_05028_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06248__B (.DIODE(_05032_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06250__A (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__06250__B (.DIODE(_03820_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06282__A (.DIODE(_04962_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06282__B (.DIODE(_04819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06283__A (.DIODE(_04809_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06284__A (.DIODE(_04964_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06284__B (.DIODE(_00254_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06286__A (.DIODE(_03809_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06286__B (.DIODE(_04827_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06292__A (.DIODE(_04812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06293__A (.DIODE(_04911_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06294__A (.DIODE(_04808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06294__B (.DIODE(_04895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06295__A (.DIODE(_00263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06295__B (.DIODE(_00264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06307__A (.DIODE(_04873_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06307__B (.DIODE(_04992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06345__A (.DIODE(_01147_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06345__B (.DIODE(_02357_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06346__A (.DIODE(_01037_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06346__B (.DIODE(_02379_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06348__A (.DIODE(_02544_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06348__B (.DIODE(_00861_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06398__A (.DIODE(_00368_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06409__A (.DIODE(_00784_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06409__B (.DIODE(_01048_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06411__B (.DIODE(_01323_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06411__C (.DIODE(_04293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06412__A (.DIODE(_01323_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06412__B (.DIODE(_04293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06415__A (.DIODE(_00740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06415__B (.DIODE(_01158_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06420__A (.DIODE(_00751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06420__B (.DIODE(_05160_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06423__A (.DIODE(_00795_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06423__B (.DIODE(_00393_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06428__A (.DIODE(_00861_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06428__B (.DIODE(_04084_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06441__A (.DIODE(_01774_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06442__A (.DIODE(_01081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06442__B (.DIODE(_00412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06443__A (.DIODE(_00850_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06443__B (.DIODE(_00204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06447__A (.DIODE(_01037_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06447__B (.DIODE(_00003_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06474__A (.DIODE(_02544_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06474__B (.DIODE(_02995_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06475__A (.DIODE(_01147_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06475__B (.DIODE(_03028_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06479__A (.DIODE(_03215_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06479__B (.DIODE(_01873_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06487__A (.DIODE(_04962_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06487__B (.DIODE(_03160_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06488__A (.DIODE(_04964_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06488__B (.DIODE(_02049_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06492__A (.DIODE(_03809_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06492__B (.DIODE(_03182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06521__A (.DIODE(_04808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06521__B (.DIODE(_05028_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06522__A (.DIODE(_04812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06522__B (.DIODE(_05031_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06526__A (.DIODE(_04818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06526__B (.DIODE(_04928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06546__A (.DIODE(_04871_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06546__B (.DIODE(_04809_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06547__A (.DIODE(_04873_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06547__B (.DIODE(_03820_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06551__A (.DIODE(_04819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06552__A (.DIODE(_04876_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06552__B (.DIODE(_00522_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06558__A (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA__06559__A (.DIODE(_00529_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06559__B (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06561__A (.DIODE(_00124_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06561__B (.DIODE(_04911_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06562__A (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__06562__B (.DIODE(_04827_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06606__A2 (.DIODE(_00141_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06611__A (.DIODE(_00581_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06618__C (.DIODE(_00581_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06633__B (.DIODE(_00602_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06639__C (.DIODE(_00368_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06640__B (.DIODE(_00610_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06645__A (.DIODE(_00615_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06645__B (.DIODE(_00368_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06664__A (.DIODE(_02049_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06664__B (.DIODE(_04260_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06665__A (.DIODE(_01873_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06665__B (.DIODE(_04293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06667__A (.DIODE(_03160_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06667__B (.DIODE(_01565_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06672__A (.DIODE(_05031_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06672__B (.DIODE(_00412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06674__A (.DIODE(_03182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06674__B (.DIODE(_00204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06677__A (.DIODE(_05028_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06677__B (.DIODE(_00003_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06685__A (.DIODE(_03820_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06686__A (.DIODE(_00656_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06686__B (.DIODE(_05029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06687__A (.DIODE(_04928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06687__B (.DIODE(_05032_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06689__A (.DIODE(_03215_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06689__B (.DIODE(_04809_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06719__A1 (.DIODE(_00263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06719__A2 (.DIODE(_00264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06721__A (.DIODE(_03809_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06721__B (.DIODE(_04911_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06722__A (.DIODE(_04962_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06722__B (.DIODE(_04828_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06723__A (.DIODE(_04964_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06723__B (.DIODE(_00522_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06761__A (.DIODE(_02544_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06761__B (.DIODE(_00751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06762__A (.DIODE(_01147_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06762__B (.DIODE(_00795_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06764__A (.DIODE(_01873_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06764__B (.DIODE(_00861_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06818__B (.DIODE(_00793_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06819__A (.DIODE(_00793_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06820__A (.DIODE(_00615_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06820__C (.DIODE(_00368_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06867__A (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__06867__B (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA__06868__A (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__06868__B (.DIODE(_00795_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06870__A (.DIODE(_02049_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06870__B (.DIODE(_00861_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06875__A (.DIODE(_03160_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06875__B (.DIODE(_01048_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06877__A (.DIODE(_02049_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06877__B (.DIODE(_01092_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06882__A (.DIODE(_03094_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06882__B (.DIODE(_01158_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06901__A (.DIODE(_04928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06901__B (.DIODE(_00003_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06902__A (.DIODE(_05028_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06902__B (.DIODE(_00412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06904__A (.DIODE(_05031_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06904__B (.DIODE(_00204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06917__A (.DIODE(_00254_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06917__B (.DIODE(_05029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06918__A (.DIODE(_00656_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06918__B (.DIODE(_05032_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06920__A (.DIODE(_03215_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06920__B (.DIODE(_04819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06970__A (.DIODE(_04812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06970__B (.DIODE(_04992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06971__A (.DIODE(_03809_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06971__B (.DIODE(_04895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06972__A (.DIODE(_04962_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06972__B (.DIODE(_04911_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06974__A (.DIODE(_04964_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06974__B (.DIODE(_04828_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07035__A (.DIODE(_02049_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07035__B (.DIODE(_00751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07036__A (.DIODE(_01873_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07036__B (.DIODE(_00795_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07038__A (.DIODE(_03160_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07038__B (.DIODE(_00861_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07043__A (.DIODE(_03094_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07043__B (.DIODE(_01048_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07045__A (.DIODE(_02753_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07045__B (.DIODE(_01092_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07049__A (.DIODE(_03226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07049__B (.DIODE(_01158_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07068__A (.DIODE(_04928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07068__B (.DIODE(_01774_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07070__A (.DIODE(_03314_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07070__B (.DIODE(_01807_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07073__A (.DIODE(_00656_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07073__B (.DIODE(_01884_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07099__A (.DIODE(_00522_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07099__B (.DIODE(_05029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07100__A (.DIODE(_00254_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07100__B (.DIODE(_05032_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07102__A (.DIODE(_03215_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07102__B (.DIODE(_04828_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07149__B (.DIODE(_01156_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07149__C (.DIODE(_01157_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07150__A (.DIODE(_01156_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07150__B (.DIODE(_01157_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07154__B (.DIODE(_01156_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07156__A1 (.DIODE(_01164_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07156__A2 (.DIODE(_00793_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07157__B (.DIODE(_00793_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07157__C (.DIODE(_01164_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07161__A2 (.DIODE(_00610_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07163__A (.DIODE(_03226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07163__B (.DIODE(_01048_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07164__A (.DIODE(_03094_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07164__B (.DIODE(_01092_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07166__A (.DIODE(_05028_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07166__B (.DIODE(_01158_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07183__A (.DIODE(_03160_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07183__B (.DIODE(_00751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07184__A (.DIODE(_02049_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07184__B (.DIODE(_02379_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07186__A (.DIODE(_03182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07186__B (.DIODE(_00861_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07213__A (.DIODE(_03820_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07213__B (.DIODE(_01774_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07214__A (.DIODE(_03402_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07214__B (.DIODE(_01807_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07216__A (.DIODE(_04809_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07216__B (.DIODE(_01884_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07243__A (.DIODE(_03182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07243__B (.DIODE(_00751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07244__A (.DIODE(_03160_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07244__B (.DIODE(_00795_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07246__A (.DIODE(_05031_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07246__B (.DIODE(_00861_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07251__A (.DIODE(_05028_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07251__B (.DIODE(_04260_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07252__A (.DIODE(_05031_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07252__B (.DIODE(_01092_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07256__A (.DIODE(_04928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07256__B (.DIODE(_01158_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07265__A (.DIODE(_00254_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07265__B (.DIODE(_00412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07266__A (.DIODE(_00656_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07266__B (.DIODE(_00204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07268__A (.DIODE(_00522_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07268__B (.DIODE(_00003_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07294__A (.DIODE(_04827_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07294__B (.DIODE(_05029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07295__A (.DIODE(_00522_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07295__B (.DIODE(_05032_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07297__A (.DIODE(_03215_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07297__B (.DIODE(_04911_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07305__A (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__07306__A (.DIODE(_04962_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07306__B (.DIODE(_04895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07307__A (.DIODE(_01330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07307__B (.DIODE(_00264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07309__A1 (.DIODE(_01330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07309__A2 (.DIODE(_00264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07325__A (.DIODE(_04911_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07325__B (.DIODE(_05029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07326__A (.DIODE(_04828_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07326__B (.DIODE(_05032_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07328__A (.DIODE(_03215_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07328__B (.DIODE(_04895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07333__A (.DIODE(_04964_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07333__B (.DIODE(_04895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07425__A (.DIODE(_03402_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07425__B (.DIODE(_01048_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07426__A (.DIODE(_03314_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07426__B (.DIODE(_01092_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07428__A (.DIODE(_00656_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07428__B (.DIODE(_01565_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07433__A (.DIODE(_00522_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07433__B (.DIODE(_00412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07435__A (.DIODE(_00254_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07435__B (.DIODE(_00204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07438__A (.DIODE(_04828_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07438__B (.DIODE(_00003_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07456__A (.DIODE(_04991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07456__B (.DIODE(_04895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07456__C (.DIODE(_05032_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07456__D (.DIODE(_05029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07491__A (.DIODE(_00861_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07492__A (.DIODE(_05028_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07492__B (.DIODE(_01535_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07493__A (.DIODE(_05031_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07493__B (.DIODE(_00751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07494__A (.DIODE(_03182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07494__B (.DIODE(_00795_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07547__A (.DIODE(_03226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07548__A (.DIODE(_00795_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07549__A (.DIODE(_03314_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07549__B (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA__07550__A2 (.DIODE(_01597_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07551__A (.DIODE(_04928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07551__B (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__07554__B (.DIODE(_05031_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07554__C (.DIODE(_00795_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07559__A (.DIODE(_00254_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07559__B (.DIODE(_01565_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07560__A (.DIODE(_00656_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07560__B (.DIODE(_04260_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07561__A (.DIODE(_04928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07561__B (.DIODE(_04293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07582__A (.DIODE(_04991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07582__B (.DIODE(_00003_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07583__A (.DIODE(_04827_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07583__B (.DIODE(_01774_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07584__A (.DIODE(_00522_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07584__B (.DIODE(_00204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07709__A (.DIODE(_01164_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07709__B (.DIODE(_00793_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07736__A (.DIODE(_03402_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07736__B (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA__07737__A (.DIODE(_03314_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07737__B (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA__07739__A (.DIODE(_03820_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07739__B (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__07745__A (.DIODE(_04809_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07745__B (.DIODE(_01048_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07746__A (.DIODE(_03820_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07746__B (.DIODE(_01092_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07751__A (.DIODE(_04819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07751__B (.DIODE(_01158_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07772__A (.DIODE(_04895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07772__B (.DIODE(_00003_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07773__A (.DIODE(_04911_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07773__B (.DIODE(_00412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07774__A (.DIODE(_04827_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07774__B (.DIODE(_00204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07787__A1 (.DIODE(_04991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07787__A2 (.DIODE(_05032_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07787__B1 (.DIODE(_04992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07787__B2 (.DIODE(_05029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07828__A (.DIODE(_00656_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07828__B (.DIODE(_00751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07829__A (.DIODE(_04928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07829__B (.DIODE(_00795_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07831__A (.DIODE(_04809_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07831__B (.DIODE(_00861_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07837__A (.DIODE(_04827_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07837__B (.DIODE(_01565_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07838__A (.DIODE(_04819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07838__B (.DIODE(_01048_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07839__A (.DIODE(_00254_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07839__B (.DIODE(_01092_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07857__A (.DIODE(_01807_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07858__A (.DIODE(_04895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07858__B (.DIODE(_00412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07859__A (.DIODE(_00264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07859__B (.DIODE(_01937_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07874__A (.DIODE(_04992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07875__A (.DIODE(_03028_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07877__B (.DIODE(_01957_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07878__A2 (.DIODE(_01957_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07946__A (.DIODE(_00522_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07946__B (.DIODE(_01535_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07947__A (.DIODE(_00254_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07947__B (.DIODE(_00751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07948__A (.DIODE(_00656_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07948__B (.DIODE(_02379_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07955__A (.DIODE(_04827_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07955__B (.DIODE(_01048_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07956__A (.DIODE(_04819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07956__B (.DIODE(_01092_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07960__A (.DIODE(_04911_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07960__B (.DIODE(_01158_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07969__A1 (.DIODE(_00264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07969__A2 (.DIODE(_01937_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07991__A (.DIODE(_04827_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07992__A (.DIODE(_01092_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07993__A (.DIODE(_04911_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07993__B (.DIODE(_04260_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07994__B (.DIODE(_02086_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07996__A2 (.DIODE(_02086_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07997__A (.DIODE(_04895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07997__B (.DIODE(_01565_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08004__A1 (.DIODE(_00254_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08004__A2 (.DIODE(_02379_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08004__B1 (.DIODE(_00522_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08004__B2 (.DIODE(_02357_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08005__A (.DIODE(_04828_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08005__B (.DIODE(_01535_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08007__A (.DIODE(_00254_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08007__B (.DIODE(_00522_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08007__C (.DIODE(_02379_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08007__D (.DIODE(_02357_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08013__A (.DIODE(_04895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08013__B (.DIODE(_00204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08097__A (.DIODE(_04991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08097__B (.DIODE(_01535_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08098__A (.DIODE(_00522_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08098__B (.DIODE(_04828_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08098__C (.DIODE(_02379_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08098__D (.DIODE(_02357_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08099__A1 (.DIODE(_00522_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08099__A2 (.DIODE(_02379_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08099__B1 (.DIODE(_04828_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08099__B2 (.DIODE(_02357_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08105__A (.DIODE(_04991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08105__B (.DIODE(_04992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08105__C (.DIODE(_04293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08105__D (.DIODE(_04260_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08107__A1 (.DIODE(_04991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08107__A2 (.DIODE(_04293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08107__B1 (.DIODE(_04992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08107__B2 (.DIODE(_04260_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08139__A (.DIODE(_04992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08139__B (.DIODE(_04293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08140__A (.DIODE(_04992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08140__B (.DIODE(_01535_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08141__A (.DIODE(_04991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08141__B (.DIODE(_02357_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08142__B (.DIODE(_01597_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08143__A2 (.DIODE(_01597_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08182__A2 (.DIODE(_01535_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08182__C1 (.DIODE(_01597_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08214__A (.DIODE(_00861_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08214__B (.DIODE(_05160_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08216__A (.DIODE(_00751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08216__B (.DIODE(_00393_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08217__A (.DIODE(_00795_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08217__B (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__08230__A (.DIODE(_00784_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08230__B (.DIODE(_01565_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08232__A (.DIODE(_01323_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08232__B (.DIODE(_01048_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08233__A (.DIODE(_04293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08233__B (.DIODE(_04084_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08246__A (.DIODE(_01081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08246__B (.DIODE(_00003_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08247__A (.DIODE(_00850_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08247__B (.DIODE(_01774_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08248__A (.DIODE(_00740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08248__B (.DIODE(_01807_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08271__A (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__08271__B (.DIODE(_02995_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08272__A (.DIODE(_01037_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08272__B (.DIODE(_03028_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08276__A (.DIODE(_03215_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08276__B (.DIODE(_02544_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08286__A (.DIODE(_03809_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08286__B (.DIODE(_02753_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08287__A (.DIODE(_01873_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08288__A (.DIODE(_04962_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08288__B (.DIODE(_02049_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08289__A (.DIODE(_01330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08291__A1 (.DIODE(_01330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08318__B (.DIODE(_02443_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08319__A (.DIODE(_02443_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08323__A (.DIODE(_04876_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08323__B (.DIODE(_04809_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08324__A (.DIODE(_03402_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08325__A (.DIODE(_04871_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08325__B (.DIODE(_03820_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08334__A (.DIODE(_00529_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08334__B (.DIODE(_04991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08335__A (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__08336__A (.DIODE(_04819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08337__A (.DIODE(_00124_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08337__B (.DIODE(_04827_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08347__A (.DIODE(_04818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08347__B (.DIODE(_05028_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08348__A (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__08348__B (.DIODE(_03226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08349__A (.DIODE(_04812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08349__B (.DIODE(_03094_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08389__B (.DIODE(_02521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08390__A (.DIODE(_02521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08393__A (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__08393__B (.DIODE(_04992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08414__A (.DIODE(_02549_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08419__A (.DIODE(_01535_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08419__B (.DIODE(_00393_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08420__A (.DIODE(_00751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08420__B (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__08422__A (.DIODE(_00795_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08434__A (.DIODE(_04260_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08434__B (.DIODE(_04084_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08435__A (.DIODE(_04293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08435__B (.DIODE(_05160_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08438__A (.DIODE(_01323_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08438__B (.DIODE(_01565_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08451__A (.DIODE(_00740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08451__B (.DIODE(_00412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08452__A (.DIODE(_00784_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08452__B (.DIODE(_00204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08455__A (.DIODE(_00850_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08455__B (.DIODE(_00003_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08477__A (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__08478__B (.DIODE(_02995_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08479__B (.DIODE(_01957_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08479__C (.DIODE(_02620_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08481__A2 (.DIODE(_01957_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08481__B1 (.DIODE(_02620_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08482__A (.DIODE(_03215_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08482__B (.DIODE(_01147_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08492__A (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__08492__B (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA__08494__A (.DIODE(_04962_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08494__B (.DIODE(_01873_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08495__A (.DIODE(_04964_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08495__B (.DIODE(_02544_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08524__A (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__08524__B (.DIODE(_03094_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08525__A (.DIODE(_04812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08525__B (.DIODE(_02753_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08528__A (.DIODE(_04818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08528__B (.DIODE(_03226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08549__A (.DIODE(_03314_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08550__A (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__08550__B (.DIODE(_03402_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08554__A (.DIODE(_04876_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08554__B (.DIODE(_03820_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08565__A (.DIODE(_00529_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08565__B (.DIODE(_04828_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08566__A (.DIODE(_00124_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08566__B (.DIODE(_04819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08607__A (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__08607__B (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__08607__C (.DIODE(_04911_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08607__D (.DIODE(_04895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08609__A1 (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__08609__A2 (.DIODE(_04991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08609__B1 (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__08609__B2 (.DIODE(_04895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08651__B (.DIODE(_02549_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08667__B (.DIODE(_00602_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08668__A_N (.DIODE(_00602_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08675__A (.DIODE(_02357_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08676__A (.DIODE(_02379_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08679__A (.DIODE(_01535_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08679__B (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__08688__A (.DIODE(_01048_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08688__B (.DIODE(_05160_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08689__A (.DIODE(_01092_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08689__B (.DIODE(_00393_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08692__A (.DIODE(_01565_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08692__B (.DIODE(_04084_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08705__A (.DIODE(_01323_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08706__A (.DIODE(_00784_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08706__B (.DIODE(_00412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08707__B (.DIODE(_01937_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08708__A2 (.DIODE(_01937_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08710__A (.DIODE(_00740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08710__B (.DIODE(_00003_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08728__A (.DIODE(_01081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08728__B (.DIODE(_02995_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08729__B (.DIODE(_01957_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08731__A2 (.DIODE(_01957_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08732__A (.DIODE(_03215_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08732__B (.DIODE(_01037_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08742__A (.DIODE(_03809_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08742__B (.DIODE(_01873_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08744__A (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__08745__A (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__08745__B (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__08746__A (.DIODE(_01330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08747__A1 (.DIODE(_01330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08779__A (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA__08780__A (.DIODE(_04808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08780__B (.DIODE(_02753_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08781__A (.DIODE(_00263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08782__A1 (.DIODE(_00263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08784__A (.DIODE(_04818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08784__B (.DIODE(_03182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08788__A (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__08789__A1 (.DIODE(_01330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08790__A (.DIODE(_01330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08810__A (.DIODE(_04871_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08810__B (.DIODE(_03314_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08814__A (.DIODE(_04876_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08814__B (.DIODE(_03402_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08822__A (.DIODE(_00529_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08822__B (.DIODE(_04819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08824__A (.DIODE(_00124_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08824__B (.DIODE(_04809_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08825__A (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__08825__B (.DIODE(_03820_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08856__B (.DIODE(_03035_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08861__A (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__08862__A (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__08862__B (.DIODE(_04911_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08866__A (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA__08866__B (.DIODE(_04895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08897__A (.DIODE(_03035_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08903__A (.DIODE(_02357_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08904__A (.DIODE(_01597_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08906__A1 (.DIODE(_01597_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08907__A (.DIODE(_01535_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08916__A (.DIODE(_01565_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08916__B (.DIODE(_05160_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08918__A (.DIODE(_04260_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08918__B (.DIODE(_00393_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08919__A (.DIODE(_04293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08919__B (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__08935__A (.DIODE(_00784_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08935__B (.DIODE(_00003_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08937__A (.DIODE(_01323_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08937__B (.DIODE(_00412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08938__A (.DIODE(_00204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08938__B (.DIODE(_04084_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08961__A (.DIODE(_03809_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08961__B (.DIODE(_02544_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08963__A (.DIODE(_04962_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08963__B (.DIODE(_01147_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08964__A (.DIODE(_04964_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08964__B (.DIODE(_01037_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08969__A (.DIODE(_03215_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08969__B (.DIODE(_01081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08971__A (.DIODE(_00850_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08971__B (.DIODE(_05029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08972__A (.DIODE(_00740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08972__B (.DIODE(_05032_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08996__A (.DIODE(_04818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08996__B (.DIODE(_03160_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08998__A (.DIODE(_04808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08998__B (.DIODE(_02049_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08999__A (.DIODE(_00263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09000__A1 (.DIODE(_00263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09020__A (.DIODE(_04876_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09020__B (.DIODE(_05028_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09022__A (.DIODE(_04873_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09022__B (.DIODE(_04871_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09022__C (.DIODE(_03094_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09022__D (.DIODE(_03226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09023__A1 (.DIODE(_04873_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09023__A2 (.DIODE(_03182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09023__B1 (.DIODE(_04871_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09023__B2 (.DIODE(_05031_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09033__A (.DIODE(_00529_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09033__B (.DIODE(_00254_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09034__A (.DIODE(_00124_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09034__B (.DIODE(_00656_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09072__A (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA__09072__B (.DIODE(_04991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09074__A (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__09074__B (.DIODE(_04828_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09081__A (.DIODE(_00656_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09106__A (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__09106__B (.DIODE(_04992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09139__A (.DIODE(_03035_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09141__A (.DIODE(_03035_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09187__A (.DIODE(_02327_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09188__A (.DIODE(_00602_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09198__A (.DIODE(_04876_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09198__B (.DIODE(_05031_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09199__A (.DIODE(_04873_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09199__B (.DIODE(_04871_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09199__C (.DIODE(_03160_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09199__D (.DIODE(_03182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09201__A1 (.DIODE(_04873_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09201__A2 (.DIODE(_03160_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09201__B1 (.DIODE(_04871_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09201__B2 (.DIODE(_03182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09209__A (.DIODE(_00529_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09209__B (.DIODE(_00656_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09210__A (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__09210__B (.DIODE(_00124_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09210__C (.DIODE(_05028_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09210__D (.DIODE(_04928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09211__A1 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__09211__A2 (.DIODE(_05028_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09211__B1 (.DIODE(_00124_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09211__B2 (.DIODE(_04928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09219__A (.DIODE(_04818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09219__B (.DIODE(_02049_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09220__A (.DIODE(_04812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09220__B (.DIODE(_04808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09220__C (.DIODE(_02544_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09220__D (.DIODE(_01873_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09221__A1 (.DIODE(_04812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09221__A2 (.DIODE(_02544_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09221__B1 (.DIODE(_04808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09221__B2 (.DIODE(_01873_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09226__A (.DIODE(_01037_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09227__A (.DIODE(_01330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09255__A (.DIODE(_01535_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09256__A (.DIODE(_02379_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09256__B (.DIODE(_02357_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09257__A1 (.DIODE(_02379_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09257__B1 (.DIODE(_02357_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09267__A (.DIODE(_01565_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09267__B (.DIODE(_00393_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09269__A (.DIODE(_04260_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09269__B (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__09270__A (.DIODE(_02086_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09271__A1 (.DIODE(_02086_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09281__A (.DIODE(_01323_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09281__B (.DIODE(_00003_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09282__A (.DIODE(_00204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09282__B (.DIODE(_00412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09282__C (.DIODE(_04084_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09282__D (.DIODE(_05160_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09283__A1 (.DIODE(_00204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09283__A2 (.DIODE(_05160_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09283__B1 (.DIODE(_00412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09283__B2 (.DIODE(_04084_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09288__A (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__09289__A (.DIODE(_02086_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09295__A (.DIODE(_04084_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09296__A (.DIODE(_01937_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09311__A (.DIODE(_03215_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09311__B (.DIODE(_00850_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09313__A (.DIODE(_00784_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09313__B (.DIODE(_00740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09313__C (.DIODE(_05032_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09313__D (.DIODE(_02995_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09315__A1 (.DIODE(_00784_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09315__A2 (.DIODE(_05032_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09315__B1 (.DIODE(_00740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09315__B2 (.DIODE(_05029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09323__A (.DIODE(_03809_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09323__B (.DIODE(_01147_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09324__A (.DIODE(_04964_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09324__B (.DIODE(_04962_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09324__C (.DIODE(_01081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09324__D (.DIODE(_01037_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09325__A1 (.DIODE(_04964_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09325__A2 (.DIODE(_01081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09325__B1 (.DIODE(_04962_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09325__B2 (.DIODE(_01037_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09361__A (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__09361__B (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__09361__C (.DIODE(_04809_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09361__D (.DIODE(_04819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09363__A1 (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__09363__A2 (.DIODE(_00254_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09363__B1 (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__09363__B2 (.DIODE(_00522_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09366__A (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA__09366__B (.DIODE(_04828_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09390__A (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__09391__A (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__09392__C (.DIODE(_00264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09393__A1 (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__09393__A2 (.DIODE(_04991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09393__B1 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__09393__B2 (.DIODE(_04992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09437__A (.DIODE(_00003_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09437__B (.DIODE(_04084_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09438__A (.DIODE(_00204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09438__B (.DIODE(_00412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09438__C (.DIODE(_05160_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09438__D (.DIODE(_00393_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09440__A1 (.DIODE(_00204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09440__A2 (.DIODE(_00393_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09440__B1 (.DIODE(_00412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09440__B2 (.DIODE(_05160_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09453__A (.DIODE(_01535_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09454__A (.DIODE(_02379_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09454__B (.DIODE(_02357_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09455__A1 (.DIODE(_02379_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09455__B1 (.DIODE(_02357_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09459__A2 (.DIODE(_01535_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09463__A (.DIODE(_01565_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09463__B (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__09464__A (.DIODE(_04293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09464__B (.DIODE(_04260_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09466__A1 (.DIODE(_04293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09466__B1 (.DIODE(_04260_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09485__A (.DIODE(_01323_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09485__B (.DIODE(_00784_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09485__C (.DIODE(_05032_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09485__D (.DIODE(_05029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09487__A1 (.DIODE(_01323_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09487__A2 (.DIODE(_05032_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09487__B1 (.DIODE(_00784_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09487__B2 (.DIODE(_05029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09489__A (.DIODE(_03215_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09489__B (.DIODE(_00740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09496__A (.DIODE(_03809_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09496__B (.DIODE(_01037_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09497__A (.DIODE(_04964_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09497__B (.DIODE(_04962_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09497__C (.DIODE(_00850_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09497__D (.DIODE(_01081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09499__A1 (.DIODE(_04964_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09499__A2 (.DIODE(_00850_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09499__B1 (.DIODE(_04962_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09499__B2 (.DIODE(_01081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09527__A2 (.DIODE(_03809_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09527__A3 (.DIODE(_01147_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09528__A (.DIODE(_04812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09528__B (.DIODE(_04808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09528__C (.DIODE(_01147_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09528__D (.DIODE(_02544_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09530__A1 (.DIODE(_04812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09530__A2 (.DIODE(_01147_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09530__B1 (.DIODE(_04808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09530__B2 (.DIODE(_02544_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09533__A (.DIODE(_04818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09533__B (.DIODE(_01873_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09547__A (.DIODE(_04876_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09547__B (.DIODE(_03182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09548__A (.DIODE(_04871_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09549__D_N (.DIODE(_03160_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09550__A1 (.DIODE(_04873_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09550__A2 (.DIODE(_02049_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09550__B1 (.DIODE(_04871_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09550__B2 (.DIODE(_03160_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09560__A (.DIODE(_00529_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09560__B (.DIODE(_04928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09562__A (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__09562__B (.DIODE(_00124_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09562__C (.DIODE(_05031_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09562__D (.DIODE(_05028_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09563__A1 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__09563__A2 (.DIODE(_05031_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09563__B1 (.DIODE(_00124_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09563__B2 (.DIODE(_05028_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09596__A2 (.DIODE(_00529_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09596__A3 (.DIODE(_00656_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09597__A (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__09597__B (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__09597__C (.DIODE(_00656_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09597__D (.DIODE(_00254_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09599__A1 (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__09599__A2 (.DIODE(_00656_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09599__B1 (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__09599__B2 (.DIODE(_00254_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09601__A (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA__09601__B (.DIODE(_00522_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09628__A (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA__09628__B (.DIODE(_04992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09629__A (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__09629__B (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__09629__C (.DIODE(_04828_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09629__D (.DIODE(_04991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09630__A1 (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__09630__A2 (.DIODE(_04828_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09630__B1 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__09630__B2 (.DIODE(_04991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09684__A (.DIODE(_04818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09684__B (.DIODE(_02544_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09685__A (.DIODE(_04808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09686__A (.DIODE(_00263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09687__A1 (.DIODE(_04812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09687__A2 (.DIODE(_01037_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09687__B1 (.DIODE(_04808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09687__B2 (.DIODE(_01147_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09709__A (.DIODE(_04876_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09709__B (.DIODE(_03160_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09711__A1 (.DIODE(_04873_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09711__A2 (.DIODE(_01873_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09711__B1 (.DIODE(_04871_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09711__B2 (.DIODE(_02049_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09720__A (.DIODE(_00529_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09720__B (.DIODE(_05028_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09722__A (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__09722__B (.DIODE(_00124_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09722__C (.DIODE(_03182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09722__D (.DIODE(_05031_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09723__A1 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__09723__A2 (.DIODE(_03182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09723__B1 (.DIODE(_00124_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09723__B2 (.DIODE(_05031_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09748__A (.DIODE(_01535_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09750__A (.DIODE(_02357_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09751__A (.DIODE(_01597_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09752__A1 (.DIODE(_01597_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09755__A2 (.DIODE(_01535_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09760__A (.DIODE(_01565_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09761__A (.DIODE(_04260_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09762__A (.DIODE(_02086_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09763__A1 (.DIODE(_02086_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09775__A (.DIODE(_00003_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09775__B (.DIODE(_05160_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09776__A (.DIODE(_00412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09776__B (.DIODE(_00393_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09777__A (.DIODE(_01937_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09779__A1 (.DIODE(_01937_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09803__A (.DIODE(_03215_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09803__B (.DIODE(_00784_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09804__A (.DIODE(_05029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09805__B (.DIODE(_01957_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09806__A1 (.DIODE(_01323_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09806__A2 (.DIODE(_05029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09806__B1 (.DIODE(_05032_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09806__B2 (.DIODE(_04084_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09816__A (.DIODE(_03809_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09816__B (.DIODE(_01081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09817__A (.DIODE(_04964_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09817__B (.DIODE(_04962_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09817__C (.DIODE(_00740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09817__D (.DIODE(_00850_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09818__A1 (.DIODE(_04964_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09818__A2 (.DIODE(_00740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09818__B1 (.DIODE(_04962_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09818__B2 (.DIODE(_00850_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09854__A (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA__09854__B (.DIODE(_00254_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09855__A (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__09857__A1 (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__09857__A2 (.DIODE(_04928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09857__B1 (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__09857__B2 (.DIODE(_00656_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09887__A (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__09887__B (.DIODE(_04992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09888__A2 (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA__09888__A3 (.DIODE(_04992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09889__A (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA__09889__B (.DIODE(_04991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09891__A1 (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__09891__A2 (.DIODE(_00522_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09891__B1 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__09891__B2 (.DIODE(_04828_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09940__A (.DIODE(_04225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09942__B (.DIODE(_04225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09951__A (.DIODE(_03215_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09951__B (.DIODE(_01323_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09953__A (.DIODE(_01957_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09953__D_N (.DIODE(_05160_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09954__A1 (.DIODE(_05032_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09954__A2 (.DIODE(_05160_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09954__B1 (.DIODE(_05029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09954__B2 (.DIODE(_04084_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09960__A (.DIODE(_03809_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09960__B (.DIODE(_00850_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09962__A (.DIODE(_04962_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09962__B (.DIODE(_00740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09963__A (.DIODE(_04964_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09963__B (.DIODE(_00784_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09980__A (.DIODE(_01565_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09981__A (.DIODE(_04293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09981__B (.DIODE(_04260_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09982__A1 (.DIODE(_04293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09982__B1 (.DIODE(_04260_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09985__A2 (.DIODE(_01535_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09986__A (.DIODE(_01535_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09987__A (.DIODE(_02357_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09988__A (.DIODE(_02379_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09998__A (.DIODE(_00003_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09998__B (.DIODE(_00393_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09999__A (.DIODE(_00412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09999__B (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__10000__A (.DIODE(_00204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10003__A2 (.DIODE(_01565_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10024__A2 (.DIODE(_03809_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10024__A3 (.DIODE(_01081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10026__A (.DIODE(_04818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10026__B (.DIODE(_01147_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10027__A (.DIODE(_00263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10028__A1 (.DIODE(_04812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10028__A2 (.DIODE(_01081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10028__B1 (.DIODE(_04808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10028__B2 (.DIODE(_01037_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10043__A (.DIODE(_04876_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10043__B (.DIODE(_02049_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10045__A1 (.DIODE(_04873_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10045__A2 (.DIODE(_02544_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10045__B1 (.DIODE(_04871_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10045__B2 (.DIODE(_01873_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10050__A (.DIODE(_00529_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10050__B (.DIODE(_05031_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10051__A (.DIODE(_00124_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10051__B (.DIODE(_03182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10052__A (.DIODE(_03160_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10052__B (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__10083__A (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA__10083__B (.DIODE(_00656_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10085__A1 (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__10085__A2 (.DIODE(_05028_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10085__B1 (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__10085__B2 (.DIODE(_04928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10111__A (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__10111__B (.DIODE(_04991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10112__A (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA__10112__B (.DIODE(_04828_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10114__A1 (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__10114__A2 (.DIODE(_00254_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10114__B1 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__10114__B2 (.DIODE(_00522_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10126__A (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__10126__B (.DIODE(_04992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10171__B (.DIODE(_04225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10172__A_N (.DIODE(_04225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10174__B (.DIODE(_04485_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10175__A (.DIODE(_04485_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10436__B (.DIODE(_02327_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10437__A (.DIODE(_02327_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10443__A1 (.DIODE(_02327_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10458__CLK (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__10459__CLK (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__10460__CLK (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__10461__CLK (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__10462__CLK (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__10463__CLK (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__10464__CLK (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__10465__CLK (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__10466__CLK (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__10467__CLK (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__10467__RESET_B (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__10468__CLK (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__10468__RESET_B (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__10469__CLK (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__10469__RESET_B (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__10470__CLK (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__10470__RESET_B (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__10471__CLK (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__10471__RESET_B (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__10472__CLK (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__10472__RESET_B (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__10473__CLK (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__10474__CLK (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__10475__CLK (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__10476__CLK (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__10477__CLK (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__10478__CLK (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__10479__CLK (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__10480__CLK (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__10481__CLK (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__10482__CLK (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__10483__CLK (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__10484__CLK (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__10485__CLK (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__10486__CLK (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__10487__CLK (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__10487__RESET_B (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__10488__CLK (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__10488__RESET_B (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__10489__CLK (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__10489__RESET_B (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__10490__CLK (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__10490__RESET_B (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__10491__CLK (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__10491__RESET_B (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__10492__CLK (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__10492__RESET_B (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__10493__CLK (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__10493__RESET_B (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__10494__CLK (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__10494__RESET_B (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__10495__CLK (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__10495__RESET_B (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__10496__CLK (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__10497__CLK (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__10498__CLK (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__10499__CLK (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__10500__CLK (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__10501__CLK (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__10502__CLK (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__10503__CLK (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__10504__CLK (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__10505__CLK (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__10505__RESET_B (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__10506__CLK (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__10506__RESET_B (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__10507__CLK (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__10507__RESET_B (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__10508__CLK (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__10508__RESET_B (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__10509__CLK (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__10509__RESET_B (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__10510__CLK (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__10510__RESET_B (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__10511__CLK (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__10511__RESET_B (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_0__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_1__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_2__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_3__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout100_A (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout101_A (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout98_A (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout99_A (.DIODE(net101));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_560 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_610 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_192 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_259 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_351 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_358 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_374 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_395 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_443 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_49 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_598 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_602 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_179 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_348 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_384 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_42 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_490 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_585 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_593 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_112 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_116 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_300 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_491 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_511 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_536 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_572 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_600 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_72 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_28 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_340 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_406 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_416 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_424 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_438 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_462 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_526 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_540 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_578 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_583 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_67 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_95 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_115 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_135 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_158 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_170 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_256 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_342 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_380 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_392 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_490 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_500 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_504 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_518 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_538 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_550 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_555 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_563 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_59 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_91 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_10 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_16 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_220 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_262 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_303 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_347 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_460 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_534 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_570 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_60 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_64 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_150 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_203 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_210 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_239 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_290 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_322 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_340 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_348 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_40 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_432 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_444 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_493 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_92 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_183 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_198 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_206 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_266 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_329 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_40 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_406 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_410 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_424 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_441 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_564 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_571 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_592 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_64 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_107 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_119 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_242 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_406 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_443 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_453 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_574 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_99 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_127 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_180 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_296 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_308 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_332 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_356 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_413 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_430 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_479 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_534 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_578 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_590 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_607 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_95 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_322 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_464 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_470 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_123 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_161 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_182 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_219 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_239 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_320 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_383 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_416 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_435 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_504 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_508 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_516 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_104 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_11 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_130 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_240 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_257 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_276 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_298 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_302 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_324 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_399 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_416 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_468 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_534 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_621 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_135 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_144 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_204 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_238 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_260 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_272 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_327 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_462 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_470 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_490 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_550 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_562 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_252 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_267 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_402 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_420 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_490 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_526 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_564 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_576 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_588 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_103 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_378 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_410 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_414 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_439 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_443 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_456 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_46 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_569 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_135 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_155 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_232 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_359 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_536 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_592 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_598 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_114 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_148 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_256 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_260 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_313 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_392 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_459 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_491 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_538 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_560 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_619 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_132 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_144 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_176 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_183 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_260 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_303 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_440 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_571 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_603 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_67 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_285 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_407 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_460 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_470 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_504 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_551 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_563 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_598 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_604 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_140 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_180 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_300 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_35 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_356 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_379 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_484 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_535 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_546 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_570 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_594 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_61 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_84 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_426 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_438 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_498 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_519 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_560 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_147 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_172 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_220 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_383 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_397 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_436 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_50 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_539 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_555 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_95 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_127 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_371 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_410 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_590 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_115 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_119 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_158 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_188 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_204 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_235 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_270 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_294 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_430 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_45 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_497 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_515 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_555 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_566 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_606 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_611 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_147 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_183 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_243 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_247 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_28 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_35 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_570 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_574 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_624 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_87 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_170 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_276 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_547 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_556 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_564 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_599 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_603 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_88 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_314 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_364 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_420 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_491 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_575 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_583 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_594 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_604 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_610 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_107 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_154 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_285 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_336 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_375 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_387 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_434 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_526 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_546 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_624 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_196 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_204 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_28 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_356 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_360 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_364 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_420 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_44 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_49 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_529 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_535 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_577 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_95 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_159 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_275 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_282 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_342 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_399 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_483 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_546 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_580 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_142 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_201 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_241 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_434 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_464 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_476 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_60 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_99 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_308 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_11 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_114 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_282 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_292 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_300 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_318 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_338 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_357 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_375 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_392 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_426 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_450 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_499 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_52 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_563 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_586 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_67 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_72 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_480 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_513 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_582 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_609 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_95 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_171 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_182 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_248 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_300 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_303 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_336 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_380 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_392 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_438 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_450 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_480 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_484 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_491 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_580 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_119 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_131 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_151 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_215 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_342 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_375 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_452 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_491 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_552 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_624 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_271 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_298 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_315 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_408 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_43 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_519 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_547 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_551 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_580 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_76 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_100 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_172 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_184 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_198 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_211 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_254 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_266 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_32 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_40 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_435 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_469 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_494 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_509 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_519 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_537 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_624 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_462 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_579 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_618 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_74 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_182 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_201 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_292 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_310 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_411 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_414 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_426 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_432 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_478 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_532 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_548 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_87 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_161 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_173 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_238 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_282 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_438 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_506 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_525 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_546 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_56 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_66 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_8 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_186 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_266 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_294 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_386 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_478 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_524 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_567 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_588 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_592 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_275 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_336 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_354 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_392 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_428 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_448 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_464 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_515 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_540 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_555 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_114 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_132 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_186 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_228 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_273 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_276 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_284 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_350 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_458 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_513 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_563 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_586 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_606 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_238 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_292 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_359 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_364 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_400 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_422 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_546 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_564 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_612 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_68 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_88 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_210 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_24 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_434 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_450 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_454 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_457 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_127 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_230 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_295 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_423 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_444 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_468 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_495 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_532 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_569 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_580 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_86 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_117 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_156 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_168 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_217 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_269 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_280 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_299 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_369 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_426 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_504 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_516 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_560 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_586 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_592 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_98 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_140 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_220 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_360 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_364 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_406 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_434 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_515 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_582 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_604 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_242 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_270 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_324 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_336 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_432 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_499 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_564 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_592 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_229 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_254 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_357 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_380 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_495 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_522 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_534 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_542 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_92 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_179 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_248 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_274 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_286 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_296 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_300 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_324 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_37 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_438 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_448 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_472 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_492 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_512 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_541 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_108 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_127 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_142 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_239 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_288 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_308 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_313 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_547 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_567 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_88 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_98 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_254 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_369 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_378 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_420 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_565 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_568 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_596 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_238 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_42 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_487 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_491 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_556 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_560 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_586 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_67 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_151 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_242 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_407 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_412 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_48 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_529 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_551 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_575 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_603 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_84 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_128 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_134 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_159 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_203 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_280 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_316 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_450 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_480 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_492 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_557 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_566 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_599 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_241 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_266 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_469 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_591 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_67 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_71 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_91 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_151 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_159 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_25 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_392 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_564 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_621 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_74 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_78 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_236 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_248 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_270 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_285 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_459 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_471 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_487 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_49 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_515 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_580 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_584 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_592 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_13 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_392 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_440 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_526 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_542 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_550 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_58 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_582 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_98 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_134 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_217 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_235 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_263 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_444 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_46 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_464 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_497 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_588 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_603 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_95 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_155 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_173 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_216 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_360 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_426 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_434 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_522 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_526 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_19 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_214 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_246 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_308 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_423 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_509 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_532 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_577 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_582 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_590 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_94 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_275 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_495 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_594 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_64 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_152 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_338 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_342 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_434 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_520 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_524 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_563 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_592 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_596 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_600 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_618 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_99 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_210 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_367 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_402 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_422 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_426 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_604 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_208 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_264 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_378 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_434 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_438 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_444 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_49 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_506 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_539 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_568 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_584 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_602 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_95 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_126 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_247 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_319 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_357 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_369 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_420 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_462 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_494 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_498 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_550 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_568 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_576 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_580 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_588 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_210 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_272 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_282 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_380 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_397 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_434 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_438 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_544 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_604 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_620 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_106 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_131 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_196 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_208 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_240 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_276 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_351 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_382 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_464 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_524 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_572 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_583 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_620 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_105 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_302 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_322 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_33 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_351 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_395 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_416 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_538 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_542 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_562 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_611 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_7 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_230 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_255 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_271 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_340 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_400 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_427 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_463 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_535 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_567 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_582 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_272 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_288 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_313 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_338 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_472 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_563 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_140 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_147 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_155 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_172 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_375 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_379 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_471 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_99 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_308 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_358 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_366 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_464 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_476 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_519 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_554 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_571 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_575 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_315 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_319 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_388 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_392 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_442 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_455 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_464 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_470 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_507 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_536 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_562 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_579 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_596 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_63 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_144 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_17 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_288 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_356 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_42 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_459 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_523 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_590 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_112 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_217 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_274 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_292 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_322 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_351 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_399 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_484 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_496 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_56 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_80 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_94 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_100 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_212 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_410 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_422 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_464 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_481 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_515 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_525 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_535 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_571 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_88 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_11 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_154 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_204 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_280 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_319 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_518 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_596 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_117 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_247 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_255 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_264 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_302 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_434 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_46 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_466 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_484 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_229 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_382 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_394 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_428 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_441 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_464 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_513 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_565 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_609 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_180 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_330 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_368 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_372 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_380 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_40 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_416 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_434 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_581 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_234 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_322 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_35 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_414 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_448 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_463 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_562 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_59 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_605 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_12 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_299 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_311 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_409 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_43 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_436 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_541 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_581 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_154 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_162 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_168 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_176 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_381 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_408 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_495 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_506 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_563 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_576 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_64 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_201 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_219 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_336 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_402 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_451 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_459 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_508 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_598 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_606 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_61 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_622 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_178 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_234 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_302 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_424 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_462 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_492 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_526 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_557 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_570 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_590 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_323 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_356 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_493 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_560 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_564 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_616 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_301 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_36 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_364 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_388 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_420 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_436 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_470 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_522 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_588 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_176 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_226 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_381 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_441 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_451 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_459 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_207 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_228 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_232 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_31 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_320 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_351 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_43 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_478 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_490 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_571 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_583 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_620 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_171 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_215 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_271 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_399 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_49 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_510 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_602 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_610 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_182 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_235 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_36 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_422 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_463 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_491 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_554 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_566 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_10 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_190 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_210 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_214 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_295 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_410 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_458 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_46 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_470 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_479 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_487 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_523 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_588 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_600 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_364 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_43 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_485 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_516 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_576 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_93 ();
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_148 ();
 sky130_fd_sc_hd__decap_3 PHY_149 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_150 ();
 sky130_fd_sc_hd__decap_3 PHY_151 ();
 sky130_fd_sc_hd__decap_3 PHY_152 ();
 sky130_fd_sc_hd__decap_3 PHY_153 ();
 sky130_fd_sc_hd__decap_3 PHY_154 ();
 sky130_fd_sc_hd__decap_3 PHY_155 ();
 sky130_fd_sc_hd__decap_3 PHY_156 ();
 sky130_fd_sc_hd__decap_3 PHY_157 ();
 sky130_fd_sc_hd__decap_3 PHY_158 ();
 sky130_fd_sc_hd__decap_3 PHY_159 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_160 ();
 sky130_fd_sc_hd__decap_3 PHY_161 ();
 sky130_fd_sc_hd__decap_3 PHY_162 ();
 sky130_fd_sc_hd__decap_3 PHY_163 ();
 sky130_fd_sc_hd__decap_3 PHY_164 ();
 sky130_fd_sc_hd__decap_3 PHY_165 ();
 sky130_fd_sc_hd__decap_3 PHY_166 ();
 sky130_fd_sc_hd__decap_3 PHY_167 ();
 sky130_fd_sc_hd__decap_3 PHY_168 ();
 sky130_fd_sc_hd__decap_3 PHY_169 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_170 ();
 sky130_fd_sc_hd__decap_3 PHY_171 ();
 sky130_fd_sc_hd__decap_3 PHY_172 ();
 sky130_fd_sc_hd__decap_3 PHY_173 ();
 sky130_fd_sc_hd__decap_3 PHY_174 ();
 sky130_fd_sc_hd__decap_3 PHY_175 ();
 sky130_fd_sc_hd__decap_3 PHY_176 ();
 sky130_fd_sc_hd__decap_3 PHY_177 ();
 sky130_fd_sc_hd__decap_3 PHY_178 ();
 sky130_fd_sc_hd__decap_3 PHY_179 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_180 ();
 sky130_fd_sc_hd__decap_3 PHY_181 ();
 sky130_fd_sc_hd__decap_3 PHY_182 ();
 sky130_fd_sc_hd__decap_3 PHY_183 ();
 sky130_fd_sc_hd__decap_3 PHY_184 ();
 sky130_fd_sc_hd__decap_3 PHY_185 ();
 sky130_fd_sc_hd__decap_3 PHY_186 ();
 sky130_fd_sc_hd__decap_3 PHY_187 ();
 sky130_fd_sc_hd__decap_3 PHY_188 ();
 sky130_fd_sc_hd__decap_3 PHY_189 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_190 ();
 sky130_fd_sc_hd__decap_3 PHY_191 ();
 sky130_fd_sc_hd__decap_3 PHY_192 ();
 sky130_fd_sc_hd__decap_3 PHY_193 ();
 sky130_fd_sc_hd__decap_3 PHY_194 ();
 sky130_fd_sc_hd__decap_3 PHY_195 ();
 sky130_fd_sc_hd__decap_3 PHY_196 ();
 sky130_fd_sc_hd__decap_3 PHY_197 ();
 sky130_fd_sc_hd__decap_3 PHY_198 ();
 sky130_fd_sc_hd__decap_3 PHY_199 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_200 ();
 sky130_fd_sc_hd__decap_3 PHY_201 ();
 sky130_fd_sc_hd__decap_3 PHY_202 ();
 sky130_fd_sc_hd__decap_3 PHY_203 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_999 ();
 sky130_fd_sc_hd__clkbuf_8 _05202_ (.A(net10),
    .X(_00740_));
 sky130_fd_sc_hd__buf_12 _05203_ (.A(net44),
    .X(_00751_));
 sky130_fd_sc_hd__nand2_1 _05204_ (.A(_00740_),
    .B(_00751_),
    .Y(_00762_));
 sky130_fd_sc_hd__inv_2 _05205_ (.A(_00762_),
    .Y(_00773_));
 sky130_fd_sc_hd__buf_4 _05206_ (.A(net11),
    .X(_00784_));
 sky130_fd_sc_hd__buf_12 _05207_ (.A(net33),
    .X(_00795_));
 sky130_fd_sc_hd__nand2_1 _05208_ (.A(_00784_),
    .B(_00795_),
    .Y(_00806_));
 sky130_fd_sc_hd__nand2_1 _05209_ (.A(_00773_),
    .B(_00806_),
    .Y(_00817_));
 sky130_fd_sc_hd__inv_2 _05210_ (.A(_00806_),
    .Y(_00828_));
 sky130_fd_sc_hd__nand2_1 _05211_ (.A(_00828_),
    .B(_00762_),
    .Y(_00839_));
 sky130_fd_sc_hd__clkbuf_8 _05212_ (.A(net9),
    .X(_00850_));
 sky130_fd_sc_hd__buf_8 _05213_ (.A(net55),
    .X(_00861_));
 sky130_fd_sc_hd__nand2_1 _05214_ (.A(_00850_),
    .B(_00861_),
    .Y(_00872_));
 sky130_fd_sc_hd__nand3_1 _05215_ (.A(_00817_),
    .B(_00839_),
    .C(_00872_),
    .Y(_00883_));
 sky130_fd_sc_hd__nand2_1 _05216_ (.A(_00773_),
    .B(_00828_),
    .Y(_00894_));
 sky130_fd_sc_hd__inv_2 _05217_ (.A(_00872_),
    .Y(_00905_));
 sky130_fd_sc_hd__nand2_1 _05218_ (.A(_00762_),
    .B(_00806_),
    .Y(_00916_));
 sky130_fd_sc_hd__nand3_1 _05219_ (.A(_00894_),
    .B(_00905_),
    .C(_00916_),
    .Y(_00927_));
 sky130_fd_sc_hd__nand2_1 _05220_ (.A(_00883_),
    .B(_00927_),
    .Y(_00938_));
 sky130_fd_sc_hd__nand2_2 _05221_ (.A(_00850_),
    .B(_00751_),
    .Y(_00949_));
 sky130_fd_sc_hd__nand2_2 _05222_ (.A(_00740_),
    .B(_00795_),
    .Y(_00960_));
 sky130_fd_sc_hd__nand2_1 _05223_ (.A(_00949_),
    .B(_00960_),
    .Y(_00971_));
 sky130_fd_sc_hd__nand2_1 _05224_ (.A(net8),
    .B(net55),
    .Y(_00982_));
 sky130_fd_sc_hd__inv_2 _05225_ (.A(_00982_),
    .Y(_00993_));
 sky130_fd_sc_hd__nor2_1 _05226_ (.A(_00949_),
    .B(_00960_),
    .Y(_01004_));
 sky130_fd_sc_hd__a21oi_2 _05227_ (.A1(_00971_),
    .A2(_00993_),
    .B1(_01004_),
    .Y(_01015_));
 sky130_fd_sc_hd__nand2_1 _05228_ (.A(_00938_),
    .B(_01015_),
    .Y(_01026_));
 sky130_fd_sc_hd__buf_8 _05229_ (.A(net7),
    .X(_01037_));
 sky130_fd_sc_hd__buf_8 _05230_ (.A(net59),
    .X(_01048_));
 sky130_fd_sc_hd__nand2_2 _05231_ (.A(_01037_),
    .B(_01048_),
    .Y(_01059_));
 sky130_fd_sc_hd__inv_2 _05232_ (.A(_01059_),
    .Y(_01070_));
 sky130_fd_sc_hd__clkbuf_8 _05233_ (.A(net8),
    .X(_01081_));
 sky130_fd_sc_hd__buf_8 _05234_ (.A(net58),
    .X(_01092_));
 sky130_fd_sc_hd__nand2_1 _05235_ (.A(_01081_),
    .B(_01092_),
    .Y(_01103_));
 sky130_fd_sc_hd__nand2_1 _05236_ (.A(_01070_),
    .B(_01103_),
    .Y(_01114_));
 sky130_fd_sc_hd__inv_2 _05237_ (.A(_01103_),
    .Y(_01125_));
 sky130_fd_sc_hd__nand2_1 _05238_ (.A(_01125_),
    .B(_01059_),
    .Y(_01136_));
 sky130_fd_sc_hd__buf_8 _05239_ (.A(net6),
    .X(_01147_));
 sky130_fd_sc_hd__buf_6 _05240_ (.A(net60),
    .X(_01158_));
 sky130_fd_sc_hd__nand2_1 _05241_ (.A(_01147_),
    .B(_01158_),
    .Y(_01169_));
 sky130_fd_sc_hd__nand3_1 _05242_ (.A(_01114_),
    .B(_01136_),
    .C(_01169_),
    .Y(_01180_));
 sky130_fd_sc_hd__nand2_1 _05243_ (.A(_01070_),
    .B(_01125_),
    .Y(_01191_));
 sky130_fd_sc_hd__inv_2 _05244_ (.A(_01169_),
    .Y(_01202_));
 sky130_fd_sc_hd__nand2_1 _05245_ (.A(_01059_),
    .B(_01103_),
    .Y(_01213_));
 sky130_fd_sc_hd__nand3_1 _05246_ (.A(_01191_),
    .B(_01202_),
    .C(_01213_),
    .Y(_01224_));
 sky130_fd_sc_hd__nand2_1 _05247_ (.A(_01180_),
    .B(_01224_),
    .Y(_01235_));
 sky130_fd_sc_hd__inv_2 _05248_ (.A(_01235_),
    .Y(_01246_));
 sky130_fd_sc_hd__nor2_1 _05249_ (.A(_01015_),
    .B(_00938_),
    .Y(_01257_));
 sky130_fd_sc_hd__a21oi_1 _05250_ (.A1(_01026_),
    .A2(_01246_),
    .B1(_01257_),
    .Y(_01268_));
 sky130_fd_sc_hd__nor2_1 _05251_ (.A(_00762_),
    .B(_00806_),
    .Y(_01279_));
 sky130_fd_sc_hd__a21o_1 _05252_ (.A1(_00916_),
    .A2(_00905_),
    .B1(_01279_),
    .X(_01290_));
 sky130_fd_sc_hd__nand2_1 _05253_ (.A(_00784_),
    .B(_00751_),
    .Y(_01301_));
 sky130_fd_sc_hd__inv_2 _05254_ (.A(_01301_),
    .Y(_01312_));
 sky130_fd_sc_hd__buf_4 _05255_ (.A(net13),
    .X(_01323_));
 sky130_fd_sc_hd__nand2_1 _05256_ (.A(_01323_),
    .B(_00795_),
    .Y(_01334_));
 sky130_fd_sc_hd__inv_2 _05257_ (.A(_01334_),
    .Y(_01345_));
 sky130_fd_sc_hd__nand2_1 _05258_ (.A(_01312_),
    .B(_01345_),
    .Y(_01356_));
 sky130_fd_sc_hd__nand2_1 _05259_ (.A(_00740_),
    .B(_00861_),
    .Y(_01367_));
 sky130_fd_sc_hd__inv_2 _05260_ (.A(_01367_),
    .Y(_01378_));
 sky130_fd_sc_hd__nand2_1 _05261_ (.A(_01301_),
    .B(_01334_),
    .Y(_01389_));
 sky130_fd_sc_hd__nand3_1 _05262_ (.A(_01356_),
    .B(_01378_),
    .C(_01389_),
    .Y(_01400_));
 sky130_fd_sc_hd__nand2_1 _05263_ (.A(_01312_),
    .B(_01334_),
    .Y(_01411_));
 sky130_fd_sc_hd__nand2_1 _05264_ (.A(_01345_),
    .B(_01301_),
    .Y(_01422_));
 sky130_fd_sc_hd__nand3_1 _05265_ (.A(_01411_),
    .B(_01422_),
    .C(_01367_),
    .Y(_01433_));
 sky130_fd_sc_hd__nand3_1 _05266_ (.A(_01290_),
    .B(_01400_),
    .C(_01433_),
    .Y(_01444_));
 sky130_fd_sc_hd__nand2_1 _05267_ (.A(_01433_),
    .B(_01400_),
    .Y(_01455_));
 sky130_fd_sc_hd__a21oi_1 _05268_ (.A1(_00916_),
    .A2(_00905_),
    .B1(_01279_),
    .Y(_01466_));
 sky130_fd_sc_hd__nand2_1 _05269_ (.A(_01455_),
    .B(_01466_),
    .Y(_01477_));
 sky130_fd_sc_hd__nand2_1 _05270_ (.A(_01081_),
    .B(_01048_),
    .Y(_01488_));
 sky130_fd_sc_hd__inv_2 _05271_ (.A(_01488_),
    .Y(_01499_));
 sky130_fd_sc_hd__nand2_1 _05272_ (.A(_00850_),
    .B(_01092_),
    .Y(_01510_));
 sky130_fd_sc_hd__inv_2 _05273_ (.A(_01510_),
    .Y(_01521_));
 sky130_fd_sc_hd__nand2_1 _05274_ (.A(_01499_),
    .B(_01521_),
    .Y(_01532_));
 sky130_fd_sc_hd__nand2_1 _05275_ (.A(_01488_),
    .B(_01510_),
    .Y(_01543_));
 sky130_fd_sc_hd__nand2_1 _05276_ (.A(_01532_),
    .B(_01543_),
    .Y(_01554_));
 sky130_fd_sc_hd__buf_8 _05277_ (.A(_01158_),
    .X(_01565_));
 sky130_fd_sc_hd__nand2_1 _05278_ (.A(_01037_),
    .B(_01565_),
    .Y(_01576_));
 sky130_fd_sc_hd__nand2_1 _05279_ (.A(_01554_),
    .B(_01576_),
    .Y(_01587_));
 sky130_fd_sc_hd__inv_2 _05280_ (.A(_01576_),
    .Y(_01598_));
 sky130_fd_sc_hd__nand3_1 _05281_ (.A(_01532_),
    .B(_01598_),
    .C(_01543_),
    .Y(_01609_));
 sky130_fd_sc_hd__nand2_1 _05282_ (.A(_01587_),
    .B(_01609_),
    .Y(_01620_));
 sky130_fd_sc_hd__inv_2 _05283_ (.A(_01620_),
    .Y(_01631_));
 sky130_fd_sc_hd__nand3_1 _05284_ (.A(_01444_),
    .B(_01477_),
    .C(_01631_),
    .Y(_01642_));
 sky130_fd_sc_hd__nand2_1 _05285_ (.A(_01455_),
    .B(_01290_),
    .Y(_01653_));
 sky130_fd_sc_hd__nand3_1 _05286_ (.A(_01466_),
    .B(_01433_),
    .C(_01400_),
    .Y(_01664_));
 sky130_fd_sc_hd__nand3_1 _05287_ (.A(_01653_),
    .B(_01664_),
    .C(_01620_),
    .Y(_01675_));
 sky130_fd_sc_hd__nand3_1 _05288_ (.A(_01268_),
    .B(_01642_),
    .C(_01675_),
    .Y(_01686_));
 sky130_fd_sc_hd__inv_2 _05289_ (.A(_01015_),
    .Y(_01697_));
 sky130_fd_sc_hd__nand3_1 _05290_ (.A(_01697_),
    .B(_00927_),
    .C(_00883_),
    .Y(_01708_));
 sky130_fd_sc_hd__nand3_1 _05291_ (.A(_01708_),
    .B(_01026_),
    .C(_01246_),
    .Y(_01719_));
 sky130_fd_sc_hd__nand2_1 _05292_ (.A(_01719_),
    .B(_01708_),
    .Y(_01730_));
 sky130_fd_sc_hd__nand2_1 _05293_ (.A(_01642_),
    .B(_01675_),
    .Y(_01741_));
 sky130_fd_sc_hd__nand2_1 _05294_ (.A(_01730_),
    .B(_01741_),
    .Y(_01752_));
 sky130_fd_sc_hd__nand2_1 _05295_ (.A(_01686_),
    .B(_01752_),
    .Y(_01763_));
 sky130_fd_sc_hd__clkbuf_8 _05296_ (.A(net62),
    .X(_01774_));
 sky130_fd_sc_hd__nand2_1 _05297_ (.A(net5),
    .B(_01774_),
    .Y(_01785_));
 sky130_fd_sc_hd__inv_2 _05298_ (.A(_01785_),
    .Y(_01796_));
 sky130_fd_sc_hd__clkbuf_8 _05299_ (.A(net61),
    .X(_01807_));
 sky130_fd_sc_hd__nand2_1 _05300_ (.A(net6),
    .B(_01807_),
    .Y(_01818_));
 sky130_fd_sc_hd__inv_2 _05301_ (.A(_01818_),
    .Y(_01829_));
 sky130_fd_sc_hd__nand2_1 _05302_ (.A(_01796_),
    .B(_01829_),
    .Y(_01840_));
 sky130_fd_sc_hd__nand2_1 _05303_ (.A(_01785_),
    .B(_01818_),
    .Y(_01851_));
 sky130_fd_sc_hd__nand2_1 _05304_ (.A(_01840_),
    .B(_01851_),
    .Y(_01862_));
 sky130_fd_sc_hd__buf_6 _05305_ (.A(net4),
    .X(_01873_));
 sky130_fd_sc_hd__buf_6 _05306_ (.A(net63),
    .X(_01884_));
 sky130_fd_sc_hd__nand2_1 _05307_ (.A(_01873_),
    .B(_01884_),
    .Y(_01895_));
 sky130_fd_sc_hd__nand2_1 _05308_ (.A(_01862_),
    .B(_01895_),
    .Y(_01906_));
 sky130_fd_sc_hd__nand3b_2 _05309_ (.A_N(_01895_),
    .B(_01840_),
    .C(_01851_),
    .Y(_01917_));
 sky130_fd_sc_hd__nand2_1 _05310_ (.A(_01906_),
    .B(_01917_),
    .Y(_01928_));
 sky130_fd_sc_hd__nor2_1 _05311_ (.A(_01059_),
    .B(_01103_),
    .Y(_01939_));
 sky130_fd_sc_hd__a21oi_1 _05312_ (.A1(_01213_),
    .A2(_01202_),
    .B1(_01939_),
    .Y(_01950_));
 sky130_fd_sc_hd__nand2_1 _05313_ (.A(_01928_),
    .B(_01950_),
    .Y(_01961_));
 sky130_fd_sc_hd__a21o_1 _05314_ (.A1(_01213_),
    .A2(_01202_),
    .B1(_01939_),
    .X(_01972_));
 sky130_fd_sc_hd__nand3_1 _05315_ (.A(_01972_),
    .B(_01917_),
    .C(_01906_),
    .Y(_01983_));
 sky130_fd_sc_hd__nand2_1 _05316_ (.A(net5),
    .B(_01807_),
    .Y(_01994_));
 sky130_fd_sc_hd__inv_2 _05317_ (.A(_01994_),
    .Y(_02005_));
 sky130_fd_sc_hd__nand2_1 _05318_ (.A(net4),
    .B(_01774_),
    .Y(_02016_));
 sky130_fd_sc_hd__inv_2 _05319_ (.A(_02016_),
    .Y(_02027_));
 sky130_fd_sc_hd__nand2_1 _05320_ (.A(_02005_),
    .B(_02027_),
    .Y(_02038_));
 sky130_fd_sc_hd__buf_6 _05321_ (.A(net3),
    .X(_02049_));
 sky130_fd_sc_hd__nand2_1 _05322_ (.A(_02049_),
    .B(_01884_),
    .Y(_02060_));
 sky130_fd_sc_hd__inv_2 _05323_ (.A(_02060_),
    .Y(_02071_));
 sky130_fd_sc_hd__nand2_1 _05324_ (.A(_01994_),
    .B(_02016_),
    .Y(_02082_));
 sky130_fd_sc_hd__nand3_2 _05325_ (.A(_02038_),
    .B(_02071_),
    .C(_02082_),
    .Y(_02093_));
 sky130_fd_sc_hd__nand2_1 _05326_ (.A(_02093_),
    .B(_02038_),
    .Y(_02104_));
 sky130_fd_sc_hd__nand3_1 _05327_ (.A(_01961_),
    .B(_01983_),
    .C(_02104_),
    .Y(_02115_));
 sky130_fd_sc_hd__nand2_1 _05328_ (.A(_01928_),
    .B(_01972_),
    .Y(_02126_));
 sky130_fd_sc_hd__nand3_1 _05329_ (.A(_01906_),
    .B(_01917_),
    .C(_01950_),
    .Y(_02137_));
 sky130_fd_sc_hd__inv_2 _05330_ (.A(_02104_),
    .Y(_02148_));
 sky130_fd_sc_hd__nand3_1 _05331_ (.A(_02126_),
    .B(_02137_),
    .C(_02148_),
    .Y(_02159_));
 sky130_fd_sc_hd__nand2_1 _05332_ (.A(_02115_),
    .B(_02159_),
    .Y(_02170_));
 sky130_fd_sc_hd__inv_2 _05333_ (.A(_02170_),
    .Y(_02181_));
 sky130_fd_sc_hd__nand2_1 _05334_ (.A(_01763_),
    .B(_02181_),
    .Y(_02192_));
 sky130_fd_sc_hd__nand3_1 _05335_ (.A(_01686_),
    .B(_01752_),
    .C(_02170_),
    .Y(_02203_));
 sky130_fd_sc_hd__nand2_1 _05336_ (.A(_02192_),
    .B(_02203_),
    .Y(_02214_));
 sky130_fd_sc_hd__nand2_1 _05337_ (.A(_00938_),
    .B(_01697_),
    .Y(_02225_));
 sky130_fd_sc_hd__nand3_1 _05338_ (.A(_01015_),
    .B(_00883_),
    .C(_00927_),
    .Y(_02236_));
 sky130_fd_sc_hd__nand3_1 _05339_ (.A(_02225_),
    .B(_02236_),
    .C(_01235_),
    .Y(_02247_));
 sky130_fd_sc_hd__nand2_1 _05340_ (.A(_01719_),
    .B(_02247_),
    .Y(_02258_));
 sky130_fd_sc_hd__inv_2 _05341_ (.A(_00949_),
    .Y(_02269_));
 sky130_fd_sc_hd__nand2_1 _05342_ (.A(_02269_),
    .B(_00960_),
    .Y(_02280_));
 sky130_fd_sc_hd__inv_2 _05343_ (.A(_00960_),
    .Y(_02291_));
 sky130_fd_sc_hd__nand2_1 _05344_ (.A(_02291_),
    .B(_00949_),
    .Y(_02302_));
 sky130_fd_sc_hd__nand3_1 _05345_ (.A(_02280_),
    .B(_02302_),
    .C(_00982_),
    .Y(_02313_));
 sky130_fd_sc_hd__nand2_1 _05346_ (.A(_02269_),
    .B(_02291_),
    .Y(_02324_));
 sky130_fd_sc_hd__nand3_1 _05347_ (.A(_02324_),
    .B(_00993_),
    .C(_00971_),
    .Y(_02335_));
 sky130_fd_sc_hd__nand2_1 _05348_ (.A(_02313_),
    .B(_02335_),
    .Y(_02346_));
 sky130_fd_sc_hd__buf_8 _05349_ (.A(_00751_),
    .X(_02357_));
 sky130_fd_sc_hd__nand2_2 _05350_ (.A(_01081_),
    .B(_02357_),
    .Y(_02368_));
 sky130_fd_sc_hd__buf_12 _05351_ (.A(_00795_),
    .X(_02379_));
 sky130_fd_sc_hd__nand2_2 _05352_ (.A(_00850_),
    .B(_02379_),
    .Y(_02390_));
 sky130_fd_sc_hd__nand2_1 _05353_ (.A(_02368_),
    .B(_02390_),
    .Y(_02401_));
 sky130_fd_sc_hd__nand2_1 _05354_ (.A(_01037_),
    .B(_00861_),
    .Y(_02412_));
 sky130_fd_sc_hd__inv_2 _05355_ (.A(_02412_),
    .Y(_02423_));
 sky130_fd_sc_hd__nor2_1 _05356_ (.A(_02368_),
    .B(_02390_),
    .Y(_02434_));
 sky130_fd_sc_hd__a21oi_2 _05357_ (.A1(_02401_),
    .A2(_02423_),
    .B1(_02434_),
    .Y(_02445_));
 sky130_fd_sc_hd__nand2_1 _05358_ (.A(_02346_),
    .B(_02445_),
    .Y(_02456_));
 sky130_fd_sc_hd__nand2_1 _05359_ (.A(_01147_),
    .B(_01048_),
    .Y(_02467_));
 sky130_fd_sc_hd__inv_2 _05360_ (.A(_02467_),
    .Y(_02478_));
 sky130_fd_sc_hd__nand2_1 _05361_ (.A(net7),
    .B(_01092_),
    .Y(_02489_));
 sky130_fd_sc_hd__nand2_1 _05362_ (.A(_02478_),
    .B(_02489_),
    .Y(_02500_));
 sky130_fd_sc_hd__inv_2 _05363_ (.A(_02489_),
    .Y(_02511_));
 sky130_fd_sc_hd__nand2_1 _05364_ (.A(_02511_),
    .B(_02467_),
    .Y(_02522_));
 sky130_fd_sc_hd__nand2_1 _05365_ (.A(_02500_),
    .B(_02522_),
    .Y(_02533_));
 sky130_fd_sc_hd__buf_8 _05366_ (.A(net5),
    .X(_02544_));
 sky130_fd_sc_hd__nand2_1 _05367_ (.A(_02544_),
    .B(_01158_),
    .Y(_02555_));
 sky130_fd_sc_hd__inv_2 _05368_ (.A(_02555_),
    .Y(_02566_));
 sky130_fd_sc_hd__nand2_1 _05369_ (.A(_02533_),
    .B(_02566_),
    .Y(_02577_));
 sky130_fd_sc_hd__nand3_1 _05370_ (.A(_02500_),
    .B(_02522_),
    .C(_02555_),
    .Y(_02588_));
 sky130_fd_sc_hd__nand2_1 _05371_ (.A(_02577_),
    .B(_02588_),
    .Y(_02599_));
 sky130_fd_sc_hd__inv_2 _05372_ (.A(_02599_),
    .Y(_02610_));
 sky130_fd_sc_hd__nor2_1 _05373_ (.A(_02445_),
    .B(_02346_),
    .Y(_02621_));
 sky130_fd_sc_hd__a21oi_1 _05374_ (.A1(_02456_),
    .A2(_02610_),
    .B1(_02621_),
    .Y(_02632_));
 sky130_fd_sc_hd__nand2_1 _05375_ (.A(_02258_),
    .B(_02632_),
    .Y(_02643_));
 sky130_fd_sc_hd__nand2_1 _05376_ (.A(_02038_),
    .B(_02082_),
    .Y(_02654_));
 sky130_fd_sc_hd__nand2_1 _05377_ (.A(_02654_),
    .B(_02060_),
    .Y(_02665_));
 sky130_fd_sc_hd__nand2_1 _05378_ (.A(_02665_),
    .B(_02093_),
    .Y(_02676_));
 sky130_fd_sc_hd__nand2_1 _05379_ (.A(_02467_),
    .B(_02489_),
    .Y(_02687_));
 sky130_fd_sc_hd__nor2_1 _05380_ (.A(_02467_),
    .B(_02489_),
    .Y(_02698_));
 sky130_fd_sc_hd__a21oi_1 _05381_ (.A1(_02687_),
    .A2(_02566_),
    .B1(_02698_),
    .Y(_02709_));
 sky130_fd_sc_hd__nand2_1 _05382_ (.A(_02676_),
    .B(_02709_),
    .Y(_02720_));
 sky130_fd_sc_hd__a21o_1 _05383_ (.A1(_02687_),
    .A2(_02566_),
    .B1(_02698_),
    .X(_02731_));
 sky130_fd_sc_hd__nand3_1 _05384_ (.A(_02731_),
    .B(_02093_),
    .C(_02665_),
    .Y(_02742_));
 sky130_fd_sc_hd__buf_6 _05385_ (.A(net2),
    .X(_02753_));
 sky130_fd_sc_hd__nand2_1 _05386_ (.A(_02753_),
    .B(_01884_),
    .Y(_02764_));
 sky130_fd_sc_hd__nand2_1 _05387_ (.A(net3),
    .B(_01774_),
    .Y(_02775_));
 sky130_fd_sc_hd__inv_2 _05388_ (.A(_02775_),
    .Y(_02786_));
 sky130_fd_sc_hd__nand2_1 _05389_ (.A(net4),
    .B(_01807_),
    .Y(_02797_));
 sky130_fd_sc_hd__inv_2 _05390_ (.A(_02797_),
    .Y(_02808_));
 sky130_fd_sc_hd__nand2_1 _05391_ (.A(_02786_),
    .B(_02808_),
    .Y(_02819_));
 sky130_fd_sc_hd__nand2_1 _05392_ (.A(_02775_),
    .B(_02797_),
    .Y(_02830_));
 sky130_fd_sc_hd__nand3b_1 _05393_ (.A_N(_02764_),
    .B(_02819_),
    .C(_02830_),
    .Y(_02841_));
 sky130_fd_sc_hd__nand2_1 _05394_ (.A(_02841_),
    .B(_02819_),
    .Y(_02852_));
 sky130_fd_sc_hd__nand3_1 _05395_ (.A(_02720_),
    .B(_02742_),
    .C(_02852_),
    .Y(_02863_));
 sky130_fd_sc_hd__nand2_1 _05396_ (.A(_02676_),
    .B(_02731_),
    .Y(_02874_));
 sky130_fd_sc_hd__nand3_1 _05397_ (.A(_02665_),
    .B(_02709_),
    .C(_02093_),
    .Y(_02885_));
 sky130_fd_sc_hd__inv_2 _05398_ (.A(_02852_),
    .Y(_02896_));
 sky130_fd_sc_hd__nand3_1 _05399_ (.A(_02874_),
    .B(_02885_),
    .C(_02896_),
    .Y(_02907_));
 sky130_fd_sc_hd__nand2_1 _05400_ (.A(_02863_),
    .B(_02907_),
    .Y(_02918_));
 sky130_fd_sc_hd__inv_2 _05401_ (.A(_02918_),
    .Y(_02929_));
 sky130_fd_sc_hd__nor2_1 _05402_ (.A(_02632_),
    .B(_02258_),
    .Y(_02940_));
 sky130_fd_sc_hd__a21oi_2 _05403_ (.A1(_02643_),
    .A2(_02929_),
    .B1(_02940_),
    .Y(_02951_));
 sky130_fd_sc_hd__nand2_1 _05404_ (.A(_02214_),
    .B(_02951_),
    .Y(_02962_));
 sky130_fd_sc_hd__nor2_1 _05405_ (.A(_02709_),
    .B(_02676_),
    .Y(_02973_));
 sky130_fd_sc_hd__a21oi_1 _05406_ (.A1(_02720_),
    .A2(_02852_),
    .B1(_02973_),
    .Y(_02984_));
 sky130_fd_sc_hd__buf_6 _05407_ (.A(net34),
    .X(_02995_));
 sky130_fd_sc_hd__nand2_1 _05408_ (.A(_02753_),
    .B(_02995_),
    .Y(_03006_));
 sky130_fd_sc_hd__inv_2 _05409_ (.A(_03006_),
    .Y(_03017_));
 sky130_fd_sc_hd__buf_4 _05410_ (.A(net64),
    .X(_03028_));
 sky130_fd_sc_hd__nand2_1 _05411_ (.A(net3),
    .B(_03028_),
    .Y(_03039_));
 sky130_fd_sc_hd__inv_2 _05412_ (.A(_03039_),
    .Y(_03050_));
 sky130_fd_sc_hd__nand2_1 _05413_ (.A(_03017_),
    .B(_03050_),
    .Y(_03061_));
 sky130_fd_sc_hd__nand2_1 _05414_ (.A(_03006_),
    .B(_03039_),
    .Y(_03072_));
 sky130_fd_sc_hd__nand2_1 _05415_ (.A(_03061_),
    .B(_03072_),
    .Y(_03083_));
 sky130_fd_sc_hd__clkbuf_8 _05416_ (.A(net32),
    .X(_03094_));
 sky130_fd_sc_hd__nand2_1 _05417_ (.A(net35),
    .B(_03094_),
    .Y(_03105_));
 sky130_fd_sc_hd__nand2_1 _05418_ (.A(_03083_),
    .B(_03105_),
    .Y(_03116_));
 sky130_fd_sc_hd__inv_2 _05419_ (.A(_03105_),
    .Y(_03127_));
 sky130_fd_sc_hd__nand3_1 _05420_ (.A(_03061_),
    .B(_03127_),
    .C(_03072_),
    .Y(_03138_));
 sky130_fd_sc_hd__nand2_1 _05421_ (.A(_03116_),
    .B(_03138_),
    .Y(_03149_));
 sky130_fd_sc_hd__buf_8 _05422_ (.A(_02753_),
    .X(_03160_));
 sky130_fd_sc_hd__nand2_1 _05423_ (.A(_03160_),
    .B(_03028_),
    .Y(_03171_));
 sky130_fd_sc_hd__clkbuf_8 _05424_ (.A(_03094_),
    .X(_03182_));
 sky130_fd_sc_hd__nand2_1 _05425_ (.A(_03182_),
    .B(_02995_),
    .Y(_03193_));
 sky130_fd_sc_hd__nand2_1 _05426_ (.A(_03171_),
    .B(_03193_),
    .Y(_03204_));
 sky130_fd_sc_hd__clkbuf_8 _05427_ (.A(net35),
    .X(_03215_));
 sky130_fd_sc_hd__clkbuf_8 _05428_ (.A(net31),
    .X(_03226_));
 sky130_fd_sc_hd__nand2_1 _05429_ (.A(_03215_),
    .B(_03226_),
    .Y(_03237_));
 sky130_fd_sc_hd__inv_2 _05430_ (.A(_03237_),
    .Y(_03248_));
 sky130_fd_sc_hd__nor2_1 _05431_ (.A(_03171_),
    .B(_03193_),
    .Y(_03259_));
 sky130_fd_sc_hd__a21oi_1 _05432_ (.A1(_03204_),
    .A2(_03248_),
    .B1(_03259_),
    .Y(_03270_));
 sky130_fd_sc_hd__nand2_1 _05433_ (.A(_03149_),
    .B(_03270_),
    .Y(_03281_));
 sky130_fd_sc_hd__a21o_1 _05434_ (.A1(_03204_),
    .A2(_03248_),
    .B1(_03259_),
    .X(_03292_));
 sky130_fd_sc_hd__nand3_1 _05435_ (.A(_03292_),
    .B(_03138_),
    .C(_03116_),
    .Y(_03303_));
 sky130_fd_sc_hd__clkbuf_8 _05436_ (.A(net30),
    .X(_03314_));
 sky130_fd_sc_hd__nand2_1 _05437_ (.A(net37),
    .B(_03314_),
    .Y(_03325_));
 sky130_fd_sc_hd__inv_2 _05438_ (.A(_03325_),
    .Y(_03336_));
 sky130_fd_sc_hd__nand2_1 _05439_ (.A(net36),
    .B(_03226_),
    .Y(_03347_));
 sky130_fd_sc_hd__inv_2 _05440_ (.A(_03347_),
    .Y(_03358_));
 sky130_fd_sc_hd__nand2_1 _05441_ (.A(_03336_),
    .B(_03358_),
    .Y(_03369_));
 sky130_fd_sc_hd__nand2_1 _05442_ (.A(_03325_),
    .B(_03347_),
    .Y(_03380_));
 sky130_fd_sc_hd__nand2_1 _05443_ (.A(_03369_),
    .B(_03380_),
    .Y(_03391_));
 sky130_fd_sc_hd__clkbuf_8 _05444_ (.A(net29),
    .X(_03402_));
 sky130_fd_sc_hd__nand2_1 _05445_ (.A(net38),
    .B(_03402_),
    .Y(_03413_));
 sky130_fd_sc_hd__nand2_1 _05446_ (.A(_03391_),
    .B(_03413_),
    .Y(_03424_));
 sky130_fd_sc_hd__inv_2 _05447_ (.A(_03413_),
    .Y(_03435_));
 sky130_fd_sc_hd__nand3_1 _05448_ (.A(_03369_),
    .B(_03435_),
    .C(_03380_),
    .Y(_03446_));
 sky130_fd_sc_hd__nand2_1 _05449_ (.A(_03424_),
    .B(_03446_),
    .Y(_03457_));
 sky130_fd_sc_hd__inv_2 _05450_ (.A(_03457_),
    .Y(_03468_));
 sky130_fd_sc_hd__nand3_2 _05451_ (.A(_03281_),
    .B(_03303_),
    .C(_03468_),
    .Y(_03479_));
 sky130_fd_sc_hd__nand2_1 _05452_ (.A(_03149_),
    .B(_03292_),
    .Y(_03490_));
 sky130_fd_sc_hd__nand3_1 _05453_ (.A(_03116_),
    .B(_03270_),
    .C(_03138_),
    .Y(_03501_));
 sky130_fd_sc_hd__nand3_1 _05454_ (.A(_03490_),
    .B(_03501_),
    .C(_03457_),
    .Y(_03512_));
 sky130_fd_sc_hd__nand3_1 _05455_ (.A(_02984_),
    .B(_03479_),
    .C(_03512_),
    .Y(_03523_));
 sky130_fd_sc_hd__nand2_1 _05456_ (.A(_03479_),
    .B(_03512_),
    .Y(_03534_));
 sky130_fd_sc_hd__a21oi_1 _05457_ (.A1(_02665_),
    .A2(_02093_),
    .B1(_02731_),
    .Y(_03545_));
 sky130_fd_sc_hd__o21ai_1 _05458_ (.A1(_02896_),
    .A2(_03545_),
    .B1(_02742_),
    .Y(_03556_));
 sky130_fd_sc_hd__nand2_1 _05459_ (.A(_03534_),
    .B(_03556_),
    .Y(_03567_));
 sky130_fd_sc_hd__nand2_1 _05460_ (.A(_03523_),
    .B(_03567_),
    .Y(_03578_));
 sky130_fd_sc_hd__nand3b_1 _05461_ (.A_N(_03259_),
    .B(_03248_),
    .C(_03204_),
    .Y(_03589_));
 sky130_fd_sc_hd__nand2b_1 _05462_ (.A_N(_03193_),
    .B(_03171_),
    .Y(_03600_));
 sky130_fd_sc_hd__nand2b_1 _05463_ (.A_N(_03171_),
    .B(_03193_),
    .Y(_03611_));
 sky130_fd_sc_hd__nand3_1 _05464_ (.A(_03600_),
    .B(_03611_),
    .C(_03237_),
    .Y(_03622_));
 sky130_fd_sc_hd__nand2_1 _05465_ (.A(_03589_),
    .B(_03622_),
    .Y(_03633_));
 sky130_fd_sc_hd__nand2_1 _05466_ (.A(_03226_),
    .B(_02995_),
    .Y(_03644_));
 sky130_fd_sc_hd__nand2_1 _05467_ (.A(_03094_),
    .B(_03028_),
    .Y(_03655_));
 sky130_fd_sc_hd__nand2_1 _05468_ (.A(_03644_),
    .B(_03655_),
    .Y(_03666_));
 sky130_fd_sc_hd__nand2_1 _05469_ (.A(net35),
    .B(_03314_),
    .Y(_03677_));
 sky130_fd_sc_hd__inv_2 _05470_ (.A(_03677_),
    .Y(_03688_));
 sky130_fd_sc_hd__nor2_1 _05471_ (.A(_03644_),
    .B(_03655_),
    .Y(_03699_));
 sky130_fd_sc_hd__a21oi_2 _05472_ (.A1(_03666_),
    .A2(_03688_),
    .B1(_03699_),
    .Y(_03710_));
 sky130_fd_sc_hd__nand2_1 _05473_ (.A(_03633_),
    .B(_03710_),
    .Y(_03721_));
 sky130_fd_sc_hd__inv_2 _05474_ (.A(_03710_),
    .Y(_03732_));
 sky130_fd_sc_hd__nand3_1 _05475_ (.A(_03589_),
    .B(_03732_),
    .C(_03622_),
    .Y(_03743_));
 sky130_fd_sc_hd__nand2_1 _05476_ (.A(net37),
    .B(_03402_),
    .Y(_03754_));
 sky130_fd_sc_hd__nand2_1 _05477_ (.A(net36),
    .B(_03314_),
    .Y(_03765_));
 sky130_fd_sc_hd__nor2_1 _05478_ (.A(_03754_),
    .B(_03765_),
    .Y(_03776_));
 sky130_fd_sc_hd__nand2_1 _05479_ (.A(_03754_),
    .B(_03765_),
    .Y(_03787_));
 sky130_fd_sc_hd__inv_2 _05480_ (.A(_03787_),
    .Y(_03798_));
 sky130_fd_sc_hd__clkbuf_8 _05481_ (.A(net38),
    .X(_03809_));
 sky130_fd_sc_hd__buf_6 _05482_ (.A(net28),
    .X(_03820_));
 sky130_fd_sc_hd__nand2_1 _05483_ (.A(_03809_),
    .B(_03820_),
    .Y(_03831_));
 sky130_fd_sc_hd__o21ai_1 _05484_ (.A1(_03776_),
    .A2(_03798_),
    .B1(_03831_),
    .Y(_03842_));
 sky130_fd_sc_hd__inv_2 _05485_ (.A(_03831_),
    .Y(_03853_));
 sky130_fd_sc_hd__nand3b_1 _05486_ (.A_N(_03776_),
    .B(_03853_),
    .C(_03787_),
    .Y(_03864_));
 sky130_fd_sc_hd__nand2_1 _05487_ (.A(_03842_),
    .B(_03864_),
    .Y(_03875_));
 sky130_fd_sc_hd__inv_2 _05488_ (.A(_03875_),
    .Y(_03886_));
 sky130_fd_sc_hd__nand3_1 _05489_ (.A(_03721_),
    .B(_03743_),
    .C(_03886_),
    .Y(_03897_));
 sky130_fd_sc_hd__nand2_1 _05490_ (.A(_03897_),
    .B(_03743_),
    .Y(_03908_));
 sky130_fd_sc_hd__nand2_1 _05491_ (.A(_03578_),
    .B(_03908_),
    .Y(_03919_));
 sky130_fd_sc_hd__inv_2 _05492_ (.A(_03908_),
    .Y(_03930_));
 sky130_fd_sc_hd__nand3_1 _05493_ (.A(_03523_),
    .B(_03567_),
    .C(_03930_),
    .Y(_03941_));
 sky130_fd_sc_hd__nand2_1 _05494_ (.A(_03919_),
    .B(_03941_),
    .Y(_03952_));
 sky130_fd_sc_hd__inv_2 _05495_ (.A(_03952_),
    .Y(_03963_));
 sky130_fd_sc_hd__nor2_1 _05496_ (.A(_02951_),
    .B(_02214_),
    .Y(_03974_));
 sky130_fd_sc_hd__a21oi_2 _05497_ (.A1(_02962_),
    .A2(_03963_),
    .B1(_03974_),
    .Y(_03985_));
 sky130_fd_sc_hd__nand2_1 _05498_ (.A(_01741_),
    .B(_01268_),
    .Y(_03996_));
 sky130_fd_sc_hd__inv_2 _05499_ (.A(_03996_),
    .Y(_04007_));
 sky130_fd_sc_hd__nor2_1 _05500_ (.A(_01268_),
    .B(_01741_),
    .Y(_04018_));
 sky130_fd_sc_hd__o21bai_1 _05501_ (.A1(_02170_),
    .A2(_04007_),
    .B1_N(_04018_),
    .Y(_04029_));
 sky130_fd_sc_hd__nand2_1 _05502_ (.A(_01642_),
    .B(_01444_),
    .Y(_04040_));
 sky130_fd_sc_hd__nor2_1 _05503_ (.A(_01301_),
    .B(_01334_),
    .Y(_04051_));
 sky130_fd_sc_hd__a21oi_2 _05504_ (.A1(_01389_),
    .A2(_01378_),
    .B1(_04051_),
    .Y(_04062_));
 sky130_fd_sc_hd__inv_2 _05505_ (.A(_04062_),
    .Y(_04073_));
 sky130_fd_sc_hd__buf_4 _05506_ (.A(net14),
    .X(_04084_));
 sky130_fd_sc_hd__nand2_1 _05507_ (.A(_02379_),
    .B(_04084_),
    .Y(_04095_));
 sky130_fd_sc_hd__inv_2 _05508_ (.A(_04095_),
    .Y(_04106_));
 sky130_fd_sc_hd__nand2_1 _05509_ (.A(_01323_),
    .B(_00751_),
    .Y(_04117_));
 sky130_fd_sc_hd__inv_2 _05510_ (.A(_04117_),
    .Y(_04128_));
 sky130_fd_sc_hd__nand2_1 _05511_ (.A(_04106_),
    .B(_04128_),
    .Y(_04139_));
 sky130_fd_sc_hd__nand2_1 _05512_ (.A(_00784_),
    .B(_00861_),
    .Y(_04150_));
 sky130_fd_sc_hd__inv_2 _05513_ (.A(_04150_),
    .Y(_04161_));
 sky130_fd_sc_hd__nand2_1 _05514_ (.A(_04095_),
    .B(_04117_),
    .Y(_04172_));
 sky130_fd_sc_hd__nand3_1 _05515_ (.A(_04139_),
    .B(_04161_),
    .C(_04172_),
    .Y(_04183_));
 sky130_fd_sc_hd__nand2_1 _05516_ (.A(_04128_),
    .B(_04095_),
    .Y(_04194_));
 sky130_fd_sc_hd__nand2_1 _05517_ (.A(_04106_),
    .B(_04117_),
    .Y(_04205_));
 sky130_fd_sc_hd__nand3_1 _05518_ (.A(_04194_),
    .B(_04205_),
    .C(_04150_),
    .Y(_04216_));
 sky130_fd_sc_hd__nand3_1 _05519_ (.A(_04073_),
    .B(_04183_),
    .C(_04216_),
    .Y(_04227_));
 sky130_fd_sc_hd__nand2_1 _05520_ (.A(_04216_),
    .B(_04183_),
    .Y(_04238_));
 sky130_fd_sc_hd__nand2_1 _05521_ (.A(_04238_),
    .B(_04062_),
    .Y(_04249_));
 sky130_fd_sc_hd__buf_8 _05522_ (.A(_01048_),
    .X(_04260_));
 sky130_fd_sc_hd__nand2_1 _05523_ (.A(_00850_),
    .B(_04260_),
    .Y(_04271_));
 sky130_fd_sc_hd__inv_2 _05524_ (.A(_04271_),
    .Y(_04282_));
 sky130_fd_sc_hd__buf_8 _05525_ (.A(_01092_),
    .X(_04293_));
 sky130_fd_sc_hd__nand2_1 _05526_ (.A(_00740_),
    .B(_04293_),
    .Y(_04304_));
 sky130_fd_sc_hd__inv_2 _05527_ (.A(_04304_),
    .Y(_04315_));
 sky130_fd_sc_hd__nand2_1 _05528_ (.A(_04282_),
    .B(_04315_),
    .Y(_04326_));
 sky130_fd_sc_hd__nand2_1 _05529_ (.A(_04271_),
    .B(_04304_),
    .Y(_04337_));
 sky130_fd_sc_hd__nand2_1 _05530_ (.A(_04326_),
    .B(_04337_),
    .Y(_04348_));
 sky130_fd_sc_hd__nand2_1 _05531_ (.A(_01081_),
    .B(_01158_),
    .Y(_04359_));
 sky130_fd_sc_hd__nand2_1 _05532_ (.A(_04348_),
    .B(_04359_),
    .Y(_04370_));
 sky130_fd_sc_hd__inv_2 _05533_ (.A(_04359_),
    .Y(_04381_));
 sky130_fd_sc_hd__nand3_1 _05534_ (.A(_04326_),
    .B(_04381_),
    .C(_04337_),
    .Y(_04392_));
 sky130_fd_sc_hd__nand2_1 _05535_ (.A(_04370_),
    .B(_04392_),
    .Y(_04403_));
 sky130_fd_sc_hd__inv_2 _05536_ (.A(_04403_),
    .Y(_04414_));
 sky130_fd_sc_hd__nand3_2 _05537_ (.A(_04227_),
    .B(_04249_),
    .C(_04414_),
    .Y(_04425_));
 sky130_fd_sc_hd__nand2_1 _05538_ (.A(_04238_),
    .B(_04073_),
    .Y(_04436_));
 sky130_fd_sc_hd__nand3_1 _05539_ (.A(_04062_),
    .B(_04216_),
    .C(_04183_),
    .Y(_04447_));
 sky130_fd_sc_hd__nand3_1 _05540_ (.A(_04436_),
    .B(_04447_),
    .C(_04403_),
    .Y(_04458_));
 sky130_fd_sc_hd__nand3_1 _05541_ (.A(_04040_),
    .B(_04425_),
    .C(_04458_),
    .Y(_04469_));
 sky130_fd_sc_hd__nand2_1 _05542_ (.A(_01147_),
    .B(_01774_),
    .Y(_04480_));
 sky130_fd_sc_hd__inv_2 _05543_ (.A(_04480_),
    .Y(_04490_));
 sky130_fd_sc_hd__nand2_1 _05544_ (.A(net7),
    .B(_01807_),
    .Y(_04500_));
 sky130_fd_sc_hd__inv_2 _05545_ (.A(_04500_),
    .Y(_04510_));
 sky130_fd_sc_hd__nand2_1 _05546_ (.A(_04490_),
    .B(_04510_),
    .Y(_04520_));
 sky130_fd_sc_hd__nand2_1 _05547_ (.A(_04480_),
    .B(_04500_),
    .Y(_04529_));
 sky130_fd_sc_hd__nand2_1 _05548_ (.A(_04520_),
    .B(_04529_),
    .Y(_04539_));
 sky130_fd_sc_hd__nand2_1 _05549_ (.A(_02544_),
    .B(_01884_),
    .Y(_04549_));
 sky130_fd_sc_hd__nand2_1 _05550_ (.A(_04539_),
    .B(_04549_),
    .Y(_04558_));
 sky130_fd_sc_hd__inv_2 _05551_ (.A(_04549_),
    .Y(_04568_));
 sky130_fd_sc_hd__nand3_2 _05552_ (.A(_04520_),
    .B(_04568_),
    .C(_04529_),
    .Y(_04578_));
 sky130_fd_sc_hd__nand2_1 _05553_ (.A(_04558_),
    .B(_04578_),
    .Y(_04588_));
 sky130_fd_sc_hd__nor2_1 _05554_ (.A(_01488_),
    .B(_01510_),
    .Y(_04598_));
 sky130_fd_sc_hd__a21oi_2 _05555_ (.A1(_01543_),
    .A2(_01598_),
    .B1(_04598_),
    .Y(_04607_));
 sky130_fd_sc_hd__nand2_1 _05556_ (.A(_04588_),
    .B(_04607_),
    .Y(_04617_));
 sky130_fd_sc_hd__a21o_1 _05557_ (.A1(_01543_),
    .A2(_01598_),
    .B1(_04598_),
    .X(_04627_));
 sky130_fd_sc_hd__nand3_1 _05558_ (.A(_04627_),
    .B(_04578_),
    .C(_04558_),
    .Y(_04636_));
 sky130_fd_sc_hd__nand2_2 _05559_ (.A(_01917_),
    .B(_01840_),
    .Y(_04646_));
 sky130_fd_sc_hd__nand3_1 _05560_ (.A(_04617_),
    .B(_04636_),
    .C(_04646_),
    .Y(_04655_));
 sky130_fd_sc_hd__nand2_1 _05561_ (.A(_04588_),
    .B(_04627_),
    .Y(_04663_));
 sky130_fd_sc_hd__nand3_1 _05562_ (.A(_04558_),
    .B(_04607_),
    .C(_04578_),
    .Y(_04672_));
 sky130_fd_sc_hd__inv_2 _05563_ (.A(_04646_),
    .Y(_04680_));
 sky130_fd_sc_hd__nand3_1 _05564_ (.A(_04663_),
    .B(_04672_),
    .C(_04680_),
    .Y(_04689_));
 sky130_fd_sc_hd__nand2_1 _05565_ (.A(_04655_),
    .B(_04689_),
    .Y(_04696_));
 sky130_fd_sc_hd__inv_2 _05566_ (.A(_04696_),
    .Y(_04704_));
 sky130_fd_sc_hd__nand2_1 _05567_ (.A(_04425_),
    .B(_04458_),
    .Y(_04712_));
 sky130_fd_sc_hd__nor2_1 _05568_ (.A(_01466_),
    .B(_01455_),
    .Y(_04721_));
 sky130_fd_sc_hd__a21oi_2 _05569_ (.A1(_01477_),
    .A2(_01631_),
    .B1(_04721_),
    .Y(_04730_));
 sky130_fd_sc_hd__nand2_1 _05570_ (.A(_04712_),
    .B(_04730_),
    .Y(_04738_));
 sky130_fd_sc_hd__nand3_1 _05571_ (.A(_04469_),
    .B(_04704_),
    .C(_04738_),
    .Y(_04744_));
 sky130_fd_sc_hd__nand3_1 _05572_ (.A(_04730_),
    .B(_04425_),
    .C(_04458_),
    .Y(_04745_));
 sky130_fd_sc_hd__nand2_1 _05573_ (.A(_04712_),
    .B(_04040_),
    .Y(_04746_));
 sky130_fd_sc_hd__nand3_1 _05574_ (.A(_04745_),
    .B(_04746_),
    .C(_04696_),
    .Y(_04747_));
 sky130_fd_sc_hd__nand3_1 _05575_ (.A(_04029_),
    .B(_04744_),
    .C(_04747_),
    .Y(_04748_));
 sky130_fd_sc_hd__nor2_1 _05576_ (.A(_01950_),
    .B(_01928_),
    .Y(_04749_));
 sky130_fd_sc_hd__a21oi_2 _05577_ (.A1(_01961_),
    .A2(_02104_),
    .B1(_04749_),
    .Y(_04750_));
 sky130_fd_sc_hd__nand2_1 _05578_ (.A(net3),
    .B(_02995_),
    .Y(_04751_));
 sky130_fd_sc_hd__inv_2 _05579_ (.A(_04751_),
    .Y(_04752_));
 sky130_fd_sc_hd__nand2_1 _05580_ (.A(net4),
    .B(_03028_),
    .Y(_04753_));
 sky130_fd_sc_hd__inv_2 _05581_ (.A(_04753_),
    .Y(_04754_));
 sky130_fd_sc_hd__nand2_1 _05582_ (.A(_04752_),
    .B(_04754_),
    .Y(_04755_));
 sky130_fd_sc_hd__nand2_1 _05583_ (.A(_04751_),
    .B(_04753_),
    .Y(_04756_));
 sky130_fd_sc_hd__nand2_1 _05584_ (.A(_04755_),
    .B(_04756_),
    .Y(_04757_));
 sky130_fd_sc_hd__nand2_1 _05585_ (.A(net35),
    .B(_02753_),
    .Y(_04758_));
 sky130_fd_sc_hd__nand2_1 _05586_ (.A(_04757_),
    .B(_04758_),
    .Y(_04759_));
 sky130_fd_sc_hd__inv_2 _05587_ (.A(_04758_),
    .Y(_04760_));
 sky130_fd_sc_hd__nand3_1 _05588_ (.A(_04755_),
    .B(_04760_),
    .C(_04756_),
    .Y(_04761_));
 sky130_fd_sc_hd__nand2_1 _05589_ (.A(_04759_),
    .B(_04761_),
    .Y(_04762_));
 sky130_fd_sc_hd__nor2_1 _05590_ (.A(_03006_),
    .B(_03039_),
    .Y(_04763_));
 sky130_fd_sc_hd__a21oi_1 _05591_ (.A1(_03072_),
    .A2(_03127_),
    .B1(_04763_),
    .Y(_04764_));
 sky130_fd_sc_hd__nand2_1 _05592_ (.A(_04762_),
    .B(_04764_),
    .Y(_04765_));
 sky130_fd_sc_hd__a21o_1 _05593_ (.A1(_03072_),
    .A2(_03127_),
    .B1(_04763_),
    .X(_04766_));
 sky130_fd_sc_hd__nand3_1 _05594_ (.A(_04766_),
    .B(_04761_),
    .C(_04759_),
    .Y(_04767_));
 sky130_fd_sc_hd__nand2_1 _05595_ (.A(net37),
    .B(_03226_),
    .Y(_04768_));
 sky130_fd_sc_hd__inv_2 _05596_ (.A(_04768_),
    .Y(_04769_));
 sky130_fd_sc_hd__nand2_1 _05597_ (.A(net36),
    .B(_03094_),
    .Y(_04770_));
 sky130_fd_sc_hd__inv_2 _05598_ (.A(_04770_),
    .Y(_04771_));
 sky130_fd_sc_hd__nand2_1 _05599_ (.A(_04769_),
    .B(_04771_),
    .Y(_04772_));
 sky130_fd_sc_hd__nand2_1 _05600_ (.A(_04768_),
    .B(_04770_),
    .Y(_04773_));
 sky130_fd_sc_hd__nand2_1 _05601_ (.A(_04772_),
    .B(_04773_),
    .Y(_04774_));
 sky130_fd_sc_hd__nand2_1 _05602_ (.A(net38),
    .B(_03314_),
    .Y(_04775_));
 sky130_fd_sc_hd__nand2_1 _05603_ (.A(_04774_),
    .B(_04775_),
    .Y(_04776_));
 sky130_fd_sc_hd__inv_2 _05604_ (.A(_04775_),
    .Y(_04777_));
 sky130_fd_sc_hd__nand3_1 _05605_ (.A(_04772_),
    .B(_04777_),
    .C(_04773_),
    .Y(_04778_));
 sky130_fd_sc_hd__nand2_1 _05606_ (.A(_04776_),
    .B(_04778_),
    .Y(_04779_));
 sky130_fd_sc_hd__inv_2 _05607_ (.A(_04779_),
    .Y(_04780_));
 sky130_fd_sc_hd__nand3_1 _05608_ (.A(_04765_),
    .B(_04767_),
    .C(_04780_),
    .Y(_04781_));
 sky130_fd_sc_hd__nand2_1 _05609_ (.A(_04762_),
    .B(_04766_),
    .Y(_04782_));
 sky130_fd_sc_hd__nand3_1 _05610_ (.A(_04759_),
    .B(_04764_),
    .C(_04761_),
    .Y(_04783_));
 sky130_fd_sc_hd__nand3_1 _05611_ (.A(_04782_),
    .B(_04783_),
    .C(_04779_),
    .Y(_04784_));
 sky130_fd_sc_hd__nand3_1 _05612_ (.A(_04750_),
    .B(_04781_),
    .C(_04784_),
    .Y(_04785_));
 sky130_fd_sc_hd__nand2_1 _05613_ (.A(_04781_),
    .B(_04784_),
    .Y(_04786_));
 sky130_fd_sc_hd__nand2_1 _05614_ (.A(_02115_),
    .B(_01983_),
    .Y(_04787_));
 sky130_fd_sc_hd__nand2_1 _05615_ (.A(_04786_),
    .B(_04787_),
    .Y(_04788_));
 sky130_fd_sc_hd__nand2_1 _05616_ (.A(_04785_),
    .B(_04788_),
    .Y(_04789_));
 sky130_fd_sc_hd__nand2_2 _05617_ (.A(_03479_),
    .B(_03303_),
    .Y(_04790_));
 sky130_fd_sc_hd__nand2_1 _05618_ (.A(_04789_),
    .B(_04790_),
    .Y(_04791_));
 sky130_fd_sc_hd__inv_2 _05619_ (.A(_04790_),
    .Y(_04792_));
 sky130_fd_sc_hd__nand3_1 _05620_ (.A(_04785_),
    .B(_04788_),
    .C(_04792_),
    .Y(_04793_));
 sky130_fd_sc_hd__nand2_1 _05621_ (.A(_04791_),
    .B(_04793_),
    .Y(_04794_));
 sky130_fd_sc_hd__inv_2 _05622_ (.A(_04794_),
    .Y(_04795_));
 sky130_fd_sc_hd__nand2_1 _05623_ (.A(_04744_),
    .B(_04747_),
    .Y(_04796_));
 sky130_fd_sc_hd__a21oi_1 _05624_ (.A1(_03996_),
    .A2(_02181_),
    .B1(_04018_),
    .Y(_04797_));
 sky130_fd_sc_hd__nand2_1 _05625_ (.A(_04796_),
    .B(_04797_),
    .Y(_04798_));
 sky130_fd_sc_hd__nand3_1 _05626_ (.A(_04748_),
    .B(_04795_),
    .C(_04798_),
    .Y(_04799_));
 sky130_fd_sc_hd__nand2_1 _05627_ (.A(_04796_),
    .B(_04029_),
    .Y(_04800_));
 sky130_fd_sc_hd__nand3_1 _05628_ (.A(_04797_),
    .B(_04744_),
    .C(_04747_),
    .Y(_04801_));
 sky130_fd_sc_hd__nand3_1 _05629_ (.A(_04800_),
    .B(_04801_),
    .C(_04794_),
    .Y(_04802_));
 sky130_fd_sc_hd__nand3_1 _05630_ (.A(_03985_),
    .B(_04799_),
    .C(_04802_),
    .Y(_04803_));
 sky130_fd_sc_hd__nand2_1 _05631_ (.A(_04799_),
    .B(_04802_),
    .Y(_04804_));
 sky130_fd_sc_hd__a21o_1 _05632_ (.A1(_02962_),
    .A2(_03963_),
    .B1(_03974_),
    .X(_04805_));
 sky130_fd_sc_hd__nand2_1 _05633_ (.A(_04804_),
    .B(_04805_),
    .Y(_04806_));
 sky130_fd_sc_hd__nand2_1 _05634_ (.A(_04803_),
    .B(_04806_),
    .Y(_04807_));
 sky130_fd_sc_hd__clkbuf_8 _05635_ (.A(net40),
    .X(_04808_));
 sky130_fd_sc_hd__buf_6 _05636_ (.A(net27),
    .X(_04809_));
 sky130_fd_sc_hd__nand2_1 _05637_ (.A(_04808_),
    .B(_04809_),
    .Y(_04810_));
 sky130_fd_sc_hd__inv_2 _05638_ (.A(_04810_),
    .Y(_04811_));
 sky130_fd_sc_hd__clkbuf_8 _05639_ (.A(net39),
    .X(_04812_));
 sky130_fd_sc_hd__nand2_1 _05640_ (.A(_04812_),
    .B(_03820_),
    .Y(_04813_));
 sky130_fd_sc_hd__inv_2 _05641_ (.A(_04813_),
    .Y(_04814_));
 sky130_fd_sc_hd__nand2_1 _05642_ (.A(_04811_),
    .B(_04814_),
    .Y(_04815_));
 sky130_fd_sc_hd__nand2_1 _05643_ (.A(_04810_),
    .B(_04813_),
    .Y(_04816_));
 sky130_fd_sc_hd__nand2_1 _05644_ (.A(_04815_),
    .B(_04816_),
    .Y(_04817_));
 sky130_fd_sc_hd__clkbuf_8 _05645_ (.A(net41),
    .X(_04818_));
 sky130_fd_sc_hd__buf_6 _05646_ (.A(net26),
    .X(_04819_));
 sky130_fd_sc_hd__nand2_1 _05647_ (.A(_04818_),
    .B(_04819_),
    .Y(_04820_));
 sky130_fd_sc_hd__nand2_1 _05648_ (.A(_04817_),
    .B(_04820_),
    .Y(_04821_));
 sky130_fd_sc_hd__inv_2 _05649_ (.A(_04820_),
    .Y(_04822_));
 sky130_fd_sc_hd__nand3_2 _05650_ (.A(_04815_),
    .B(_04822_),
    .C(_04816_),
    .Y(_04823_));
 sky130_fd_sc_hd__nand2_1 _05651_ (.A(_04821_),
    .B(_04823_),
    .Y(_04824_));
 sky130_fd_sc_hd__a21oi_1 _05652_ (.A1(_03787_),
    .A2(_03853_),
    .B1(_03776_),
    .Y(_04825_));
 sky130_fd_sc_hd__nand2_1 _05653_ (.A(_04824_),
    .B(_04825_),
    .Y(_04826_));
 sky130_fd_sc_hd__clkbuf_8 _05654_ (.A(net23),
    .X(_04827_));
 sky130_fd_sc_hd__clkbuf_8 _05655_ (.A(_04827_),
    .X(_04828_));
 sky130_fd_sc_hd__nand2_1 _05656_ (.A(_04818_),
    .B(_04828_),
    .Y(_04829_));
 sky130_fd_sc_hd__nand2_1 _05657_ (.A(_04812_),
    .B(_04809_),
    .Y(_04830_));
 sky130_fd_sc_hd__inv_2 _05658_ (.A(_04830_),
    .Y(_04831_));
 sky130_fd_sc_hd__nand2_1 _05659_ (.A(_04808_),
    .B(_04819_),
    .Y(_04832_));
 sky130_fd_sc_hd__inv_2 _05660_ (.A(_04832_),
    .Y(_04833_));
 sky130_fd_sc_hd__nand2_1 _05661_ (.A(_04831_),
    .B(_04833_),
    .Y(_04834_));
 sky130_fd_sc_hd__nand2_1 _05662_ (.A(_04830_),
    .B(_04832_),
    .Y(_04835_));
 sky130_fd_sc_hd__nand3b_1 _05663_ (.A_N(_04829_),
    .B(_04834_),
    .C(_04835_),
    .Y(_04836_));
 sky130_fd_sc_hd__nand2_1 _05664_ (.A(_04836_),
    .B(_04834_),
    .Y(_04837_));
 sky130_fd_sc_hd__nor2_1 _05665_ (.A(_04825_),
    .B(_04824_),
    .Y(_04838_));
 sky130_fd_sc_hd__a21oi_1 _05666_ (.A1(_04826_),
    .A2(_04837_),
    .B1(_04838_),
    .Y(_04839_));
 sky130_fd_sc_hd__nand2_1 _05667_ (.A(net40),
    .B(_03820_),
    .Y(_04840_));
 sky130_fd_sc_hd__inv_2 _05668_ (.A(_04840_),
    .Y(_04841_));
 sky130_fd_sc_hd__nand2_1 _05669_ (.A(net39),
    .B(_03402_),
    .Y(_04842_));
 sky130_fd_sc_hd__inv_2 _05670_ (.A(_04842_),
    .Y(_04843_));
 sky130_fd_sc_hd__nand2_1 _05671_ (.A(_04841_),
    .B(_04843_),
    .Y(_04844_));
 sky130_fd_sc_hd__nand2_1 _05672_ (.A(_04840_),
    .B(_04842_),
    .Y(_04845_));
 sky130_fd_sc_hd__nand2_1 _05673_ (.A(_04844_),
    .B(_04845_),
    .Y(_04846_));
 sky130_fd_sc_hd__nand2_1 _05674_ (.A(_04818_),
    .B(_04809_),
    .Y(_04847_));
 sky130_fd_sc_hd__nand2_1 _05675_ (.A(_04846_),
    .B(_04847_),
    .Y(_04848_));
 sky130_fd_sc_hd__nand3b_2 _05676_ (.A_N(_04847_),
    .B(_04844_),
    .C(_04845_),
    .Y(_04849_));
 sky130_fd_sc_hd__nand2_1 _05677_ (.A(_04848_),
    .B(_04849_),
    .Y(_04850_));
 sky130_fd_sc_hd__nor2_1 _05678_ (.A(_03325_),
    .B(_03347_),
    .Y(_04851_));
 sky130_fd_sc_hd__a21oi_1 _05679_ (.A1(_03380_),
    .A2(_03435_),
    .B1(_04851_),
    .Y(_04852_));
 sky130_fd_sc_hd__nand2_1 _05680_ (.A(_04850_),
    .B(_04852_),
    .Y(_04853_));
 sky130_fd_sc_hd__a21o_1 _05681_ (.A1(_03380_),
    .A2(_03435_),
    .B1(_04851_),
    .X(_04854_));
 sky130_fd_sc_hd__nand3_1 _05682_ (.A(_04854_),
    .B(_04849_),
    .C(_04848_),
    .Y(_04855_));
 sky130_fd_sc_hd__nand2_1 _05683_ (.A(_04823_),
    .B(_04815_),
    .Y(_04856_));
 sky130_fd_sc_hd__nand3_1 _05684_ (.A(_04853_),
    .B(_04855_),
    .C(_04856_),
    .Y(_04857_));
 sky130_fd_sc_hd__nand2_1 _05685_ (.A(_04850_),
    .B(_04854_),
    .Y(_04858_));
 sky130_fd_sc_hd__nand3_1 _05686_ (.A(_04848_),
    .B(_04849_),
    .C(_04852_),
    .Y(_04859_));
 sky130_fd_sc_hd__inv_2 _05687_ (.A(_04856_),
    .Y(_04860_));
 sky130_fd_sc_hd__nand3_1 _05688_ (.A(_04858_),
    .B(_04859_),
    .C(_04860_),
    .Y(_04861_));
 sky130_fd_sc_hd__nand3_1 _05689_ (.A(_04839_),
    .B(_04857_),
    .C(_04861_),
    .Y(_04862_));
 sky130_fd_sc_hd__nand2_1 _05690_ (.A(_04857_),
    .B(_04861_),
    .Y(_04863_));
 sky130_fd_sc_hd__inv_2 _05691_ (.A(_04837_),
    .Y(_04864_));
 sky130_fd_sc_hd__a21o_1 _05692_ (.A1(_03787_),
    .A2(_03853_),
    .B1(_03776_),
    .X(_04865_));
 sky130_fd_sc_hd__a21oi_1 _05693_ (.A1(_04821_),
    .A2(_04823_),
    .B1(_04865_),
    .Y(_04866_));
 sky130_fd_sc_hd__nand3_1 _05694_ (.A(_04865_),
    .B(_04823_),
    .C(_04821_),
    .Y(_04867_));
 sky130_fd_sc_hd__o21ai_1 _05695_ (.A1(_04864_),
    .A2(_04866_),
    .B1(_04867_),
    .Y(_04868_));
 sky130_fd_sc_hd__nand2_1 _05696_ (.A(_04863_),
    .B(_04868_),
    .Y(_04869_));
 sky130_fd_sc_hd__nand2_1 _05697_ (.A(_04862_),
    .B(_04869_),
    .Y(_04870_));
 sky130_fd_sc_hd__buf_4 _05698_ (.A(net43),
    .X(_04871_));
 sky130_fd_sc_hd__nand2_1 _05699_ (.A(_04871_),
    .B(net12),
    .Y(_04872_));
 sky130_fd_sc_hd__buf_4 _05700_ (.A(net42),
    .X(_04873_));
 sky130_fd_sc_hd__nand2_1 _05701_ (.A(_04873_),
    .B(_04827_),
    .Y(_04874_));
 sky130_fd_sc_hd__nand2_1 _05702_ (.A(_04872_),
    .B(_04874_),
    .Y(_04875_));
 sky130_fd_sc_hd__buf_4 _05703_ (.A(net45),
    .X(_04876_));
 sky130_fd_sc_hd__nand2_1 _05704_ (.A(_04876_),
    .B(net1),
    .Y(_04877_));
 sky130_fd_sc_hd__inv_2 _05705_ (.A(_04877_),
    .Y(_04878_));
 sky130_fd_sc_hd__nor2_1 _05706_ (.A(_04872_),
    .B(_04874_),
    .Y(_04879_));
 sky130_fd_sc_hd__a21oi_1 _05707_ (.A1(_04875_),
    .A2(_04878_),
    .B1(_04879_),
    .Y(_04880_));
 sky130_fd_sc_hd__nand2_1 _05708_ (.A(_04871_),
    .B(_04827_),
    .Y(_04881_));
 sky130_fd_sc_hd__nand2_1 _05709_ (.A(_04873_),
    .B(_04819_),
    .Y(_04882_));
 sky130_fd_sc_hd__nor2_1 _05710_ (.A(_04881_),
    .B(_04882_),
    .Y(_04883_));
 sky130_fd_sc_hd__inv_2 _05711_ (.A(_04883_),
    .Y(_04884_));
 sky130_fd_sc_hd__nand2_1 _05712_ (.A(_04881_),
    .B(_04882_),
    .Y(_04885_));
 sky130_fd_sc_hd__nand2_1 _05713_ (.A(_04884_),
    .B(_04885_),
    .Y(_04886_));
 sky130_fd_sc_hd__nand2_1 _05714_ (.A(_04876_),
    .B(net12),
    .Y(_04887_));
 sky130_fd_sc_hd__nand2_1 _05715_ (.A(_04886_),
    .B(_04887_),
    .Y(_04888_));
 sky130_fd_sc_hd__inv_2 _05716_ (.A(_04887_),
    .Y(_04889_));
 sky130_fd_sc_hd__nand3_1 _05717_ (.A(_04884_),
    .B(_04885_),
    .C(_04889_),
    .Y(_04890_));
 sky130_fd_sc_hd__nand3b_1 _05718_ (.A_N(_04880_),
    .B(_04888_),
    .C(_04890_),
    .Y(_04891_));
 sky130_fd_sc_hd__nand2_1 _05719_ (.A(_04888_),
    .B(_04890_),
    .Y(_04892_));
 sky130_fd_sc_hd__nand2_1 _05720_ (.A(_04892_),
    .B(_04880_),
    .Y(_04893_));
 sky130_fd_sc_hd__nand2_1 _05721_ (.A(_04891_),
    .B(_04893_),
    .Y(_04894_));
 sky130_fd_sc_hd__clkbuf_8 _05722_ (.A(net1),
    .X(_04895_));
 sky130_fd_sc_hd__nand2_1 _05723_ (.A(net46),
    .B(_04895_),
    .Y(_04896_));
 sky130_fd_sc_hd__nand2_1 _05724_ (.A(_04894_),
    .B(_04896_),
    .Y(_04897_));
 sky130_fd_sc_hd__nand3b_1 _05725_ (.A_N(_04896_),
    .B(_04891_),
    .C(_04893_),
    .Y(_04898_));
 sky130_fd_sc_hd__nand2_1 _05726_ (.A(_04897_),
    .B(_04898_),
    .Y(_04899_));
 sky130_fd_sc_hd__inv_2 _05727_ (.A(_04899_),
    .Y(_04900_));
 sky130_fd_sc_hd__nand2_1 _05728_ (.A(_04870_),
    .B(_04900_),
    .Y(_04901_));
 sky130_fd_sc_hd__nand3_1 _05729_ (.A(_04862_),
    .B(_04869_),
    .C(_04899_),
    .Y(_04902_));
 sky130_fd_sc_hd__nand2_1 _05730_ (.A(_04901_),
    .B(_04902_),
    .Y(_04903_));
 sky130_fd_sc_hd__nand2_1 _05731_ (.A(_03534_),
    .B(_02984_),
    .Y(_04904_));
 sky130_fd_sc_hd__nor2_1 _05732_ (.A(_02984_),
    .B(_03534_),
    .Y(_04905_));
 sky130_fd_sc_hd__a21oi_2 _05733_ (.A1(_04904_),
    .A2(_03908_),
    .B1(_04905_),
    .Y(_04906_));
 sky130_fd_sc_hd__inv_2 _05734_ (.A(_04906_),
    .Y(_04907_));
 sky130_fd_sc_hd__nand2_1 _05735_ (.A(_04903_),
    .B(_04907_),
    .Y(_04908_));
 sky130_fd_sc_hd__nand3_1 _05736_ (.A(_04906_),
    .B(_04901_),
    .C(_04902_),
    .Y(_04909_));
 sky130_fd_sc_hd__nand2_1 _05737_ (.A(_04908_),
    .B(_04909_),
    .Y(_04910_));
 sky130_fd_sc_hd__clkbuf_8 _05738_ (.A(net12),
    .X(_04911_));
 sky130_fd_sc_hd__and4_1 _05739_ (.A(_04873_),
    .B(_04871_),
    .C(_04911_),
    .D(net1),
    .X(_04912_));
 sky130_fd_sc_hd__inv_2 _05740_ (.A(_04912_),
    .Y(_04913_));
 sky130_fd_sc_hd__nor2b_1 _05741_ (.A(_04879_),
    .B_N(_04875_),
    .Y(_04914_));
 sky130_fd_sc_hd__xor2_1 _05742_ (.A(_04877_),
    .B(_04914_),
    .X(_04915_));
 sky130_fd_sc_hd__or2_2 _05743_ (.A(_04913_),
    .B(_04915_),
    .X(_04916_));
 sky130_fd_sc_hd__nand2_1 _05744_ (.A(_04915_),
    .B(_04913_),
    .Y(_04917_));
 sky130_fd_sc_hd__nand2_1 _05745_ (.A(_04916_),
    .B(_04917_),
    .Y(_04918_));
 sky130_fd_sc_hd__inv_2 _05746_ (.A(_04918_),
    .Y(_04919_));
 sky130_fd_sc_hd__nand2_1 _05747_ (.A(_04826_),
    .B(_04867_),
    .Y(_04920_));
 sky130_fd_sc_hd__nand2_1 _05748_ (.A(_04920_),
    .B(_04864_),
    .Y(_04921_));
 sky130_fd_sc_hd__nand3_1 _05749_ (.A(_04826_),
    .B(_04867_),
    .C(_04837_),
    .Y(_04922_));
 sky130_fd_sc_hd__nand2_1 _05750_ (.A(_04921_),
    .B(_04922_),
    .Y(_04923_));
 sky130_fd_sc_hd__nand2_1 _05751_ (.A(_04834_),
    .B(_04835_),
    .Y(_04924_));
 sky130_fd_sc_hd__nand2_1 _05752_ (.A(_04924_),
    .B(_04829_),
    .Y(_04925_));
 sky130_fd_sc_hd__nand2_1 _05753_ (.A(_04925_),
    .B(_04836_),
    .Y(_04926_));
 sky130_fd_sc_hd__nand2_1 _05754_ (.A(net37),
    .B(_03820_),
    .Y(_04927_));
 sky130_fd_sc_hd__clkbuf_8 _05755_ (.A(_03402_),
    .X(_04928_));
 sky130_fd_sc_hd__nand2_1 _05756_ (.A(net36),
    .B(_04928_),
    .Y(_04929_));
 sky130_fd_sc_hd__nand2_1 _05757_ (.A(_04927_),
    .B(_04929_),
    .Y(_04930_));
 sky130_fd_sc_hd__nand2_1 _05758_ (.A(net38),
    .B(_04809_),
    .Y(_04931_));
 sky130_fd_sc_hd__inv_2 _05759_ (.A(_04931_),
    .Y(_04932_));
 sky130_fd_sc_hd__nor2_1 _05760_ (.A(_04927_),
    .B(_04929_),
    .Y(_04933_));
 sky130_fd_sc_hd__a21oi_2 _05761_ (.A1(_04930_),
    .A2(_04932_),
    .B1(_04933_),
    .Y(_04934_));
 sky130_fd_sc_hd__nand2_1 _05762_ (.A(_04926_),
    .B(_04934_),
    .Y(_04935_));
 sky130_fd_sc_hd__nand2_1 _05763_ (.A(_04808_),
    .B(_04827_),
    .Y(_04936_));
 sky130_fd_sc_hd__nand2_1 _05764_ (.A(_04812_),
    .B(_04819_),
    .Y(_04937_));
 sky130_fd_sc_hd__nand2b_1 _05765_ (.A_N(_04936_),
    .B(_04937_),
    .Y(_04938_));
 sky130_fd_sc_hd__nand2b_1 _05766_ (.A_N(_04937_),
    .B(_04936_),
    .Y(_04939_));
 sky130_fd_sc_hd__nand2_1 _05767_ (.A(_04938_),
    .B(_04939_),
    .Y(_04940_));
 sky130_fd_sc_hd__nand2_1 _05768_ (.A(_04818_),
    .B(_04911_),
    .Y(_04941_));
 sky130_fd_sc_hd__inv_2 _05769_ (.A(_04941_),
    .Y(_04942_));
 sky130_fd_sc_hd__nand2_1 _05770_ (.A(_04940_),
    .B(_04942_),
    .Y(_04943_));
 sky130_fd_sc_hd__o21ai_2 _05771_ (.A1(_04936_),
    .A2(_04937_),
    .B1(_04943_),
    .Y(_04944_));
 sky130_fd_sc_hd__inv_2 _05772_ (.A(_04934_),
    .Y(_04945_));
 sky130_fd_sc_hd__nand3_1 _05773_ (.A(_04945_),
    .B(_04836_),
    .C(_04925_),
    .Y(_04946_));
 sky130_fd_sc_hd__inv_2 _05774_ (.A(_04946_),
    .Y(_04947_));
 sky130_fd_sc_hd__a21oi_2 _05775_ (.A1(_04935_),
    .A2(_04944_),
    .B1(_04947_),
    .Y(_04948_));
 sky130_fd_sc_hd__nand2_1 _05776_ (.A(_04923_),
    .B(_04948_),
    .Y(_04949_));
 sky130_fd_sc_hd__nor2_1 _05777_ (.A(_04948_),
    .B(_04923_),
    .Y(_04950_));
 sky130_fd_sc_hd__a21oi_1 _05778_ (.A1(_04919_),
    .A2(_04949_),
    .B1(_04950_),
    .Y(_04951_));
 sky130_fd_sc_hd__inv_2 _05779_ (.A(_04951_),
    .Y(_04952_));
 sky130_fd_sc_hd__nand2_1 _05780_ (.A(_04910_),
    .B(_04952_),
    .Y(_04953_));
 sky130_fd_sc_hd__nand3_1 _05781_ (.A(_04908_),
    .B(_04909_),
    .C(_04951_),
    .Y(_04954_));
 sky130_fd_sc_hd__nand2_1 _05782_ (.A(_04953_),
    .B(_04954_),
    .Y(_04955_));
 sky130_fd_sc_hd__inv_2 _05783_ (.A(_04955_),
    .Y(_04956_));
 sky130_fd_sc_hd__nand2_1 _05784_ (.A(_04807_),
    .B(_04956_),
    .Y(_04957_));
 sky130_fd_sc_hd__nand3_1 _05785_ (.A(_04803_),
    .B(_04806_),
    .C(_04955_),
    .Y(_04958_));
 sky130_fd_sc_hd__nand2_1 _05786_ (.A(_04957_),
    .B(_04958_),
    .Y(_04959_));
 sky130_fd_sc_hd__nand3_1 _05787_ (.A(_04938_),
    .B(_04939_),
    .C(_04941_),
    .Y(_04960_));
 sky130_fd_sc_hd__nand2_1 _05788_ (.A(_04943_),
    .B(_04960_),
    .Y(_04961_));
 sky130_fd_sc_hd__clkbuf_8 _05789_ (.A(net37),
    .X(_04962_));
 sky130_fd_sc_hd__nand2_1 _05790_ (.A(_04962_),
    .B(_04809_),
    .Y(_04963_));
 sky130_fd_sc_hd__clkbuf_8 _05791_ (.A(net36),
    .X(_04964_));
 sky130_fd_sc_hd__nand2_1 _05792_ (.A(_04964_),
    .B(_03820_),
    .Y(_04965_));
 sky130_fd_sc_hd__nand2_1 _05793_ (.A(_04963_),
    .B(_04965_),
    .Y(_04966_));
 sky130_fd_sc_hd__nand2_1 _05794_ (.A(_03809_),
    .B(_04819_),
    .Y(_04967_));
 sky130_fd_sc_hd__inv_2 _05795_ (.A(_04967_),
    .Y(_04968_));
 sky130_fd_sc_hd__nor2_1 _05796_ (.A(_04963_),
    .B(_04965_),
    .Y(_04969_));
 sky130_fd_sc_hd__a21oi_1 _05797_ (.A1(_04966_),
    .A2(_04968_),
    .B1(_04969_),
    .Y(_04970_));
 sky130_fd_sc_hd__nand2_1 _05798_ (.A(_04961_),
    .B(_04970_),
    .Y(_04971_));
 sky130_fd_sc_hd__nand2_1 _05799_ (.A(_04818_),
    .B(_04895_),
    .Y(_04972_));
 sky130_fd_sc_hd__nand2_1 _05800_ (.A(_04808_),
    .B(_04911_),
    .Y(_04973_));
 sky130_fd_sc_hd__inv_2 _05801_ (.A(_04973_),
    .Y(_04974_));
 sky130_fd_sc_hd__nand2_1 _05802_ (.A(_04812_),
    .B(_04827_),
    .Y(_04975_));
 sky130_fd_sc_hd__inv_2 _05803_ (.A(_04975_),
    .Y(_04976_));
 sky130_fd_sc_hd__nand2_1 _05804_ (.A(_04974_),
    .B(_04976_),
    .Y(_04977_));
 sky130_fd_sc_hd__nand2_1 _05805_ (.A(_04973_),
    .B(_04975_),
    .Y(_04978_));
 sky130_fd_sc_hd__nand3b_2 _05806_ (.A_N(_04972_),
    .B(_04977_),
    .C(_04978_),
    .Y(_04979_));
 sky130_fd_sc_hd__nand2_1 _05807_ (.A(_04979_),
    .B(_04977_),
    .Y(_04980_));
 sky130_fd_sc_hd__inv_2 _05808_ (.A(_04970_),
    .Y(_04981_));
 sky130_fd_sc_hd__nand3_1 _05809_ (.A(_04981_),
    .B(_04943_),
    .C(_04960_),
    .Y(_04982_));
 sky130_fd_sc_hd__a21boi_1 _05810_ (.A1(_04971_),
    .A2(_04980_),
    .B1_N(_04982_),
    .Y(_04983_));
 sky130_fd_sc_hd__nand2_1 _05811_ (.A(_04946_),
    .B(_04935_),
    .Y(_04984_));
 sky130_fd_sc_hd__inv_2 _05812_ (.A(_04944_),
    .Y(_04985_));
 sky130_fd_sc_hd__nand2_1 _05813_ (.A(_04984_),
    .B(_04985_),
    .Y(_04986_));
 sky130_fd_sc_hd__nand3_1 _05814_ (.A(_04946_),
    .B(_04935_),
    .C(_04944_),
    .Y(_04987_));
 sky130_fd_sc_hd__nand2_1 _05815_ (.A(_04986_),
    .B(_04987_),
    .Y(_04988_));
 sky130_fd_sc_hd__nor2_1 _05816_ (.A(_04983_),
    .B(_04988_),
    .Y(_04989_));
 sky130_fd_sc_hd__inv_2 _05817_ (.A(_04989_),
    .Y(_04990_));
 sky130_fd_sc_hd__buf_4 _05818_ (.A(_04911_),
    .X(_04991_));
 sky130_fd_sc_hd__clkbuf_8 _05819_ (.A(_04895_),
    .X(_04992_));
 sky130_fd_sc_hd__a22o_1 _05820_ (.A1(_04873_),
    .A2(_04991_),
    .B1(_04871_),
    .B2(_04992_),
    .X(_04993_));
 sky130_fd_sc_hd__and2_1 _05821_ (.A(_04913_),
    .B(_04993_),
    .X(_04994_));
 sky130_fd_sc_hd__nand2_1 _05822_ (.A(_04988_),
    .B(_04983_),
    .Y(_04995_));
 sky130_fd_sc_hd__nand3_1 _05823_ (.A(_04990_),
    .B(_04994_),
    .C(_04995_),
    .Y(_04996_));
 sky130_fd_sc_hd__nand2_1 _05824_ (.A(_04996_),
    .B(_04990_),
    .Y(_04997_));
 sky130_fd_sc_hd__nand2_1 _05825_ (.A(_03633_),
    .B(_03732_),
    .Y(_04998_));
 sky130_fd_sc_hd__nand3_1 _05826_ (.A(_03589_),
    .B(_03622_),
    .C(_03710_),
    .Y(_04999_));
 sky130_fd_sc_hd__nand3_1 _05827_ (.A(_04998_),
    .B(_03875_),
    .C(_04999_),
    .Y(_05000_));
 sky130_fd_sc_hd__nand2_1 _05828_ (.A(_03897_),
    .B(_05000_),
    .Y(_05001_));
 sky130_fd_sc_hd__nand2_1 _05829_ (.A(_02819_),
    .B(_02830_),
    .Y(_05002_));
 sky130_fd_sc_hd__nand2_1 _05830_ (.A(_05002_),
    .B(_02764_),
    .Y(_05003_));
 sky130_fd_sc_hd__nand2_1 _05831_ (.A(_05003_),
    .B(_02841_),
    .Y(_05004_));
 sky130_fd_sc_hd__nand2_1 _05832_ (.A(_01873_),
    .B(_01565_),
    .Y(_05005_));
 sky130_fd_sc_hd__inv_2 _05833_ (.A(_05005_),
    .Y(_05006_));
 sky130_fd_sc_hd__nand2_1 _05834_ (.A(net5),
    .B(_01048_),
    .Y(_05007_));
 sky130_fd_sc_hd__nand2_1 _05835_ (.A(net6),
    .B(_01092_),
    .Y(_05008_));
 sky130_fd_sc_hd__nand2_1 _05836_ (.A(_05007_),
    .B(_05008_),
    .Y(_05009_));
 sky130_fd_sc_hd__inv_2 _05837_ (.A(_05007_),
    .Y(_05010_));
 sky130_fd_sc_hd__inv_2 _05838_ (.A(_05008_),
    .Y(_05011_));
 sky130_fd_sc_hd__nand2_1 _05839_ (.A(_05010_),
    .B(_05011_),
    .Y(_05012_));
 sky130_fd_sc_hd__a21boi_1 _05840_ (.A1(_05006_),
    .A2(_05009_),
    .B1_N(_05012_),
    .Y(_05013_));
 sky130_fd_sc_hd__nand2_1 _05841_ (.A(_05004_),
    .B(_05013_),
    .Y(_05014_));
 sky130_fd_sc_hd__nand2_1 _05842_ (.A(_02753_),
    .B(_01774_),
    .Y(_05015_));
 sky130_fd_sc_hd__inv_2 _05843_ (.A(_05015_),
    .Y(_05016_));
 sky130_fd_sc_hd__nand2_1 _05844_ (.A(_02049_),
    .B(_01807_),
    .Y(_05017_));
 sky130_fd_sc_hd__inv_2 _05845_ (.A(_05017_),
    .Y(_05018_));
 sky130_fd_sc_hd__nand2_1 _05846_ (.A(_05016_),
    .B(_05018_),
    .Y(_05019_));
 sky130_fd_sc_hd__nand2_1 _05847_ (.A(_03182_),
    .B(_01884_),
    .Y(_05020_));
 sky130_fd_sc_hd__inv_2 _05848_ (.A(_05020_),
    .Y(_05021_));
 sky130_fd_sc_hd__nand2_1 _05849_ (.A(_05015_),
    .B(_05017_),
    .Y(_05022_));
 sky130_fd_sc_hd__nand3_1 _05850_ (.A(_05019_),
    .B(_05021_),
    .C(_05022_),
    .Y(_05023_));
 sky130_fd_sc_hd__nand2_1 _05851_ (.A(_05023_),
    .B(_05019_),
    .Y(_05024_));
 sky130_fd_sc_hd__nor2_1 _05852_ (.A(_05013_),
    .B(_05004_),
    .Y(_05025_));
 sky130_fd_sc_hd__a21oi_2 _05853_ (.A1(_05014_),
    .A2(_05024_),
    .B1(_05025_),
    .Y(_05026_));
 sky130_fd_sc_hd__nand2_1 _05854_ (.A(_05001_),
    .B(_05026_),
    .Y(_05027_));
 sky130_fd_sc_hd__buf_6 _05855_ (.A(_03314_),
    .X(_05028_));
 sky130_fd_sc_hd__buf_6 _05856_ (.A(_02995_),
    .X(_05029_));
 sky130_fd_sc_hd__nand2_2 _05857_ (.A(_05028_),
    .B(_05029_),
    .Y(_05030_));
 sky130_fd_sc_hd__clkbuf_8 _05858_ (.A(_03226_),
    .X(_05031_));
 sky130_fd_sc_hd__clkbuf_8 _05859_ (.A(_03028_),
    .X(_05032_));
 sky130_fd_sc_hd__nand2_2 _05860_ (.A(_05031_),
    .B(_05032_),
    .Y(_05033_));
 sky130_fd_sc_hd__nand2_1 _05861_ (.A(_05030_),
    .B(_05033_),
    .Y(_05034_));
 sky130_fd_sc_hd__nand2_1 _05862_ (.A(net35),
    .B(_04928_),
    .Y(_05035_));
 sky130_fd_sc_hd__inv_2 _05863_ (.A(_05035_),
    .Y(_05036_));
 sky130_fd_sc_hd__nor2_1 _05864_ (.A(_05030_),
    .B(_05033_),
    .Y(_05037_));
 sky130_fd_sc_hd__a21oi_2 _05865_ (.A1(_05034_),
    .A2(_05036_),
    .B1(_05037_),
    .Y(_05038_));
 sky130_fd_sc_hd__inv_2 _05866_ (.A(_03644_),
    .Y(_05039_));
 sky130_fd_sc_hd__inv_2 _05867_ (.A(_03655_),
    .Y(_05040_));
 sky130_fd_sc_hd__nand2_1 _05868_ (.A(_05039_),
    .B(_05040_),
    .Y(_05041_));
 sky130_fd_sc_hd__nand2_1 _05869_ (.A(_05041_),
    .B(_03666_),
    .Y(_05042_));
 sky130_fd_sc_hd__nand2_1 _05870_ (.A(_05042_),
    .B(_03677_),
    .Y(_05043_));
 sky130_fd_sc_hd__nand3_1 _05871_ (.A(_05041_),
    .B(_03688_),
    .C(_03666_),
    .Y(_05044_));
 sky130_fd_sc_hd__nand2_1 _05872_ (.A(_05043_),
    .B(_05044_),
    .Y(_05045_));
 sky130_fd_sc_hd__inv_2 _05873_ (.A(_05038_),
    .Y(_05046_));
 sky130_fd_sc_hd__nand2_1 _05874_ (.A(_05045_),
    .B(_05046_),
    .Y(_05047_));
 sky130_fd_sc_hd__nand3_1 _05875_ (.A(_05043_),
    .B(_05038_),
    .C(_05044_),
    .Y(_05048_));
 sky130_fd_sc_hd__nand2_1 _05876_ (.A(_05047_),
    .B(_05048_),
    .Y(_05049_));
 sky130_fd_sc_hd__inv_2 _05877_ (.A(_04930_),
    .Y(_05050_));
 sky130_fd_sc_hd__o21ai_1 _05878_ (.A1(_04933_),
    .A2(_05050_),
    .B1(_04931_),
    .Y(_05051_));
 sky130_fd_sc_hd__nand3b_1 _05879_ (.A_N(_04933_),
    .B(_04932_),
    .C(_04930_),
    .Y(_05052_));
 sky130_fd_sc_hd__nand2_1 _05880_ (.A(_05051_),
    .B(_05052_),
    .Y(_05053_));
 sky130_fd_sc_hd__inv_2 _05881_ (.A(_05053_),
    .Y(_05054_));
 sky130_fd_sc_hd__nand2_1 _05882_ (.A(_05049_),
    .B(_05054_),
    .Y(_05055_));
 sky130_fd_sc_hd__o21ai_2 _05883_ (.A1(_05038_),
    .A2(_05045_),
    .B1(_05055_),
    .Y(_05056_));
 sky130_fd_sc_hd__nor2_1 _05884_ (.A(_05026_),
    .B(_05001_),
    .Y(_05057_));
 sky130_fd_sc_hd__a21oi_2 _05885_ (.A1(_05027_),
    .A2(_05056_),
    .B1(_05057_),
    .Y(_05058_));
 sky130_fd_sc_hd__nand3_1 _05886_ (.A(_04948_),
    .B(_04922_),
    .C(_04921_),
    .Y(_05059_));
 sky130_fd_sc_hd__inv_2 _05887_ (.A(_04948_),
    .Y(_05060_));
 sky130_fd_sc_hd__nand2_1 _05888_ (.A(_05060_),
    .B(_04923_),
    .Y(_05061_));
 sky130_fd_sc_hd__nand2_1 _05889_ (.A(_05059_),
    .B(_05061_),
    .Y(_05062_));
 sky130_fd_sc_hd__nand2_1 _05890_ (.A(_05062_),
    .B(_04919_),
    .Y(_05063_));
 sky130_fd_sc_hd__nand3_1 _05891_ (.A(_05059_),
    .B(_05061_),
    .C(_04918_),
    .Y(_05064_));
 sky130_fd_sc_hd__nand3_1 _05892_ (.A(_05058_),
    .B(_05063_),
    .C(_05064_),
    .Y(_05065_));
 sky130_fd_sc_hd__nand2_1 _05893_ (.A(_05063_),
    .B(_05064_),
    .Y(_05066_));
 sky130_fd_sc_hd__inv_2 _05894_ (.A(_05058_),
    .Y(_05067_));
 sky130_fd_sc_hd__nand2_1 _05895_ (.A(_05066_),
    .B(_05067_),
    .Y(_05068_));
 sky130_fd_sc_hd__nand3b_1 _05896_ (.A_N(_04997_),
    .B(_05065_),
    .C(_05068_),
    .Y(_05069_));
 sky130_fd_sc_hd__nand2_1 _05897_ (.A(_05068_),
    .B(_05065_),
    .Y(_05070_));
 sky130_fd_sc_hd__nand2_1 _05898_ (.A(_05070_),
    .B(_04997_),
    .Y(_05071_));
 sky130_fd_sc_hd__nand2_1 _05899_ (.A(_05069_),
    .B(_05071_),
    .Y(_05072_));
 sky130_fd_sc_hd__inv_2 _05900_ (.A(_05072_),
    .Y(_05073_));
 sky130_fd_sc_hd__inv_2 _05901_ (.A(_02951_),
    .Y(_05074_));
 sky130_fd_sc_hd__nand2_1 _05902_ (.A(_02214_),
    .B(_05074_),
    .Y(_05075_));
 sky130_fd_sc_hd__nand3_1 _05903_ (.A(_02951_),
    .B(_02192_),
    .C(_02203_),
    .Y(_05076_));
 sky130_fd_sc_hd__nand2_1 _05904_ (.A(_05075_),
    .B(_05076_),
    .Y(_05077_));
 sky130_fd_sc_hd__nand2_1 _05905_ (.A(_05077_),
    .B(_03963_),
    .Y(_05078_));
 sky130_fd_sc_hd__nand3_1 _05906_ (.A(_05075_),
    .B(_05076_),
    .C(_03952_),
    .Y(_05079_));
 sky130_fd_sc_hd__nand2_1 _05907_ (.A(_05078_),
    .B(_05079_),
    .Y(_05080_));
 sky130_fd_sc_hd__nand3_1 _05908_ (.A(_02632_),
    .B(_01719_),
    .C(_02247_),
    .Y(_05081_));
 sky130_fd_sc_hd__inv_2 _05909_ (.A(_02445_),
    .Y(_05082_));
 sky130_fd_sc_hd__nand3_1 _05910_ (.A(_05082_),
    .B(_02335_),
    .C(_02313_),
    .Y(_05083_));
 sky130_fd_sc_hd__nand3_1 _05911_ (.A(_05083_),
    .B(_02456_),
    .C(_02610_),
    .Y(_05084_));
 sky130_fd_sc_hd__nand2_1 _05912_ (.A(_05084_),
    .B(_05083_),
    .Y(_05085_));
 sky130_fd_sc_hd__nand2_1 _05913_ (.A(_02258_),
    .B(_05085_),
    .Y(_05086_));
 sky130_fd_sc_hd__nand2_1 _05914_ (.A(_05081_),
    .B(_05086_),
    .Y(_05087_));
 sky130_fd_sc_hd__nand2_1 _05915_ (.A(_05087_),
    .B(_02929_),
    .Y(_05088_));
 sky130_fd_sc_hd__nand3_1 _05916_ (.A(_05081_),
    .B(_05086_),
    .C(_02918_),
    .Y(_05089_));
 sky130_fd_sc_hd__nand2_1 _05917_ (.A(_05088_),
    .B(_05089_),
    .Y(_05090_));
 sky130_fd_sc_hd__nand3_1 _05918_ (.A(_05012_),
    .B(_05006_),
    .C(_05009_),
    .Y(_05091_));
 sky130_fd_sc_hd__nand2_1 _05919_ (.A(_05091_),
    .B(_05012_),
    .Y(_05092_));
 sky130_fd_sc_hd__nand3_1 _05920_ (.A(_05092_),
    .B(_02841_),
    .C(_05003_),
    .Y(_05093_));
 sky130_fd_sc_hd__nand2_1 _05921_ (.A(_05093_),
    .B(_05014_),
    .Y(_05094_));
 sky130_fd_sc_hd__inv_2 _05922_ (.A(_05024_),
    .Y(_05095_));
 sky130_fd_sc_hd__nand2_1 _05923_ (.A(_05094_),
    .B(_05095_),
    .Y(_05096_));
 sky130_fd_sc_hd__nand3_1 _05924_ (.A(_05093_),
    .B(_05014_),
    .C(_05024_),
    .Y(_05097_));
 sky130_fd_sc_hd__nand2_1 _05925_ (.A(_05096_),
    .B(_05097_),
    .Y(_05098_));
 sky130_fd_sc_hd__inv_2 _05926_ (.A(_05098_),
    .Y(_05099_));
 sky130_fd_sc_hd__nand2_1 _05927_ (.A(_02346_),
    .B(_05082_),
    .Y(_05100_));
 sky130_fd_sc_hd__nand3_1 _05928_ (.A(_02445_),
    .B(_02313_),
    .C(_02335_),
    .Y(_05101_));
 sky130_fd_sc_hd__nand3_1 _05929_ (.A(_05100_),
    .B(_05101_),
    .C(_02599_),
    .Y(_05102_));
 sky130_fd_sc_hd__nand2_1 _05930_ (.A(_05084_),
    .B(_05102_),
    .Y(_05103_));
 sky130_fd_sc_hd__inv_2 _05931_ (.A(_02368_),
    .Y(_05104_));
 sky130_fd_sc_hd__nand2_1 _05932_ (.A(_05104_),
    .B(_02390_),
    .Y(_05105_));
 sky130_fd_sc_hd__inv_2 _05933_ (.A(_02390_),
    .Y(_05106_));
 sky130_fd_sc_hd__nand2_1 _05934_ (.A(_05106_),
    .B(_02368_),
    .Y(_05107_));
 sky130_fd_sc_hd__nand3_1 _05935_ (.A(_05105_),
    .B(_05107_),
    .C(_02412_),
    .Y(_05108_));
 sky130_fd_sc_hd__nand2_1 _05936_ (.A(_05104_),
    .B(_05106_),
    .Y(_05109_));
 sky130_fd_sc_hd__nand3_1 _05937_ (.A(_05109_),
    .B(_02423_),
    .C(_02401_),
    .Y(_05110_));
 sky130_fd_sc_hd__nand2_1 _05938_ (.A(_05108_),
    .B(_05110_),
    .Y(_05111_));
 sky130_fd_sc_hd__nand2_1 _05939_ (.A(_01037_),
    .B(_02357_),
    .Y(_05112_));
 sky130_fd_sc_hd__nand2_1 _05940_ (.A(_01081_),
    .B(_02379_),
    .Y(_05113_));
 sky130_fd_sc_hd__nand2_1 _05941_ (.A(_05112_),
    .B(_05113_),
    .Y(_05114_));
 sky130_fd_sc_hd__nand2_1 _05942_ (.A(_01147_),
    .B(_00861_),
    .Y(_05115_));
 sky130_fd_sc_hd__inv_2 _05943_ (.A(_05115_),
    .Y(_05116_));
 sky130_fd_sc_hd__nor2_1 _05944_ (.A(_05112_),
    .B(_05113_),
    .Y(_05117_));
 sky130_fd_sc_hd__a21oi_2 _05945_ (.A1(_05114_),
    .A2(_05116_),
    .B1(_05117_),
    .Y(_05118_));
 sky130_fd_sc_hd__nand2_1 _05946_ (.A(_05111_),
    .B(_05118_),
    .Y(_05119_));
 sky130_fd_sc_hd__nand2_1 _05947_ (.A(_05010_),
    .B(_05008_),
    .Y(_05120_));
 sky130_fd_sc_hd__nand2_1 _05948_ (.A(_05011_),
    .B(_05007_),
    .Y(_05121_));
 sky130_fd_sc_hd__nand3_1 _05949_ (.A(_05120_),
    .B(_05121_),
    .C(_05005_),
    .Y(_05122_));
 sky130_fd_sc_hd__nand2_1 _05950_ (.A(_05122_),
    .B(_05091_),
    .Y(_05123_));
 sky130_fd_sc_hd__inv_2 _05951_ (.A(_05123_),
    .Y(_05124_));
 sky130_fd_sc_hd__nor2_1 _05952_ (.A(_05118_),
    .B(_05111_),
    .Y(_05125_));
 sky130_fd_sc_hd__a21oi_1 _05953_ (.A1(_05119_),
    .A2(_05124_),
    .B1(_05125_),
    .Y(_05126_));
 sky130_fd_sc_hd__nand2_1 _05954_ (.A(_05103_),
    .B(_05126_),
    .Y(_05127_));
 sky130_fd_sc_hd__nor2_1 _05955_ (.A(_05126_),
    .B(_05103_),
    .Y(_05128_));
 sky130_fd_sc_hd__a21oi_1 _05956_ (.A1(_05099_),
    .A2(_05127_),
    .B1(_05128_),
    .Y(_05129_));
 sky130_fd_sc_hd__nand2_1 _05957_ (.A(_05090_),
    .B(_05129_),
    .Y(_05130_));
 sky130_fd_sc_hd__inv_2 _05958_ (.A(_05026_),
    .Y(_05131_));
 sky130_fd_sc_hd__nand2_1 _05959_ (.A(_05001_),
    .B(_05131_),
    .Y(_05132_));
 sky130_fd_sc_hd__nand3_1 _05960_ (.A(_05026_),
    .B(_03897_),
    .C(_05000_),
    .Y(_05133_));
 sky130_fd_sc_hd__nand2_1 _05961_ (.A(_05132_),
    .B(_05133_),
    .Y(_05134_));
 sky130_fd_sc_hd__nand2_1 _05962_ (.A(_05134_),
    .B(_05056_),
    .Y(_05135_));
 sky130_fd_sc_hd__nand3b_1 _05963_ (.A_N(_05056_),
    .B(_05132_),
    .C(_05133_),
    .Y(_05136_));
 sky130_fd_sc_hd__nand2_1 _05964_ (.A(_05135_),
    .B(_05136_),
    .Y(_05137_));
 sky130_fd_sc_hd__inv_2 _05965_ (.A(_05137_),
    .Y(_05138_));
 sky130_fd_sc_hd__nor2_1 _05966_ (.A(_05129_),
    .B(_05090_),
    .Y(_05139_));
 sky130_fd_sc_hd__a21oi_1 _05967_ (.A1(_05130_),
    .A2(_05138_),
    .B1(_05139_),
    .Y(_05140_));
 sky130_fd_sc_hd__nand2_1 _05968_ (.A(_05080_),
    .B(_05140_),
    .Y(_05141_));
 sky130_fd_sc_hd__nor2_1 _05969_ (.A(_05140_),
    .B(_05080_),
    .Y(_05142_));
 sky130_fd_sc_hd__a21oi_1 _05970_ (.A1(_05073_),
    .A2(_05141_),
    .B1(_05142_),
    .Y(_05143_));
 sky130_fd_sc_hd__nand2_1 _05971_ (.A(_04959_),
    .B(_05143_),
    .Y(_05144_));
 sky130_fd_sc_hd__o21a_1 _05972_ (.A1(_05066_),
    .A2(_05058_),
    .B1(_05071_),
    .X(_05145_));
 sky130_fd_sc_hd__xor2_2 _05973_ (.A(_04916_),
    .B(_05145_),
    .X(_05146_));
 sky130_fd_sc_hd__nor2_1 _05974_ (.A(_05143_),
    .B(_04959_),
    .Y(_05147_));
 sky130_fd_sc_hd__a21oi_1 _05975_ (.A1(_05144_),
    .A2(_05146_),
    .B1(_05147_),
    .Y(_05148_));
 sky130_fd_sc_hd__nand2_1 _05976_ (.A(_04804_),
    .B(_03985_),
    .Y(_05149_));
 sky130_fd_sc_hd__nor2_1 _05977_ (.A(_03985_),
    .B(_04804_),
    .Y(_05150_));
 sky130_fd_sc_hd__a21o_1 _05978_ (.A1(_05149_),
    .A2(_04956_),
    .B1(_05150_),
    .X(_05151_));
 sky130_fd_sc_hd__nor2_1 _05979_ (.A(_04797_),
    .B(_04796_),
    .Y(_05152_));
 sky130_fd_sc_hd__a21oi_2 _05980_ (.A1(_04798_),
    .A2(_04795_),
    .B1(_05152_),
    .Y(_05153_));
 sky130_fd_sc_hd__nor2_1 _05981_ (.A(_04730_),
    .B(_04712_),
    .Y(_05154_));
 sky130_fd_sc_hd__a21o_1 _05982_ (.A1(_04738_),
    .A2(_04704_),
    .B1(_05154_),
    .X(_05155_));
 sky130_fd_sc_hd__nor2_1 _05983_ (.A(_04062_),
    .B(_04238_),
    .Y(_05156_));
 sky130_fd_sc_hd__a21oi_1 _05984_ (.A1(_04249_),
    .A2(_04414_),
    .B1(_05156_),
    .Y(_05157_));
 sky130_fd_sc_hd__nand2_1 _05985_ (.A(_00751_),
    .B(_04084_),
    .Y(_05158_));
 sky130_fd_sc_hd__inv_2 _05986_ (.A(_05158_),
    .Y(_05159_));
 sky130_fd_sc_hd__buf_4 _05987_ (.A(net15),
    .X(_05160_));
 sky130_fd_sc_hd__nand2_1 _05988_ (.A(_00795_),
    .B(_05160_),
    .Y(_05161_));
 sky130_fd_sc_hd__inv_2 _05989_ (.A(_05161_),
    .Y(_05162_));
 sky130_fd_sc_hd__nand2_1 _05990_ (.A(_05159_),
    .B(_05162_),
    .Y(_05163_));
 sky130_fd_sc_hd__nand2_1 _05991_ (.A(_05158_),
    .B(_05161_),
    .Y(_05164_));
 sky130_fd_sc_hd__nand2_1 _05992_ (.A(_05163_),
    .B(_05164_),
    .Y(_05165_));
 sky130_fd_sc_hd__nand2_1 _05993_ (.A(_01323_),
    .B(_00861_),
    .Y(_05166_));
 sky130_fd_sc_hd__nand2_1 _05994_ (.A(_05165_),
    .B(_05166_),
    .Y(_05167_));
 sky130_fd_sc_hd__inv_2 _05995_ (.A(_05166_),
    .Y(_05168_));
 sky130_fd_sc_hd__nand3_2 _05996_ (.A(_05163_),
    .B(_05168_),
    .C(_05164_),
    .Y(_05169_));
 sky130_fd_sc_hd__nand2_1 _05997_ (.A(_05167_),
    .B(_05169_),
    .Y(_05170_));
 sky130_fd_sc_hd__nor2_1 _05998_ (.A(_04095_),
    .B(_04117_),
    .Y(_05171_));
 sky130_fd_sc_hd__a21oi_1 _05999_ (.A1(_04172_),
    .A2(_04161_),
    .B1(_05171_),
    .Y(_05172_));
 sky130_fd_sc_hd__nand2_1 _06000_ (.A(_05170_),
    .B(_05172_),
    .Y(_05173_));
 sky130_fd_sc_hd__a21o_1 _06001_ (.A1(_04172_),
    .A2(_04161_),
    .B1(_05171_),
    .X(_05174_));
 sky130_fd_sc_hd__nand3_2 _06002_ (.A(_05174_),
    .B(_05169_),
    .C(_05167_),
    .Y(_05175_));
 sky130_fd_sc_hd__nand2_1 _06003_ (.A(_00740_),
    .B(_01048_),
    .Y(_05176_));
 sky130_fd_sc_hd__inv_2 _06004_ (.A(_05176_),
    .Y(_05177_));
 sky130_fd_sc_hd__nand2_1 _06005_ (.A(_00784_),
    .B(_01092_),
    .Y(_05178_));
 sky130_fd_sc_hd__inv_2 _06006_ (.A(_05178_),
    .Y(_05179_));
 sky130_fd_sc_hd__nand2_1 _06007_ (.A(_05177_),
    .B(_05179_),
    .Y(_05180_));
 sky130_fd_sc_hd__nand2_1 _06008_ (.A(_05176_),
    .B(_05178_),
    .Y(_05181_));
 sky130_fd_sc_hd__nand2_1 _06009_ (.A(_05180_),
    .B(_05181_),
    .Y(_05182_));
 sky130_fd_sc_hd__nand2_1 _06010_ (.A(_00850_),
    .B(_01158_),
    .Y(_05183_));
 sky130_fd_sc_hd__nand2_1 _06011_ (.A(_05182_),
    .B(_05183_),
    .Y(_05184_));
 sky130_fd_sc_hd__inv_2 _06012_ (.A(_05183_),
    .Y(_05185_));
 sky130_fd_sc_hd__nand3_1 _06013_ (.A(_05180_),
    .B(_05185_),
    .C(_05181_),
    .Y(_05186_));
 sky130_fd_sc_hd__nand2_1 _06014_ (.A(_05184_),
    .B(_05186_),
    .Y(_05187_));
 sky130_fd_sc_hd__inv_2 _06015_ (.A(_05187_),
    .Y(_05188_));
 sky130_fd_sc_hd__nand3_1 _06016_ (.A(_05173_),
    .B(_05175_),
    .C(_05188_),
    .Y(_05189_));
 sky130_fd_sc_hd__nand2_1 _06017_ (.A(_05170_),
    .B(_05174_),
    .Y(_05190_));
 sky130_fd_sc_hd__nand3_1 _06018_ (.A(_05167_),
    .B(_05172_),
    .C(_05169_),
    .Y(_05191_));
 sky130_fd_sc_hd__nand3_1 _06019_ (.A(_05190_),
    .B(_05191_),
    .C(_05187_),
    .Y(_05192_));
 sky130_fd_sc_hd__nand3_1 _06020_ (.A(_05157_),
    .B(_05189_),
    .C(_05192_),
    .Y(_05193_));
 sky130_fd_sc_hd__nand2_1 _06021_ (.A(_05189_),
    .B(_05192_),
    .Y(_05194_));
 sky130_fd_sc_hd__nand2_1 _06022_ (.A(_04425_),
    .B(_04227_),
    .Y(_05195_));
 sky130_fd_sc_hd__nand2_1 _06023_ (.A(_05194_),
    .B(_05195_),
    .Y(_05196_));
 sky130_fd_sc_hd__nand2_1 _06024_ (.A(_05193_),
    .B(_05196_),
    .Y(_05197_));
 sky130_fd_sc_hd__nand2_1 _06025_ (.A(_01037_),
    .B(_01774_),
    .Y(_05198_));
 sky130_fd_sc_hd__inv_2 _06026_ (.A(_05198_),
    .Y(_05199_));
 sky130_fd_sc_hd__nand2_1 _06027_ (.A(net8),
    .B(_01807_),
    .Y(_05200_));
 sky130_fd_sc_hd__inv_2 _06028_ (.A(_05200_),
    .Y(_05201_));
 sky130_fd_sc_hd__nand2_1 _06029_ (.A(_05199_),
    .B(_05201_),
    .Y(_00000_));
 sky130_fd_sc_hd__nand2_1 _06030_ (.A(_05198_),
    .B(_05200_),
    .Y(_00001_));
 sky130_fd_sc_hd__nand2_1 _06031_ (.A(_00000_),
    .B(_00001_),
    .Y(_00002_));
 sky130_fd_sc_hd__buf_6 _06032_ (.A(_01884_),
    .X(_00003_));
 sky130_fd_sc_hd__nand2_1 _06033_ (.A(_01147_),
    .B(_00003_),
    .Y(_00004_));
 sky130_fd_sc_hd__nand2_1 _06034_ (.A(_00002_),
    .B(_00004_),
    .Y(_00005_));
 sky130_fd_sc_hd__nand3b_2 _06035_ (.A_N(_00004_),
    .B(_00000_),
    .C(_00001_),
    .Y(_00006_));
 sky130_fd_sc_hd__nand2_1 _06036_ (.A(_00005_),
    .B(_00006_),
    .Y(_00007_));
 sky130_fd_sc_hd__nor2_1 _06037_ (.A(_04271_),
    .B(_04304_),
    .Y(_00008_));
 sky130_fd_sc_hd__a21oi_2 _06038_ (.A1(_04337_),
    .A2(_04381_),
    .B1(_00008_),
    .Y(_00009_));
 sky130_fd_sc_hd__inv_2 _06039_ (.A(_00009_),
    .Y(_00010_));
 sky130_fd_sc_hd__nand2_1 _06040_ (.A(_00007_),
    .B(_00010_),
    .Y(_00011_));
 sky130_fd_sc_hd__nand3_1 _06041_ (.A(_00005_),
    .B(_00006_),
    .C(_00009_),
    .Y(_00012_));
 sky130_fd_sc_hd__nand2_1 _06042_ (.A(_00011_),
    .B(_00012_),
    .Y(_00013_));
 sky130_fd_sc_hd__nand2_1 _06043_ (.A(_04578_),
    .B(_04520_),
    .Y(_00014_));
 sky130_fd_sc_hd__nand2_1 _06044_ (.A(_00013_),
    .B(_00014_),
    .Y(_00015_));
 sky130_fd_sc_hd__nand3b_1 _06045_ (.A_N(_00014_),
    .B(_00011_),
    .C(_00012_),
    .Y(_00016_));
 sky130_fd_sc_hd__nand2_1 _06046_ (.A(_00015_),
    .B(_00016_),
    .Y(_00017_));
 sky130_fd_sc_hd__inv_2 _06047_ (.A(_00017_),
    .Y(_00018_));
 sky130_fd_sc_hd__nand2_1 _06048_ (.A(_05197_),
    .B(_00018_),
    .Y(_00019_));
 sky130_fd_sc_hd__nand3_1 _06049_ (.A(_05193_),
    .B(_05196_),
    .C(_00017_),
    .Y(_00020_));
 sky130_fd_sc_hd__nand3_1 _06050_ (.A(_05155_),
    .B(_00019_),
    .C(_00020_),
    .Y(_00021_));
 sky130_fd_sc_hd__nand2_1 _06051_ (.A(_00019_),
    .B(_00020_),
    .Y(_00022_));
 sky130_fd_sc_hd__a21oi_1 _06052_ (.A1(_04738_),
    .A2(_04704_),
    .B1(_05154_),
    .Y(_00023_));
 sky130_fd_sc_hd__nand2_1 _06053_ (.A(_00022_),
    .B(_00023_),
    .Y(_00024_));
 sky130_fd_sc_hd__nand2_1 _06054_ (.A(net37),
    .B(_03094_),
    .Y(_00025_));
 sky130_fd_sc_hd__nand2_1 _06055_ (.A(_04964_),
    .B(_03160_),
    .Y(_00026_));
 sky130_fd_sc_hd__nor2_1 _06056_ (.A(_00025_),
    .B(_00026_),
    .Y(_00027_));
 sky130_fd_sc_hd__inv_2 _06057_ (.A(_00027_),
    .Y(_00028_));
 sky130_fd_sc_hd__nand2_1 _06058_ (.A(_00025_),
    .B(_00026_),
    .Y(_00029_));
 sky130_fd_sc_hd__nand2_1 _06059_ (.A(_00028_),
    .B(_00029_),
    .Y(_00030_));
 sky130_fd_sc_hd__nand2_1 _06060_ (.A(_03809_),
    .B(_03226_),
    .Y(_00031_));
 sky130_fd_sc_hd__nand2_1 _06061_ (.A(_00030_),
    .B(_00031_),
    .Y(_00032_));
 sky130_fd_sc_hd__inv_2 _06062_ (.A(_00031_),
    .Y(_00033_));
 sky130_fd_sc_hd__nand3_1 _06063_ (.A(_00028_),
    .B(_00033_),
    .C(_00029_),
    .Y(_00034_));
 sky130_fd_sc_hd__nand2_1 _06064_ (.A(_00032_),
    .B(_00034_),
    .Y(_00035_));
 sky130_fd_sc_hd__nor2_1 _06065_ (.A(_04751_),
    .B(_04753_),
    .Y(_00036_));
 sky130_fd_sc_hd__a21oi_2 _06066_ (.A1(_04756_),
    .A2(_04760_),
    .B1(_00036_),
    .Y(_00037_));
 sky130_fd_sc_hd__inv_2 _06067_ (.A(_00037_),
    .Y(_00038_));
 sky130_fd_sc_hd__nand2_1 _06068_ (.A(_01873_),
    .B(_02995_),
    .Y(_00039_));
 sky130_fd_sc_hd__inv_2 _06069_ (.A(_00039_),
    .Y(_00040_));
 sky130_fd_sc_hd__nand2_1 _06070_ (.A(_02544_),
    .B(_03028_),
    .Y(_00041_));
 sky130_fd_sc_hd__inv_2 _06071_ (.A(_00041_),
    .Y(_00042_));
 sky130_fd_sc_hd__nand2_1 _06072_ (.A(_00040_),
    .B(_00042_),
    .Y(_00043_));
 sky130_fd_sc_hd__nand2_1 _06073_ (.A(_03215_),
    .B(_02049_),
    .Y(_00044_));
 sky130_fd_sc_hd__inv_2 _06074_ (.A(_00044_),
    .Y(_00045_));
 sky130_fd_sc_hd__nand2_1 _06075_ (.A(_00039_),
    .B(_00041_),
    .Y(_00046_));
 sky130_fd_sc_hd__nand3_1 _06076_ (.A(_00043_),
    .B(_00045_),
    .C(_00046_),
    .Y(_00047_));
 sky130_fd_sc_hd__nand2_1 _06077_ (.A(_00043_),
    .B(_00046_),
    .Y(_00048_));
 sky130_fd_sc_hd__nand2_1 _06078_ (.A(_00048_),
    .B(_00044_),
    .Y(_00049_));
 sky130_fd_sc_hd__nand3_1 _06079_ (.A(_00038_),
    .B(_00047_),
    .C(_00049_),
    .Y(_00050_));
 sky130_fd_sc_hd__nand2_1 _06080_ (.A(_00049_),
    .B(_00047_),
    .Y(_00051_));
 sky130_fd_sc_hd__nand2_1 _06081_ (.A(_00051_),
    .B(_00037_),
    .Y(_00052_));
 sky130_fd_sc_hd__nand3b_1 _06082_ (.A_N(_00035_),
    .B(_00050_),
    .C(_00052_),
    .Y(_00053_));
 sky130_fd_sc_hd__nand2_1 _06083_ (.A(_00051_),
    .B(_00038_),
    .Y(_00054_));
 sky130_fd_sc_hd__nand3_1 _06084_ (.A(_00049_),
    .B(_00037_),
    .C(_00047_),
    .Y(_00055_));
 sky130_fd_sc_hd__nand3_1 _06085_ (.A(_00054_),
    .B(_00055_),
    .C(_00035_),
    .Y(_00056_));
 sky130_fd_sc_hd__nand2_1 _06086_ (.A(_00053_),
    .B(_00056_),
    .Y(_00057_));
 sky130_fd_sc_hd__nor2_1 _06087_ (.A(_04607_),
    .B(_04588_),
    .Y(_00058_));
 sky130_fd_sc_hd__a21oi_2 _06088_ (.A1(_04617_),
    .A2(_04646_),
    .B1(_00058_),
    .Y(_00059_));
 sky130_fd_sc_hd__inv_2 _06089_ (.A(_00059_),
    .Y(_00060_));
 sky130_fd_sc_hd__nand2_1 _06090_ (.A(_00057_),
    .B(_00060_),
    .Y(_00061_));
 sky130_fd_sc_hd__nand3_1 _06091_ (.A(_00059_),
    .B(_00053_),
    .C(_00056_),
    .Y(_00062_));
 sky130_fd_sc_hd__nand2_1 _06092_ (.A(_00061_),
    .B(_00062_),
    .Y(_00063_));
 sky130_fd_sc_hd__nand2_1 _06093_ (.A(_04781_),
    .B(_04767_),
    .Y(_00064_));
 sky130_fd_sc_hd__nand2_1 _06094_ (.A(_00063_),
    .B(_00064_),
    .Y(_00065_));
 sky130_fd_sc_hd__nand3b_1 _06095_ (.A_N(_00064_),
    .B(_00061_),
    .C(_00062_),
    .Y(_00066_));
 sky130_fd_sc_hd__nand2_1 _06096_ (.A(_00065_),
    .B(_00066_),
    .Y(_00067_));
 sky130_fd_sc_hd__inv_2 _06097_ (.A(_00067_),
    .Y(_00068_));
 sky130_fd_sc_hd__nand3_1 _06098_ (.A(_00021_),
    .B(_00024_),
    .C(_00068_),
    .Y(_00069_));
 sky130_fd_sc_hd__nand2_1 _06099_ (.A(_00022_),
    .B(_05155_),
    .Y(_00070_));
 sky130_fd_sc_hd__nand3_1 _06100_ (.A(_00023_),
    .B(_00019_),
    .C(_00020_),
    .Y(_00071_));
 sky130_fd_sc_hd__nand3_1 _06101_ (.A(_00070_),
    .B(_00071_),
    .C(_00067_),
    .Y(_00072_));
 sky130_fd_sc_hd__nand3_1 _06102_ (.A(_05153_),
    .B(_00069_),
    .C(_00072_),
    .Y(_00073_));
 sky130_fd_sc_hd__nand2_1 _06103_ (.A(_00069_),
    .B(_00072_),
    .Y(_00074_));
 sky130_fd_sc_hd__a21o_1 _06104_ (.A1(_04798_),
    .A2(_04795_),
    .B1(_05152_),
    .X(_00075_));
 sky130_fd_sc_hd__nand2_1 _06105_ (.A(_00074_),
    .B(_00075_),
    .Y(_00076_));
 sky130_fd_sc_hd__nand2_1 _06106_ (.A(_00073_),
    .B(_00076_),
    .Y(_00077_));
 sky130_fd_sc_hd__nor2_1 _06107_ (.A(_04852_),
    .B(_04850_),
    .Y(_00078_));
 sky130_fd_sc_hd__a21oi_1 _06108_ (.A1(_04853_),
    .A2(_04856_),
    .B1(_00078_),
    .Y(_00079_));
 sky130_fd_sc_hd__nand2_1 _06109_ (.A(_04808_),
    .B(_03402_),
    .Y(_00080_));
 sky130_fd_sc_hd__inv_2 _06110_ (.A(_00080_),
    .Y(_00081_));
 sky130_fd_sc_hd__nand2_1 _06111_ (.A(_04812_),
    .B(_03314_),
    .Y(_00082_));
 sky130_fd_sc_hd__inv_2 _06112_ (.A(_00082_),
    .Y(_00083_));
 sky130_fd_sc_hd__nand2_1 _06113_ (.A(_00081_),
    .B(_00083_),
    .Y(_00084_));
 sky130_fd_sc_hd__nand2_1 _06114_ (.A(_00080_),
    .B(_00082_),
    .Y(_00085_));
 sky130_fd_sc_hd__nand2_1 _06115_ (.A(_00084_),
    .B(_00085_),
    .Y(_00086_));
 sky130_fd_sc_hd__nand2_1 _06116_ (.A(_04818_),
    .B(_03820_),
    .Y(_00087_));
 sky130_fd_sc_hd__nand2_1 _06117_ (.A(_00086_),
    .B(_00087_),
    .Y(_00088_));
 sky130_fd_sc_hd__inv_2 _06118_ (.A(_00087_),
    .Y(_00089_));
 sky130_fd_sc_hd__nand3_1 _06119_ (.A(_00084_),
    .B(_00089_),
    .C(_00085_),
    .Y(_00090_));
 sky130_fd_sc_hd__nand2_1 _06120_ (.A(_00088_),
    .B(_00090_),
    .Y(_00091_));
 sky130_fd_sc_hd__nor2_1 _06121_ (.A(_04768_),
    .B(_04770_),
    .Y(_00092_));
 sky130_fd_sc_hd__a21oi_1 _06122_ (.A1(_04773_),
    .A2(_04777_),
    .B1(_00092_),
    .Y(_00093_));
 sky130_fd_sc_hd__nand2_1 _06123_ (.A(_00091_),
    .B(_00093_),
    .Y(_00094_));
 sky130_fd_sc_hd__a21o_1 _06124_ (.A1(_04773_),
    .A2(_04777_),
    .B1(_00092_),
    .X(_00095_));
 sky130_fd_sc_hd__nand3_1 _06125_ (.A(_00095_),
    .B(_00090_),
    .C(_00088_),
    .Y(_00096_));
 sky130_fd_sc_hd__nand2_1 _06126_ (.A(_04849_),
    .B(_04844_),
    .Y(_00097_));
 sky130_fd_sc_hd__nand3_1 _06127_ (.A(_00094_),
    .B(_00096_),
    .C(_00097_),
    .Y(_00098_));
 sky130_fd_sc_hd__nand2_1 _06128_ (.A(_00091_),
    .B(_00095_),
    .Y(_00099_));
 sky130_fd_sc_hd__nand3_1 _06129_ (.A(_00088_),
    .B(_00093_),
    .C(_00090_),
    .Y(_00100_));
 sky130_fd_sc_hd__inv_2 _06130_ (.A(_00097_),
    .Y(_00101_));
 sky130_fd_sc_hd__nand3_1 _06131_ (.A(_00099_),
    .B(_00100_),
    .C(_00101_),
    .Y(_00102_));
 sky130_fd_sc_hd__nand3_1 _06132_ (.A(_00079_),
    .B(_00098_),
    .C(_00102_),
    .Y(_00103_));
 sky130_fd_sc_hd__nand2_1 _06133_ (.A(_04857_),
    .B(_04855_),
    .Y(_00104_));
 sky130_fd_sc_hd__nand2_1 _06134_ (.A(_00098_),
    .B(_00102_),
    .Y(_00105_));
 sky130_fd_sc_hd__nand2_1 _06135_ (.A(_00104_),
    .B(_00105_),
    .Y(_00106_));
 sky130_fd_sc_hd__nand2_1 _06136_ (.A(_00103_),
    .B(_00106_),
    .Y(_00107_));
 sky130_fd_sc_hd__nand2_1 _06137_ (.A(_04871_),
    .B(_04819_),
    .Y(_00108_));
 sky130_fd_sc_hd__nand3b_1 _06138_ (.A_N(_00108_),
    .B(_04873_),
    .C(_04809_),
    .Y(_00109_));
 sky130_fd_sc_hd__inv_2 _06139_ (.A(_04873_),
    .Y(_00110_));
 sky130_fd_sc_hd__inv_2 _06140_ (.A(_04809_),
    .Y(_00111_));
 sky130_fd_sc_hd__o21ai_2 _06141_ (.A1(_00110_),
    .A2(_00111_),
    .B1(_00108_),
    .Y(_00112_));
 sky130_fd_sc_hd__nand2_1 _06142_ (.A(_00109_),
    .B(_00112_),
    .Y(_00113_));
 sky130_fd_sc_hd__nand2_1 _06143_ (.A(_04876_),
    .B(_04827_),
    .Y(_00114_));
 sky130_fd_sc_hd__nand2_1 _06144_ (.A(_00113_),
    .B(_00114_),
    .Y(_00115_));
 sky130_fd_sc_hd__inv_2 _06145_ (.A(_00114_),
    .Y(_00116_));
 sky130_fd_sc_hd__nand3_1 _06146_ (.A(_00109_),
    .B(_00112_),
    .C(_00116_),
    .Y(_00117_));
 sky130_fd_sc_hd__nand2_1 _06147_ (.A(_00115_),
    .B(_00117_),
    .Y(_00118_));
 sky130_fd_sc_hd__a21oi_2 _06148_ (.A1(_04885_),
    .A2(_04889_),
    .B1(_04883_),
    .Y(_00119_));
 sky130_fd_sc_hd__inv_2 _06149_ (.A(_00119_),
    .Y(_00120_));
 sky130_fd_sc_hd__nand2_1 _06150_ (.A(_00118_),
    .B(_00120_),
    .Y(_00121_));
 sky130_fd_sc_hd__nand3_1 _06151_ (.A(_00115_),
    .B(_00119_),
    .C(_00117_),
    .Y(_00122_));
 sky130_fd_sc_hd__nand2_1 _06152_ (.A(_00121_),
    .B(_00122_),
    .Y(_00123_));
 sky130_fd_sc_hd__clkbuf_4 _06153_ (.A(net47),
    .X(_00124_));
 sky130_fd_sc_hd__nand2_1 _06154_ (.A(_00124_),
    .B(net1),
    .Y(_00125_));
 sky130_fd_sc_hd__nand2_1 _06155_ (.A(net46),
    .B(_04911_),
    .Y(_00126_));
 sky130_fd_sc_hd__nor2_1 _06156_ (.A(_00125_),
    .B(_00126_),
    .Y(_00127_));
 sky130_fd_sc_hd__inv_2 _06157_ (.A(_00127_),
    .Y(_00128_));
 sky130_fd_sc_hd__nand2_1 _06158_ (.A(_00125_),
    .B(_00126_),
    .Y(_00129_));
 sky130_fd_sc_hd__nand2_1 _06159_ (.A(_00128_),
    .B(_00129_),
    .Y(_00130_));
 sky130_fd_sc_hd__inv_2 _06160_ (.A(_00130_),
    .Y(_00131_));
 sky130_fd_sc_hd__nand2_1 _06161_ (.A(_00123_),
    .B(_00131_),
    .Y(_00132_));
 sky130_fd_sc_hd__nand3_1 _06162_ (.A(_00121_),
    .B(_00122_),
    .C(_00130_),
    .Y(_00133_));
 sky130_fd_sc_hd__nand2_1 _06163_ (.A(_00132_),
    .B(_00133_),
    .Y(_00134_));
 sky130_fd_sc_hd__inv_2 _06164_ (.A(_00134_),
    .Y(_00135_));
 sky130_fd_sc_hd__nand2_1 _06165_ (.A(_00107_),
    .B(_00135_),
    .Y(_00136_));
 sky130_fd_sc_hd__nand3_1 _06166_ (.A(_00103_),
    .B(_00106_),
    .C(_00134_),
    .Y(_00137_));
 sky130_fd_sc_hd__nand2_1 _06167_ (.A(_00136_),
    .B(_00137_),
    .Y(_00138_));
 sky130_fd_sc_hd__nand2_1 _06168_ (.A(_04786_),
    .B(_04750_),
    .Y(_00139_));
 sky130_fd_sc_hd__nor2_1 _06169_ (.A(_04750_),
    .B(_04786_),
    .Y(_00140_));
 sky130_fd_sc_hd__a21oi_4 _06170_ (.A1(_00139_),
    .A2(_04790_),
    .B1(_00140_),
    .Y(_00141_));
 sky130_fd_sc_hd__inv_2 _06171_ (.A(_00141_),
    .Y(_00142_));
 sky130_fd_sc_hd__nand2_1 _06172_ (.A(_00138_),
    .B(_00142_),
    .Y(_00143_));
 sky130_fd_sc_hd__nand3_1 _06173_ (.A(_00141_),
    .B(_00136_),
    .C(_00137_),
    .Y(_00144_));
 sky130_fd_sc_hd__nand2_1 _06174_ (.A(_00143_),
    .B(_00144_),
    .Y(_00145_));
 sky130_fd_sc_hd__or2_1 _06175_ (.A(_04839_),
    .B(_04863_),
    .X(_00146_));
 sky130_fd_sc_hd__nand2_1 _06176_ (.A(_04901_),
    .B(_00146_),
    .Y(_00147_));
 sky130_fd_sc_hd__nand2_1 _06177_ (.A(_00145_),
    .B(_00147_),
    .Y(_00148_));
 sky130_fd_sc_hd__inv_2 _06178_ (.A(_00147_),
    .Y(_00149_));
 sky130_fd_sc_hd__nand3_1 _06179_ (.A(_00143_),
    .B(_00144_),
    .C(_00149_),
    .Y(_00150_));
 sky130_fd_sc_hd__nand2_1 _06180_ (.A(_00148_),
    .B(_00150_),
    .Y(_00151_));
 sky130_fd_sc_hd__inv_2 _06181_ (.A(_00151_),
    .Y(_00152_));
 sky130_fd_sc_hd__nand2_1 _06182_ (.A(_00077_),
    .B(_00152_),
    .Y(_00153_));
 sky130_fd_sc_hd__nand3_1 _06183_ (.A(_00073_),
    .B(_00076_),
    .C(_00151_),
    .Y(_00154_));
 sky130_fd_sc_hd__nand3_1 _06184_ (.A(_05151_),
    .B(_00153_),
    .C(_00154_),
    .Y(_00155_));
 sky130_fd_sc_hd__and2_1 _06185_ (.A(_04898_),
    .B(_04891_),
    .X(_00156_));
 sky130_fd_sc_hd__or2_1 _06186_ (.A(_04906_),
    .B(_04903_),
    .X(_00157_));
 sky130_fd_sc_hd__and2_1 _06187_ (.A(_04953_),
    .B(_00157_),
    .X(_00158_));
 sky130_fd_sc_hd__nor2_1 _06188_ (.A(_00156_),
    .B(_00158_),
    .Y(_00159_));
 sky130_fd_sc_hd__inv_2 _06189_ (.A(_00159_),
    .Y(_00160_));
 sky130_fd_sc_hd__nand2_1 _06190_ (.A(_00158_),
    .B(_00156_),
    .Y(_00161_));
 sky130_fd_sc_hd__nand2_1 _06191_ (.A(_00160_),
    .B(_00161_),
    .Y(_00162_));
 sky130_fd_sc_hd__inv_2 _06192_ (.A(_00162_),
    .Y(_00163_));
 sky130_fd_sc_hd__nand2_1 _06193_ (.A(_00153_),
    .B(_00154_),
    .Y(_00164_));
 sky130_fd_sc_hd__a21oi_1 _06194_ (.A1(_05149_),
    .A2(_04956_),
    .B1(_05150_),
    .Y(_00165_));
 sky130_fd_sc_hd__nand2_1 _06195_ (.A(_00164_),
    .B(_00165_),
    .Y(_00166_));
 sky130_fd_sc_hd__nand3_1 _06196_ (.A(_00155_),
    .B(_00163_),
    .C(_00166_),
    .Y(_00167_));
 sky130_fd_sc_hd__nand2_1 _06197_ (.A(_00164_),
    .B(_05151_),
    .Y(_00168_));
 sky130_fd_sc_hd__nand3_1 _06198_ (.A(_00165_),
    .B(_00153_),
    .C(_00154_),
    .Y(_00169_));
 sky130_fd_sc_hd__nand3_1 _06199_ (.A(_00168_),
    .B(_00169_),
    .C(_00162_),
    .Y(_00170_));
 sky130_fd_sc_hd__nand3_1 _06200_ (.A(_05148_),
    .B(_00167_),
    .C(_00170_),
    .Y(_00171_));
 sky130_fd_sc_hd__nand2_1 _06201_ (.A(_00167_),
    .B(_00170_),
    .Y(_00172_));
 sky130_fd_sc_hd__a21o_1 _06202_ (.A1(_05144_),
    .A2(_05146_),
    .B1(_05147_),
    .X(_00173_));
 sky130_fd_sc_hd__nand2_1 _06203_ (.A(_00172_),
    .B(_00173_),
    .Y(_00174_));
 sky130_fd_sc_hd__nand2_1 _06204_ (.A(_00171_),
    .B(_00174_),
    .Y(_00175_));
 sky130_fd_sc_hd__nor2_1 _06205_ (.A(_04916_),
    .B(_05145_),
    .Y(_00176_));
 sky130_fd_sc_hd__nand2_1 _06206_ (.A(_00175_),
    .B(_00176_),
    .Y(_00177_));
 sky130_fd_sc_hd__inv_2 _06207_ (.A(_00176_),
    .Y(_00178_));
 sky130_fd_sc_hd__nand3_2 _06208_ (.A(_00171_),
    .B(_00174_),
    .C(_00178_),
    .Y(_00179_));
 sky130_fd_sc_hd__inv_2 _06209_ (.A(_05141_),
    .Y(_00180_));
 sky130_fd_sc_hd__o21ai_1 _06210_ (.A1(_05142_),
    .A2(_00180_),
    .B1(_05072_),
    .Y(_00181_));
 sky130_fd_sc_hd__nand3b_1 _06211_ (.A_N(_05142_),
    .B(_05073_),
    .C(_05141_),
    .Y(_00182_));
 sky130_fd_sc_hd__nand2_1 _06212_ (.A(_00181_),
    .B(_00182_),
    .Y(_00183_));
 sky130_fd_sc_hd__nand2b_1 _06213_ (.A_N(_04988_),
    .B(_04983_),
    .Y(_00184_));
 sky130_fd_sc_hd__nand3_1 _06214_ (.A(_04971_),
    .B(_04982_),
    .C(_04980_),
    .Y(_00185_));
 sky130_fd_sc_hd__nand2_1 _06215_ (.A(_00185_),
    .B(_04982_),
    .Y(_00186_));
 sky130_fd_sc_hd__nand2_1 _06216_ (.A(_00186_),
    .B(_04988_),
    .Y(_00187_));
 sky130_fd_sc_hd__nand3b_1 _06217_ (.A_N(_04994_),
    .B(_00184_),
    .C(_00187_),
    .Y(_00188_));
 sky130_fd_sc_hd__nand2_1 _06218_ (.A(_00188_),
    .B(_04996_),
    .Y(_00189_));
 sky130_fd_sc_hd__nand3_1 _06219_ (.A(_05047_),
    .B(_05048_),
    .C(_05053_),
    .Y(_00190_));
 sky130_fd_sc_hd__nand2_1 _06220_ (.A(_05055_),
    .B(_00190_),
    .Y(_00191_));
 sky130_fd_sc_hd__nand2_1 _06221_ (.A(_05016_),
    .B(_05017_),
    .Y(_00192_));
 sky130_fd_sc_hd__nand2_1 _06222_ (.A(_05018_),
    .B(_05015_),
    .Y(_00193_));
 sky130_fd_sc_hd__nand3_1 _06223_ (.A(_00192_),
    .B(_00193_),
    .C(_05020_),
    .Y(_00194_));
 sky130_fd_sc_hd__nand2_1 _06224_ (.A(_00194_),
    .B(_05023_),
    .Y(_00195_));
 sky130_fd_sc_hd__nand2_1 _06225_ (.A(_01873_),
    .B(_04260_),
    .Y(_00196_));
 sky130_fd_sc_hd__nand2_1 _06226_ (.A(_02544_),
    .B(_04293_),
    .Y(_00197_));
 sky130_fd_sc_hd__nand2_1 _06227_ (.A(_00196_),
    .B(_00197_),
    .Y(_00198_));
 sky130_fd_sc_hd__nand2_1 _06228_ (.A(_02049_),
    .B(_01158_),
    .Y(_00199_));
 sky130_fd_sc_hd__inv_2 _06229_ (.A(_00199_),
    .Y(_00200_));
 sky130_fd_sc_hd__nor2_1 _06230_ (.A(_00196_),
    .B(_00197_),
    .Y(_00201_));
 sky130_fd_sc_hd__a21oi_2 _06231_ (.A1(_00198_),
    .A2(_00200_),
    .B1(_00201_),
    .Y(_00202_));
 sky130_fd_sc_hd__nand2_1 _06232_ (.A(_00195_),
    .B(_00202_),
    .Y(_00203_));
 sky130_fd_sc_hd__buf_6 _06233_ (.A(_01807_),
    .X(_00204_));
 sky130_fd_sc_hd__nand2_1 _06234_ (.A(_03160_),
    .B(_00204_),
    .Y(_00205_));
 sky130_fd_sc_hd__inv_2 _06235_ (.A(_00205_),
    .Y(_00206_));
 sky130_fd_sc_hd__nand2_1 _06236_ (.A(_03182_),
    .B(_01774_),
    .Y(_00207_));
 sky130_fd_sc_hd__inv_2 _06237_ (.A(_00207_),
    .Y(_00208_));
 sky130_fd_sc_hd__nand2_1 _06238_ (.A(_00206_),
    .B(_00208_),
    .Y(_00209_));
 sky130_fd_sc_hd__nand2_1 _06239_ (.A(_05031_),
    .B(_01884_),
    .Y(_00210_));
 sky130_fd_sc_hd__inv_2 _06240_ (.A(_00210_),
    .Y(_00211_));
 sky130_fd_sc_hd__nand2_1 _06241_ (.A(_00205_),
    .B(_00207_),
    .Y(_00212_));
 sky130_fd_sc_hd__nand3_1 _06242_ (.A(_00209_),
    .B(_00211_),
    .C(_00212_),
    .Y(_00213_));
 sky130_fd_sc_hd__nand2_1 _06243_ (.A(_00213_),
    .B(_00209_),
    .Y(_00214_));
 sky130_fd_sc_hd__nor2_1 _06244_ (.A(_00202_),
    .B(_00195_),
    .Y(_00215_));
 sky130_fd_sc_hd__a21oi_2 _06245_ (.A1(_00203_),
    .A2(_00214_),
    .B1(_00215_),
    .Y(_00216_));
 sky130_fd_sc_hd__nand2_1 _06246_ (.A(_00191_),
    .B(_00216_),
    .Y(_00217_));
 sky130_fd_sc_hd__nand2_1 _06247_ (.A(_04928_),
    .B(_05029_),
    .Y(_00218_));
 sky130_fd_sc_hd__nand2_2 _06248_ (.A(_05028_),
    .B(_05032_),
    .Y(_00219_));
 sky130_fd_sc_hd__nand2_1 _06249_ (.A(_00218_),
    .B(_00219_),
    .Y(_00220_));
 sky130_fd_sc_hd__nand2_1 _06250_ (.A(net35),
    .B(_03820_),
    .Y(_00221_));
 sky130_fd_sc_hd__inv_2 _06251_ (.A(_00221_),
    .Y(_00222_));
 sky130_fd_sc_hd__nor2_1 _06252_ (.A(_00218_),
    .B(_00219_),
    .Y(_00223_));
 sky130_fd_sc_hd__a21oi_2 _06253_ (.A1(_00220_),
    .A2(_00222_),
    .B1(_00223_),
    .Y(_00224_));
 sky130_fd_sc_hd__inv_2 _06254_ (.A(_05030_),
    .Y(_00225_));
 sky130_fd_sc_hd__nand2_1 _06255_ (.A(_00225_),
    .B(_05033_),
    .Y(_00226_));
 sky130_fd_sc_hd__inv_2 _06256_ (.A(_05033_),
    .Y(_00227_));
 sky130_fd_sc_hd__nand2_1 _06257_ (.A(_00227_),
    .B(_05030_),
    .Y(_00228_));
 sky130_fd_sc_hd__nand3_1 _06258_ (.A(_00226_),
    .B(_00228_),
    .C(_05035_),
    .Y(_00229_));
 sky130_fd_sc_hd__nand2_1 _06259_ (.A(_00225_),
    .B(_00227_),
    .Y(_00230_));
 sky130_fd_sc_hd__nand3_1 _06260_ (.A(_00230_),
    .B(_05036_),
    .C(_05034_),
    .Y(_00231_));
 sky130_fd_sc_hd__nand2_1 _06261_ (.A(_00229_),
    .B(_00231_),
    .Y(_00232_));
 sky130_fd_sc_hd__inv_2 _06262_ (.A(_00224_),
    .Y(_00233_));
 sky130_fd_sc_hd__nand2_1 _06263_ (.A(_00232_),
    .B(_00233_),
    .Y(_00234_));
 sky130_fd_sc_hd__nand3_1 _06264_ (.A(_00224_),
    .B(_00229_),
    .C(_00231_),
    .Y(_00235_));
 sky130_fd_sc_hd__nand2_1 _06265_ (.A(_00234_),
    .B(_00235_),
    .Y(_00236_));
 sky130_fd_sc_hd__inv_2 _06266_ (.A(_04966_),
    .Y(_00237_));
 sky130_fd_sc_hd__o21ai_1 _06267_ (.A1(_04969_),
    .A2(_00237_),
    .B1(_04967_),
    .Y(_00238_));
 sky130_fd_sc_hd__nand3b_1 _06268_ (.A_N(_04969_),
    .B(_04968_),
    .C(_04966_),
    .Y(_00239_));
 sky130_fd_sc_hd__nand2_1 _06269_ (.A(_00238_),
    .B(_00239_),
    .Y(_00240_));
 sky130_fd_sc_hd__inv_2 _06270_ (.A(_00240_),
    .Y(_00241_));
 sky130_fd_sc_hd__nand2_1 _06271_ (.A(_00236_),
    .B(_00241_),
    .Y(_00242_));
 sky130_fd_sc_hd__o21ai_2 _06272_ (.A1(_00224_),
    .A2(_00232_),
    .B1(_00242_),
    .Y(_00243_));
 sky130_fd_sc_hd__nor2_1 _06273_ (.A(_00216_),
    .B(_00191_),
    .Y(_00244_));
 sky130_fd_sc_hd__a21oi_2 _06274_ (.A1(_00217_),
    .A2(_00243_),
    .B1(_00244_),
    .Y(_00245_));
 sky130_fd_sc_hd__inv_2 _06275_ (.A(_00245_),
    .Y(_00246_));
 sky130_fd_sc_hd__nand2_1 _06276_ (.A(_00189_),
    .B(_00246_),
    .Y(_00247_));
 sky130_fd_sc_hd__nand3_1 _06277_ (.A(_00188_),
    .B(_04996_),
    .C(_00245_),
    .Y(_00248_));
 sky130_fd_sc_hd__nand2_1 _06278_ (.A(_00247_),
    .B(_00248_),
    .Y(_00249_));
 sky130_fd_sc_hd__nand2_1 _06279_ (.A(_04977_),
    .B(_04978_),
    .Y(_00250_));
 sky130_fd_sc_hd__nand2_1 _06280_ (.A(_00250_),
    .B(_04972_),
    .Y(_00251_));
 sky130_fd_sc_hd__nand2_1 _06281_ (.A(_00251_),
    .B(_04979_),
    .Y(_00252_));
 sky130_fd_sc_hd__nand2_1 _06282_ (.A(_04962_),
    .B(_04819_),
    .Y(_00253_));
 sky130_fd_sc_hd__clkbuf_8 _06283_ (.A(_04809_),
    .X(_00254_));
 sky130_fd_sc_hd__nand2_1 _06284_ (.A(_04964_),
    .B(_00254_),
    .Y(_00255_));
 sky130_fd_sc_hd__nand2_1 _06285_ (.A(_00253_),
    .B(_00255_),
    .Y(_00256_));
 sky130_fd_sc_hd__nand2_1 _06286_ (.A(_03809_),
    .B(_04827_),
    .Y(_00257_));
 sky130_fd_sc_hd__inv_2 _06287_ (.A(_00257_),
    .Y(_00258_));
 sky130_fd_sc_hd__nor2_1 _06288_ (.A(_00253_),
    .B(_00255_),
    .Y(_00259_));
 sky130_fd_sc_hd__a21o_1 _06289_ (.A1(_00256_),
    .A2(_00258_),
    .B1(_00259_),
    .X(_00260_));
 sky130_fd_sc_hd__inv_2 _06290_ (.A(_00260_),
    .Y(_00261_));
 sky130_fd_sc_hd__nand2_1 _06291_ (.A(_00252_),
    .B(_00261_),
    .Y(_00262_));
 sky130_fd_sc_hd__inv_2 _06292_ (.A(_04812_),
    .Y(_00263_));
 sky130_fd_sc_hd__inv_2 _06293_ (.A(_04911_),
    .Y(_00264_));
 sky130_fd_sc_hd__nand2_1 _06294_ (.A(_04808_),
    .B(_04895_),
    .Y(_00265_));
 sky130_fd_sc_hd__nor3_1 _06295_ (.A(_00263_),
    .B(_00264_),
    .C(_00265_),
    .Y(_00266_));
 sky130_fd_sc_hd__nand3_2 _06296_ (.A(_00260_),
    .B(_04979_),
    .C(_00251_),
    .Y(_00267_));
 sky130_fd_sc_hd__a21boi_1 _06297_ (.A1(_00262_),
    .A2(_00266_),
    .B1_N(_00267_),
    .Y(_00268_));
 sky130_fd_sc_hd__nand2_1 _06298_ (.A(_04971_),
    .B(_04982_),
    .Y(_00269_));
 sky130_fd_sc_hd__and2_1 _06299_ (.A(_04979_),
    .B(_04977_),
    .X(_00270_));
 sky130_fd_sc_hd__nand2_1 _06300_ (.A(_00269_),
    .B(_00270_),
    .Y(_00271_));
 sky130_fd_sc_hd__nand2_1 _06301_ (.A(_00271_),
    .B(_00185_),
    .Y(_00272_));
 sky130_fd_sc_hd__nand3_1 _06302_ (.A(_00268_),
    .B(_00185_),
    .C(_00271_),
    .Y(_00273_));
 sky130_fd_sc_hd__nand3_1 _06303_ (.A(_00262_),
    .B(_00267_),
    .C(_00266_),
    .Y(_00274_));
 sky130_fd_sc_hd__nand2_1 _06304_ (.A(_00274_),
    .B(_00267_),
    .Y(_00275_));
 sky130_fd_sc_hd__nand2_1 _06305_ (.A(_00272_),
    .B(_00275_),
    .Y(_00276_));
 sky130_fd_sc_hd__nand2_1 _06306_ (.A(_00273_),
    .B(_00276_),
    .Y(_00277_));
 sky130_fd_sc_hd__nand2_1 _06307_ (.A(_04873_),
    .B(_04992_),
    .Y(_00278_));
 sky130_fd_sc_hd__inv_2 _06308_ (.A(_00278_),
    .Y(_00279_));
 sky130_fd_sc_hd__nand2_1 _06309_ (.A(_00277_),
    .B(_00279_),
    .Y(_00280_));
 sky130_fd_sc_hd__o21ai_1 _06310_ (.A1(_00268_),
    .A2(_00272_),
    .B1(_00280_),
    .Y(_00281_));
 sky130_fd_sc_hd__nand2_1 _06311_ (.A(_00249_),
    .B(_00281_),
    .Y(_00282_));
 sky130_fd_sc_hd__inv_2 _06312_ (.A(_00281_),
    .Y(_00283_));
 sky130_fd_sc_hd__nand3_1 _06313_ (.A(_00247_),
    .B(_00283_),
    .C(_00248_),
    .Y(_00284_));
 sky130_fd_sc_hd__nand2_1 _06314_ (.A(_00282_),
    .B(_00284_),
    .Y(_00285_));
 sky130_fd_sc_hd__inv_2 _06315_ (.A(_00285_),
    .Y(_00286_));
 sky130_fd_sc_hd__nand3_1 _06316_ (.A(_05129_),
    .B(_05088_),
    .C(_05089_),
    .Y(_00287_));
 sky130_fd_sc_hd__a21o_1 _06317_ (.A1(_05099_),
    .A2(_05127_),
    .B1(_05128_),
    .X(_00288_));
 sky130_fd_sc_hd__nand2_1 _06318_ (.A(_05090_),
    .B(_00288_),
    .Y(_00289_));
 sky130_fd_sc_hd__nand2_1 _06319_ (.A(_00287_),
    .B(_00289_),
    .Y(_00290_));
 sky130_fd_sc_hd__nand2_1 _06320_ (.A(_00290_),
    .B(_05138_),
    .Y(_00291_));
 sky130_fd_sc_hd__nand3_1 _06321_ (.A(_00287_),
    .B(_00289_),
    .C(_05137_),
    .Y(_00292_));
 sky130_fd_sc_hd__nand2_1 _06322_ (.A(_00291_),
    .B(_00292_),
    .Y(_00293_));
 sky130_fd_sc_hd__inv_2 _06323_ (.A(_05118_),
    .Y(_00294_));
 sky130_fd_sc_hd__nand3_1 _06324_ (.A(_00294_),
    .B(_05110_),
    .C(_05108_),
    .Y(_00295_));
 sky130_fd_sc_hd__nand3_1 _06325_ (.A(_00295_),
    .B(_05119_),
    .C(_05124_),
    .Y(_00296_));
 sky130_fd_sc_hd__nand2_1 _06326_ (.A(_00296_),
    .B(_00295_),
    .Y(_00297_));
 sky130_fd_sc_hd__nand2_1 _06327_ (.A(_05103_),
    .B(_00297_),
    .Y(_00298_));
 sky130_fd_sc_hd__nand3_1 _06328_ (.A(_05126_),
    .B(_05084_),
    .C(_05102_),
    .Y(_00299_));
 sky130_fd_sc_hd__nand2_1 _06329_ (.A(_00298_),
    .B(_00299_),
    .Y(_00300_));
 sky130_fd_sc_hd__nand2_1 _06330_ (.A(_00300_),
    .B(_05099_),
    .Y(_00301_));
 sky130_fd_sc_hd__nand3_1 _06331_ (.A(_00298_),
    .B(_00299_),
    .C(_05098_),
    .Y(_00302_));
 sky130_fd_sc_hd__nand2_1 _06332_ (.A(_00301_),
    .B(_00302_),
    .Y(_00303_));
 sky130_fd_sc_hd__nand2_1 _06333_ (.A(_05111_),
    .B(_00294_),
    .Y(_00304_));
 sky130_fd_sc_hd__nand3_1 _06334_ (.A(_05118_),
    .B(_05108_),
    .C(_05110_),
    .Y(_00305_));
 sky130_fd_sc_hd__nand3_1 _06335_ (.A(_00304_),
    .B(_00305_),
    .C(_05123_),
    .Y(_00306_));
 sky130_fd_sc_hd__nand2_1 _06336_ (.A(_00296_),
    .B(_00306_),
    .Y(_00307_));
 sky130_fd_sc_hd__inv_2 _06337_ (.A(_05112_),
    .Y(_00308_));
 sky130_fd_sc_hd__nand2_1 _06338_ (.A(_00308_),
    .B(_05113_),
    .Y(_00309_));
 sky130_fd_sc_hd__inv_2 _06339_ (.A(_05113_),
    .Y(_00310_));
 sky130_fd_sc_hd__nand2_1 _06340_ (.A(_00310_),
    .B(_05112_),
    .Y(_00311_));
 sky130_fd_sc_hd__nand3_1 _06341_ (.A(_00309_),
    .B(_00311_),
    .C(_05115_),
    .Y(_00312_));
 sky130_fd_sc_hd__nand2_1 _06342_ (.A(_00308_),
    .B(_00310_),
    .Y(_00313_));
 sky130_fd_sc_hd__nand3_1 _06343_ (.A(_00313_),
    .B(_05116_),
    .C(_05114_),
    .Y(_00314_));
 sky130_fd_sc_hd__nand2_1 _06344_ (.A(_00312_),
    .B(_00314_),
    .Y(_00315_));
 sky130_fd_sc_hd__nand2_2 _06345_ (.A(_01147_),
    .B(_02357_),
    .Y(_00316_));
 sky130_fd_sc_hd__nand2_1 _06346_ (.A(_01037_),
    .B(_02379_),
    .Y(_00317_));
 sky130_fd_sc_hd__nand2_1 _06347_ (.A(_00316_),
    .B(_00317_),
    .Y(_00318_));
 sky130_fd_sc_hd__nand2_1 _06348_ (.A(_02544_),
    .B(_00861_),
    .Y(_00319_));
 sky130_fd_sc_hd__inv_2 _06349_ (.A(_00319_),
    .Y(_00320_));
 sky130_fd_sc_hd__nor2_1 _06350_ (.A(_00316_),
    .B(_00317_),
    .Y(_00321_));
 sky130_fd_sc_hd__a21oi_2 _06351_ (.A1(_00318_),
    .A2(_00320_),
    .B1(_00321_),
    .Y(_00322_));
 sky130_fd_sc_hd__nand2_1 _06352_ (.A(_00315_),
    .B(_00322_),
    .Y(_00323_));
 sky130_fd_sc_hd__inv_2 _06353_ (.A(_00196_),
    .Y(_00324_));
 sky130_fd_sc_hd__inv_2 _06354_ (.A(_00197_),
    .Y(_00325_));
 sky130_fd_sc_hd__nand2_1 _06355_ (.A(_00324_),
    .B(_00325_),
    .Y(_00326_));
 sky130_fd_sc_hd__nand2_1 _06356_ (.A(_00326_),
    .B(_00198_),
    .Y(_00327_));
 sky130_fd_sc_hd__nand2_1 _06357_ (.A(_00327_),
    .B(_00199_),
    .Y(_00328_));
 sky130_fd_sc_hd__nand3_1 _06358_ (.A(_00326_),
    .B(_00200_),
    .C(_00198_),
    .Y(_00329_));
 sky130_fd_sc_hd__nand2_1 _06359_ (.A(_00328_),
    .B(_00329_),
    .Y(_00330_));
 sky130_fd_sc_hd__inv_2 _06360_ (.A(_00330_),
    .Y(_00331_));
 sky130_fd_sc_hd__nor2_1 _06361_ (.A(_00322_),
    .B(_00315_),
    .Y(_00332_));
 sky130_fd_sc_hd__a21oi_1 _06362_ (.A1(_00323_),
    .A2(_00331_),
    .B1(_00332_),
    .Y(_00333_));
 sky130_fd_sc_hd__nand2_1 _06363_ (.A(_00307_),
    .B(_00333_),
    .Y(_00334_));
 sky130_fd_sc_hd__inv_2 _06364_ (.A(_00202_),
    .Y(_00335_));
 sky130_fd_sc_hd__nand2_1 _06365_ (.A(_00195_),
    .B(_00335_),
    .Y(_00336_));
 sky130_fd_sc_hd__nand3_1 _06366_ (.A(_00202_),
    .B(_00194_),
    .C(_05023_),
    .Y(_00337_));
 sky130_fd_sc_hd__nand2_1 _06367_ (.A(_00336_),
    .B(_00337_),
    .Y(_00338_));
 sky130_fd_sc_hd__nand2_1 _06368_ (.A(_00338_),
    .B(_00214_),
    .Y(_00339_));
 sky130_fd_sc_hd__nand3b_1 _06369_ (.A_N(_00214_),
    .B(_00336_),
    .C(_00337_),
    .Y(_00340_));
 sky130_fd_sc_hd__nand2_1 _06370_ (.A(_00339_),
    .B(_00340_),
    .Y(_00341_));
 sky130_fd_sc_hd__inv_2 _06371_ (.A(_00341_),
    .Y(_00342_));
 sky130_fd_sc_hd__nor2_1 _06372_ (.A(_00333_),
    .B(_00307_),
    .Y(_00343_));
 sky130_fd_sc_hd__a21oi_1 _06373_ (.A1(_00334_),
    .A2(_00342_),
    .B1(_00343_),
    .Y(_00344_));
 sky130_fd_sc_hd__nand2_1 _06374_ (.A(_00303_),
    .B(_00344_),
    .Y(_00345_));
 sky130_fd_sc_hd__inv_2 _06375_ (.A(_00216_),
    .Y(_00346_));
 sky130_fd_sc_hd__nand2_1 _06376_ (.A(_00191_),
    .B(_00346_),
    .Y(_00347_));
 sky130_fd_sc_hd__nand3_1 _06377_ (.A(_00216_),
    .B(_05055_),
    .C(_00190_),
    .Y(_00348_));
 sky130_fd_sc_hd__nand3b_1 _06378_ (.A_N(_00243_),
    .B(_00347_),
    .C(_00348_),
    .Y(_00349_));
 sky130_fd_sc_hd__nand2_1 _06379_ (.A(_00347_),
    .B(_00348_),
    .Y(_00350_));
 sky130_fd_sc_hd__nand2_1 _06380_ (.A(_00350_),
    .B(_00243_),
    .Y(_00351_));
 sky130_fd_sc_hd__nand2_1 _06381_ (.A(_00349_),
    .B(_00351_),
    .Y(_00352_));
 sky130_fd_sc_hd__inv_2 _06382_ (.A(_00352_),
    .Y(_00353_));
 sky130_fd_sc_hd__nor2_1 _06383_ (.A(_00344_),
    .B(_00303_),
    .Y(_00354_));
 sky130_fd_sc_hd__a21oi_1 _06384_ (.A1(_00345_),
    .A2(_00353_),
    .B1(_00354_),
    .Y(_00355_));
 sky130_fd_sc_hd__nand2_1 _06385_ (.A(_00293_),
    .B(_00355_),
    .Y(_00356_));
 sky130_fd_sc_hd__nor2_1 _06386_ (.A(_00355_),
    .B(_00293_),
    .Y(_00357_));
 sky130_fd_sc_hd__a21oi_2 _06387_ (.A1(_00286_),
    .A2(_00356_),
    .B1(_00357_),
    .Y(_00358_));
 sky130_fd_sc_hd__nand2_1 _06388_ (.A(_00183_),
    .B(_00358_),
    .Y(_00359_));
 sky130_fd_sc_hd__o21ai_2 _06389_ (.A1(_00189_),
    .A2(_00245_),
    .B1(_00282_),
    .Y(_00360_));
 sky130_fd_sc_hd__nor2_1 _06390_ (.A(_00358_),
    .B(_00183_),
    .Y(_00361_));
 sky130_fd_sc_hd__a21oi_2 _06391_ (.A1(_00359_),
    .A2(_00360_),
    .B1(_00361_),
    .Y(_00362_));
 sky130_fd_sc_hd__inv_2 _06392_ (.A(_05144_),
    .Y(_00363_));
 sky130_fd_sc_hd__o21bai_1 _06393_ (.A1(_05147_),
    .A2(_00363_),
    .B1_N(_05146_),
    .Y(_00364_));
 sky130_fd_sc_hd__nand3b_1 _06394_ (.A_N(_05147_),
    .B(_05146_),
    .C(_05144_),
    .Y(_00365_));
 sky130_fd_sc_hd__nand2_1 _06395_ (.A(_00364_),
    .B(_00365_),
    .Y(_00366_));
 sky130_fd_sc_hd__nor2_1 _06396_ (.A(_00362_),
    .B(_00366_),
    .Y(_00367_));
 sky130_fd_sc_hd__nand3_4 _06397_ (.A(_00177_),
    .B(_00179_),
    .C(_00367_),
    .Y(_00368_));
 sky130_fd_sc_hd__inv_2 _06398_ (.A(_00368_),
    .Y(_00369_));
 sky130_fd_sc_hd__nor2_1 _06399_ (.A(_00165_),
    .B(_00164_),
    .Y(_00370_));
 sky130_fd_sc_hd__a21oi_1 _06400_ (.A1(_00166_),
    .A2(_00163_),
    .B1(_00370_),
    .Y(_00371_));
 sky130_fd_sc_hd__nand2_1 _06401_ (.A(_00074_),
    .B(_05153_),
    .Y(_00372_));
 sky130_fd_sc_hd__nor2_1 _06402_ (.A(_05153_),
    .B(_00074_),
    .Y(_00373_));
 sky130_fd_sc_hd__a21o_1 _06403_ (.A1(_00372_),
    .A2(_00152_),
    .B1(_00373_),
    .X(_00374_));
 sky130_fd_sc_hd__nand2_1 _06404_ (.A(_00069_),
    .B(_00021_),
    .Y(_00375_));
 sky130_fd_sc_hd__nand2_1 _06405_ (.A(_05194_),
    .B(_05157_),
    .Y(_00376_));
 sky130_fd_sc_hd__nor2_1 _06406_ (.A(_05157_),
    .B(_05194_),
    .Y(_00377_));
 sky130_fd_sc_hd__a21o_1 _06407_ (.A1(_00376_),
    .A2(_00018_),
    .B1(_00377_),
    .X(_00378_));
 sky130_fd_sc_hd__nand2_1 _06408_ (.A(_05189_),
    .B(_05175_),
    .Y(_00379_));
 sky130_fd_sc_hd__nand2_1 _06409_ (.A(_00784_),
    .B(_01048_),
    .Y(_00380_));
 sky130_fd_sc_hd__inv_2 _06410_ (.A(_00380_),
    .Y(_00381_));
 sky130_fd_sc_hd__nand3_1 _06411_ (.A(_00381_),
    .B(_01323_),
    .C(_04293_),
    .Y(_00382_));
 sky130_fd_sc_hd__nand2_1 _06412_ (.A(_01323_),
    .B(_04293_),
    .Y(_00383_));
 sky130_fd_sc_hd__nand2_1 _06413_ (.A(_00380_),
    .B(_00383_),
    .Y(_00384_));
 sky130_fd_sc_hd__nand2_1 _06414_ (.A(_00382_),
    .B(_00384_),
    .Y(_00385_));
 sky130_fd_sc_hd__nand2_1 _06415_ (.A(_00740_),
    .B(_01158_),
    .Y(_00386_));
 sky130_fd_sc_hd__nand2_1 _06416_ (.A(_00385_),
    .B(_00386_),
    .Y(_00387_));
 sky130_fd_sc_hd__inv_2 _06417_ (.A(_00386_),
    .Y(_00388_));
 sky130_fd_sc_hd__nand3_1 _06418_ (.A(_00382_),
    .B(_00388_),
    .C(_00384_),
    .Y(_00389_));
 sky130_fd_sc_hd__nand2_1 _06419_ (.A(_00387_),
    .B(_00389_),
    .Y(_00390_));
 sky130_fd_sc_hd__nand2_1 _06420_ (.A(_00751_),
    .B(_05160_),
    .Y(_00391_));
 sky130_fd_sc_hd__inv_2 _06421_ (.A(_00391_),
    .Y(_00392_));
 sky130_fd_sc_hd__clkbuf_4 _06422_ (.A(net16),
    .X(_00393_));
 sky130_fd_sc_hd__nand2_1 _06423_ (.A(_00795_),
    .B(_00393_),
    .Y(_00394_));
 sky130_fd_sc_hd__inv_2 _06424_ (.A(_00394_),
    .Y(_00395_));
 sky130_fd_sc_hd__nand2_1 _06425_ (.A(_00392_),
    .B(_00395_),
    .Y(_00396_));
 sky130_fd_sc_hd__nand2_1 _06426_ (.A(_00391_),
    .B(_00394_),
    .Y(_00397_));
 sky130_fd_sc_hd__nand2_1 _06427_ (.A(_00396_),
    .B(_00397_),
    .Y(_00398_));
 sky130_fd_sc_hd__nand2_1 _06428_ (.A(_00861_),
    .B(_04084_),
    .Y(_00399_));
 sky130_fd_sc_hd__nand2_1 _06429_ (.A(_00398_),
    .B(_00399_),
    .Y(_00400_));
 sky130_fd_sc_hd__nand3b_1 _06430_ (.A_N(_00399_),
    .B(_00396_),
    .C(_00397_),
    .Y(_00401_));
 sky130_fd_sc_hd__nand2_1 _06431_ (.A(_00400_),
    .B(_00401_),
    .Y(_00402_));
 sky130_fd_sc_hd__nor2_1 _06432_ (.A(_05158_),
    .B(_05161_),
    .Y(_00403_));
 sky130_fd_sc_hd__a21o_1 _06433_ (.A1(_05164_),
    .A2(_05168_),
    .B1(_00403_),
    .X(_00404_));
 sky130_fd_sc_hd__inv_2 _06434_ (.A(_00404_),
    .Y(_00405_));
 sky130_fd_sc_hd__nand2_1 _06435_ (.A(_00402_),
    .B(_00405_),
    .Y(_00406_));
 sky130_fd_sc_hd__nand3_1 _06436_ (.A(_00404_),
    .B(_00401_),
    .C(_00400_),
    .Y(_00407_));
 sky130_fd_sc_hd__nand3b_1 _06437_ (.A_N(_00390_),
    .B(_00406_),
    .C(_00407_),
    .Y(_00408_));
 sky130_fd_sc_hd__nand2_1 _06438_ (.A(_00406_),
    .B(_00407_),
    .Y(_00409_));
 sky130_fd_sc_hd__nand2_1 _06439_ (.A(_00409_),
    .B(_00390_),
    .Y(_00410_));
 sky130_fd_sc_hd__nand3_1 _06440_ (.A(_00379_),
    .B(_00408_),
    .C(_00410_),
    .Y(_00411_));
 sky130_fd_sc_hd__buf_12 _06441_ (.A(_01774_),
    .X(_00412_));
 sky130_fd_sc_hd__nand2_1 _06442_ (.A(_01081_),
    .B(_00412_),
    .Y(_00413_));
 sky130_fd_sc_hd__nand2_1 _06443_ (.A(_00850_),
    .B(_00204_),
    .Y(_00414_));
 sky130_fd_sc_hd__or2_1 _06444_ (.A(_00413_),
    .B(_00414_),
    .X(_00415_));
 sky130_fd_sc_hd__nand2_1 _06445_ (.A(_00413_),
    .B(_00414_),
    .Y(_00416_));
 sky130_fd_sc_hd__nand2_1 _06446_ (.A(_00415_),
    .B(_00416_),
    .Y(_00417_));
 sky130_fd_sc_hd__nand2_1 _06447_ (.A(_01037_),
    .B(_00003_),
    .Y(_00418_));
 sky130_fd_sc_hd__nand2_1 _06448_ (.A(_00417_),
    .B(_00418_),
    .Y(_00419_));
 sky130_fd_sc_hd__nand3b_1 _06449_ (.A_N(_00418_),
    .B(_00415_),
    .C(_00416_),
    .Y(_00420_));
 sky130_fd_sc_hd__nand2_1 _06450_ (.A(_00419_),
    .B(_00420_),
    .Y(_00421_));
 sky130_fd_sc_hd__inv_2 _06451_ (.A(_05180_),
    .Y(_00422_));
 sky130_fd_sc_hd__a21oi_2 _06452_ (.A1(_05181_),
    .A2(_05185_),
    .B1(_00422_),
    .Y(_00423_));
 sky130_fd_sc_hd__inv_2 _06453_ (.A(_00423_),
    .Y(_00424_));
 sky130_fd_sc_hd__nand2_1 _06454_ (.A(_00421_),
    .B(_00424_),
    .Y(_00425_));
 sky130_fd_sc_hd__nand3_1 _06455_ (.A(_00423_),
    .B(_00419_),
    .C(_00420_),
    .Y(_00426_));
 sky130_fd_sc_hd__nand2_1 _06456_ (.A(_00425_),
    .B(_00426_),
    .Y(_00427_));
 sky130_fd_sc_hd__nand2_2 _06457_ (.A(_00006_),
    .B(_00000_),
    .Y(_00428_));
 sky130_fd_sc_hd__nand2_1 _06458_ (.A(_00427_),
    .B(_00428_),
    .Y(_00429_));
 sky130_fd_sc_hd__nand3b_1 _06459_ (.A_N(_00428_),
    .B(_00425_),
    .C(_00426_),
    .Y(_00430_));
 sky130_fd_sc_hd__nand2_1 _06460_ (.A(_00429_),
    .B(_00430_),
    .Y(_00431_));
 sky130_fd_sc_hd__inv_2 _06461_ (.A(_00431_),
    .Y(_00432_));
 sky130_fd_sc_hd__nand2_1 _06462_ (.A(_00408_),
    .B(_00410_),
    .Y(_00433_));
 sky130_fd_sc_hd__inv_2 _06463_ (.A(_05175_),
    .Y(_00434_));
 sky130_fd_sc_hd__a21oi_1 _06464_ (.A1(_05173_),
    .A2(_05188_),
    .B1(_00434_),
    .Y(_00435_));
 sky130_fd_sc_hd__nand2_1 _06465_ (.A(_00433_),
    .B(_00435_),
    .Y(_00436_));
 sky130_fd_sc_hd__nand3_2 _06466_ (.A(_00411_),
    .B(_00432_),
    .C(_00436_),
    .Y(_00437_));
 sky130_fd_sc_hd__nand3_1 _06467_ (.A(_00435_),
    .B(_00408_),
    .C(_00410_),
    .Y(_00438_));
 sky130_fd_sc_hd__nand2_1 _06468_ (.A(_00433_),
    .B(_00379_),
    .Y(_00439_));
 sky130_fd_sc_hd__nand3_1 _06469_ (.A(_00438_),
    .B(_00439_),
    .C(_00431_),
    .Y(_00440_));
 sky130_fd_sc_hd__nand3_1 _06470_ (.A(_00378_),
    .B(_00437_),
    .C(_00440_),
    .Y(_00441_));
 sky130_fd_sc_hd__nand2_1 _06471_ (.A(_00437_),
    .B(_00440_),
    .Y(_00442_));
 sky130_fd_sc_hd__a21oi_1 _06472_ (.A1(_00376_),
    .A2(_00018_),
    .B1(_00377_),
    .Y(_00443_));
 sky130_fd_sc_hd__nand2_1 _06473_ (.A(_00442_),
    .B(_00443_),
    .Y(_00444_));
 sky130_fd_sc_hd__nand2_1 _06474_ (.A(_02544_),
    .B(_02995_),
    .Y(_00445_));
 sky130_fd_sc_hd__nand2_1 _06475_ (.A(_01147_),
    .B(_03028_),
    .Y(_00446_));
 sky130_fd_sc_hd__or2_1 _06476_ (.A(_00445_),
    .B(_00446_),
    .X(_00447_));
 sky130_fd_sc_hd__nand2_1 _06477_ (.A(_00445_),
    .B(_00446_),
    .Y(_00448_));
 sky130_fd_sc_hd__nand2_1 _06478_ (.A(_00447_),
    .B(_00448_),
    .Y(_00449_));
 sky130_fd_sc_hd__nand2_1 _06479_ (.A(_03215_),
    .B(_01873_),
    .Y(_00450_));
 sky130_fd_sc_hd__nand2_1 _06480_ (.A(_00449_),
    .B(_00450_),
    .Y(_00451_));
 sky130_fd_sc_hd__inv_2 _06481_ (.A(_00450_),
    .Y(_00452_));
 sky130_fd_sc_hd__nand3_2 _06482_ (.A(_00447_),
    .B(_00448_),
    .C(_00452_),
    .Y(_00453_));
 sky130_fd_sc_hd__nand2_1 _06483_ (.A(_00451_),
    .B(_00453_),
    .Y(_00454_));
 sky130_fd_sc_hd__nor2_1 _06484_ (.A(_00039_),
    .B(_00041_),
    .Y(_00455_));
 sky130_fd_sc_hd__a21oi_2 _06485_ (.A1(_00046_),
    .A2(_00045_),
    .B1(_00455_),
    .Y(_00456_));
 sky130_fd_sc_hd__nand2_1 _06486_ (.A(_00454_),
    .B(_00456_),
    .Y(_00457_));
 sky130_fd_sc_hd__nand2_1 _06487_ (.A(_04962_),
    .B(_03160_),
    .Y(_00458_));
 sky130_fd_sc_hd__nand2_1 _06488_ (.A(_04964_),
    .B(_02049_),
    .Y(_00459_));
 sky130_fd_sc_hd__or2_1 _06489_ (.A(_00458_),
    .B(_00459_),
    .X(_00460_));
 sky130_fd_sc_hd__nand2_1 _06490_ (.A(_00458_),
    .B(_00459_),
    .Y(_00461_));
 sky130_fd_sc_hd__nand2_1 _06491_ (.A(_00460_),
    .B(_00461_),
    .Y(_00462_));
 sky130_fd_sc_hd__nand2_1 _06492_ (.A(_03809_),
    .B(_03182_),
    .Y(_00463_));
 sky130_fd_sc_hd__nand2_1 _06493_ (.A(_00462_),
    .B(_00463_),
    .Y(_00464_));
 sky130_fd_sc_hd__nand3b_1 _06494_ (.A_N(_00463_),
    .B(_00460_),
    .C(_00461_),
    .Y(_00465_));
 sky130_fd_sc_hd__nand2_1 _06495_ (.A(_00464_),
    .B(_00465_),
    .Y(_00466_));
 sky130_fd_sc_hd__inv_2 _06496_ (.A(_00466_),
    .Y(_00467_));
 sky130_fd_sc_hd__inv_2 _06497_ (.A(_00456_),
    .Y(_00468_));
 sky130_fd_sc_hd__nand3_1 _06498_ (.A(_00451_),
    .B(_00468_),
    .C(_00453_),
    .Y(_00469_));
 sky130_fd_sc_hd__nand3_1 _06499_ (.A(_00457_),
    .B(_00467_),
    .C(_00469_),
    .Y(_00470_));
 sky130_fd_sc_hd__nand2_1 _06500_ (.A(_00454_),
    .B(_00468_),
    .Y(_00471_));
 sky130_fd_sc_hd__nand3_1 _06501_ (.A(_00451_),
    .B(_00453_),
    .C(_00456_),
    .Y(_00472_));
 sky130_fd_sc_hd__nand3_1 _06502_ (.A(_00471_),
    .B(_00466_),
    .C(_00472_),
    .Y(_00473_));
 sky130_fd_sc_hd__nand2_1 _06503_ (.A(_00470_),
    .B(_00473_),
    .Y(_00474_));
 sky130_fd_sc_hd__nand2_1 _06504_ (.A(_00007_),
    .B(_00009_),
    .Y(_00475_));
 sky130_fd_sc_hd__nor2_1 _06505_ (.A(_00009_),
    .B(_00007_),
    .Y(_00476_));
 sky130_fd_sc_hd__a21oi_2 _06506_ (.A1(_00475_),
    .A2(_00014_),
    .B1(_00476_),
    .Y(_00477_));
 sky130_fd_sc_hd__inv_2 _06507_ (.A(_00477_),
    .Y(_00478_));
 sky130_fd_sc_hd__nand2_1 _06508_ (.A(_00474_),
    .B(_00478_),
    .Y(_00479_));
 sky130_fd_sc_hd__nand3_1 _06509_ (.A(_00477_),
    .B(_00470_),
    .C(_00473_),
    .Y(_00480_));
 sky130_fd_sc_hd__nand2_1 _06510_ (.A(_00479_),
    .B(_00480_),
    .Y(_00481_));
 sky130_fd_sc_hd__nand2_1 _06511_ (.A(_00053_),
    .B(_00050_),
    .Y(_00482_));
 sky130_fd_sc_hd__nand2_1 _06512_ (.A(_00481_),
    .B(_00482_),
    .Y(_00483_));
 sky130_fd_sc_hd__nand3b_1 _06513_ (.A_N(_00482_),
    .B(_00479_),
    .C(_00480_),
    .Y(_00484_));
 sky130_fd_sc_hd__nand2_1 _06514_ (.A(_00483_),
    .B(_00484_),
    .Y(_00485_));
 sky130_fd_sc_hd__inv_2 _06515_ (.A(_00485_),
    .Y(_00486_));
 sky130_fd_sc_hd__nand3_2 _06516_ (.A(_00441_),
    .B(_00444_),
    .C(_00486_),
    .Y(_00487_));
 sky130_fd_sc_hd__nand2_1 _06517_ (.A(_00442_),
    .B(_00378_),
    .Y(_00488_));
 sky130_fd_sc_hd__nand3_1 _06518_ (.A(_00443_),
    .B(_00437_),
    .C(_00440_),
    .Y(_00489_));
 sky130_fd_sc_hd__nand3_1 _06519_ (.A(_00488_),
    .B(_00489_),
    .C(_00485_),
    .Y(_00490_));
 sky130_fd_sc_hd__nand3_1 _06520_ (.A(_00375_),
    .B(_00487_),
    .C(_00490_),
    .Y(_00491_));
 sky130_fd_sc_hd__nand2_1 _06521_ (.A(_04808_),
    .B(_05028_),
    .Y(_00492_));
 sky130_fd_sc_hd__nand2_1 _06522_ (.A(_04812_),
    .B(_05031_),
    .Y(_00493_));
 sky130_fd_sc_hd__or2_1 _06523_ (.A(_00492_),
    .B(_00493_),
    .X(_00494_));
 sky130_fd_sc_hd__nand2_1 _06524_ (.A(_00492_),
    .B(_00493_),
    .Y(_00495_));
 sky130_fd_sc_hd__nand2_1 _06525_ (.A(_00494_),
    .B(_00495_),
    .Y(_00496_));
 sky130_fd_sc_hd__nand2_1 _06526_ (.A(_04818_),
    .B(_04928_),
    .Y(_00497_));
 sky130_fd_sc_hd__nand2_1 _06527_ (.A(_00496_),
    .B(_00497_),
    .Y(_00498_));
 sky130_fd_sc_hd__nand3b_2 _06528_ (.A_N(_00497_),
    .B(_00494_),
    .C(_00495_),
    .Y(_00499_));
 sky130_fd_sc_hd__nand2_1 _06529_ (.A(_00498_),
    .B(_00499_),
    .Y(_00500_));
 sky130_fd_sc_hd__a21oi_2 _06530_ (.A1(_00029_),
    .A2(_00033_),
    .B1(_00027_),
    .Y(_00501_));
 sky130_fd_sc_hd__nand2_1 _06531_ (.A(_00500_),
    .B(_00501_),
    .Y(_00502_));
 sky130_fd_sc_hd__inv_2 _06532_ (.A(_00501_),
    .Y(_00503_));
 sky130_fd_sc_hd__nand3_1 _06533_ (.A(_00498_),
    .B(_00499_),
    .C(_00503_),
    .Y(_00504_));
 sky130_fd_sc_hd__nand2_1 _06534_ (.A(_00090_),
    .B(_00084_),
    .Y(_00505_));
 sky130_fd_sc_hd__nand3_1 _06535_ (.A(_00502_),
    .B(_00504_),
    .C(_00505_),
    .Y(_00506_));
 sky130_fd_sc_hd__nand2_1 _06536_ (.A(_00500_),
    .B(_00503_),
    .Y(_00507_));
 sky130_fd_sc_hd__nand3_1 _06537_ (.A(_00498_),
    .B(_00499_),
    .C(_00501_),
    .Y(_00508_));
 sky130_fd_sc_hd__inv_2 _06538_ (.A(_00505_),
    .Y(_00509_));
 sky130_fd_sc_hd__nand3_1 _06539_ (.A(_00507_),
    .B(_00508_),
    .C(_00509_),
    .Y(_00510_));
 sky130_fd_sc_hd__nand2_1 _06540_ (.A(_00506_),
    .B(_00510_),
    .Y(_00511_));
 sky130_fd_sc_hd__a21boi_2 _06541_ (.A1(_00097_),
    .A2(_00094_),
    .B1_N(_00096_),
    .Y(_00512_));
 sky130_fd_sc_hd__inv_2 _06542_ (.A(_00512_),
    .Y(_00513_));
 sky130_fd_sc_hd__nand2_1 _06543_ (.A(_00511_),
    .B(_00513_),
    .Y(_00514_));
 sky130_fd_sc_hd__nand3_1 _06544_ (.A(_00512_),
    .B(_00506_),
    .C(_00510_),
    .Y(_00515_));
 sky130_fd_sc_hd__nand2_1 _06545_ (.A(_00514_),
    .B(_00515_),
    .Y(_00516_));
 sky130_fd_sc_hd__nand2_1 _06546_ (.A(_04871_),
    .B(_04809_),
    .Y(_00517_));
 sky130_fd_sc_hd__nand2_1 _06547_ (.A(_04873_),
    .B(_03820_),
    .Y(_00518_));
 sky130_fd_sc_hd__or2_1 _06548_ (.A(_00517_),
    .B(_00518_),
    .X(_00519_));
 sky130_fd_sc_hd__nand2_1 _06549_ (.A(_00517_),
    .B(_00518_),
    .Y(_00520_));
 sky130_fd_sc_hd__nand2_1 _06550_ (.A(_00519_),
    .B(_00520_),
    .Y(_00521_));
 sky130_fd_sc_hd__clkbuf_8 _06551_ (.A(_04819_),
    .X(_00522_));
 sky130_fd_sc_hd__nand2_1 _06552_ (.A(_04876_),
    .B(_00522_),
    .Y(_00523_));
 sky130_fd_sc_hd__nand2_1 _06553_ (.A(_00521_),
    .B(_00523_),
    .Y(_00524_));
 sky130_fd_sc_hd__nand3b_1 _06554_ (.A_N(_00523_),
    .B(_00519_),
    .C(_00520_),
    .Y(_00525_));
 sky130_fd_sc_hd__nand2_1 _06555_ (.A(_00524_),
    .B(_00525_),
    .Y(_00526_));
 sky130_fd_sc_hd__a21boi_2 _06556_ (.A1(_00116_),
    .A2(_00112_),
    .B1_N(_00109_),
    .Y(_00527_));
 sky130_fd_sc_hd__or2_1 _06557_ (.A(_00526_),
    .B(_00527_),
    .X(_00528_));
 sky130_fd_sc_hd__clkbuf_4 _06558_ (.A(net48),
    .X(_00529_));
 sky130_fd_sc_hd__nand2_1 _06559_ (.A(_00529_),
    .B(net1),
    .Y(_00530_));
 sky130_fd_sc_hd__inv_2 _06560_ (.A(_00530_),
    .Y(_00531_));
 sky130_fd_sc_hd__nand2_1 _06561_ (.A(_00124_),
    .B(_04911_),
    .Y(_00532_));
 sky130_fd_sc_hd__nand2_1 _06562_ (.A(net46),
    .B(_04827_),
    .Y(_00533_));
 sky130_fd_sc_hd__or2_1 _06563_ (.A(_00532_),
    .B(_00533_),
    .X(_00534_));
 sky130_fd_sc_hd__nand2_1 _06564_ (.A(_00532_),
    .B(_00533_),
    .Y(_00535_));
 sky130_fd_sc_hd__nand2_1 _06565_ (.A(_00534_),
    .B(_00535_),
    .Y(_00536_));
 sky130_fd_sc_hd__xor2_1 _06566_ (.A(_00531_),
    .B(_00536_),
    .X(_00537_));
 sky130_fd_sc_hd__inv_2 _06567_ (.A(_00537_),
    .Y(_00538_));
 sky130_fd_sc_hd__nand2_1 _06568_ (.A(_00527_),
    .B(_00526_),
    .Y(_00539_));
 sky130_fd_sc_hd__nand3_1 _06569_ (.A(_00528_),
    .B(_00538_),
    .C(_00539_),
    .Y(_00540_));
 sky130_fd_sc_hd__or2b_1 _06570_ (.A(_00527_),
    .B_N(_00526_),
    .X(_00541_));
 sky130_fd_sc_hd__or2b_1 _06571_ (.A(_00526_),
    .B_N(_00527_),
    .X(_00542_));
 sky130_fd_sc_hd__nand3_1 _06572_ (.A(_00541_),
    .B(_00542_),
    .C(_00537_),
    .Y(_00543_));
 sky130_fd_sc_hd__nand2_1 _06573_ (.A(_00540_),
    .B(_00543_),
    .Y(_00544_));
 sky130_fd_sc_hd__inv_2 _06574_ (.A(_00544_),
    .Y(_00545_));
 sky130_fd_sc_hd__nand2_1 _06575_ (.A(_00516_),
    .B(_00545_),
    .Y(_00546_));
 sky130_fd_sc_hd__nand3_1 _06576_ (.A(_00544_),
    .B(_00514_),
    .C(_00515_),
    .Y(_00547_));
 sky130_fd_sc_hd__nand2_1 _06577_ (.A(_00546_),
    .B(_00547_),
    .Y(_00548_));
 sky130_fd_sc_hd__nand2_1 _06578_ (.A(_00057_),
    .B(_00059_),
    .Y(_00549_));
 sky130_fd_sc_hd__nor2_1 _06579_ (.A(_00059_),
    .B(_00057_),
    .Y(_00550_));
 sky130_fd_sc_hd__a21oi_2 _06580_ (.A1(_00549_),
    .A2(_00064_),
    .B1(_00550_),
    .Y(_00551_));
 sky130_fd_sc_hd__inv_2 _06581_ (.A(_00551_),
    .Y(_00552_));
 sky130_fd_sc_hd__nand2_1 _06582_ (.A(_00548_),
    .B(_00552_),
    .Y(_00553_));
 sky130_fd_sc_hd__nand3_1 _06583_ (.A(_00546_),
    .B(_00551_),
    .C(_00547_),
    .Y(_00554_));
 sky130_fd_sc_hd__nand2_1 _06584_ (.A(_00553_),
    .B(_00554_),
    .Y(_00555_));
 sky130_fd_sc_hd__nor2_1 _06585_ (.A(_00079_),
    .B(_00105_),
    .Y(_00556_));
 sky130_fd_sc_hd__inv_2 _06586_ (.A(_00136_),
    .Y(_00557_));
 sky130_fd_sc_hd__nor2_1 _06587_ (.A(_00556_),
    .B(_00557_),
    .Y(_00558_));
 sky130_fd_sc_hd__inv_2 _06588_ (.A(_00558_),
    .Y(_00559_));
 sky130_fd_sc_hd__nand2_1 _06589_ (.A(_00555_),
    .B(_00559_),
    .Y(_00560_));
 sky130_fd_sc_hd__nand3_1 _06590_ (.A(_00553_),
    .B(_00554_),
    .C(_00558_),
    .Y(_00561_));
 sky130_fd_sc_hd__nand2_1 _06591_ (.A(_00560_),
    .B(_00561_),
    .Y(_00562_));
 sky130_fd_sc_hd__inv_2 _06592_ (.A(_00562_),
    .Y(_00563_));
 sky130_fd_sc_hd__nand2_1 _06593_ (.A(_00487_),
    .B(_00490_),
    .Y(_00564_));
 sky130_fd_sc_hd__nor2_1 _06594_ (.A(_00023_),
    .B(_00022_),
    .Y(_00565_));
 sky130_fd_sc_hd__a21oi_1 _06595_ (.A1(_00024_),
    .A2(_00068_),
    .B1(_00565_),
    .Y(_00566_));
 sky130_fd_sc_hd__nand2_1 _06596_ (.A(_00564_),
    .B(_00566_),
    .Y(_00567_));
 sky130_fd_sc_hd__nand3_2 _06597_ (.A(_00491_),
    .B(_00563_),
    .C(_00567_),
    .Y(_00568_));
 sky130_fd_sc_hd__nand3_1 _06598_ (.A(_00566_),
    .B(_00487_),
    .C(_00490_),
    .Y(_00569_));
 sky130_fd_sc_hd__nand2_1 _06599_ (.A(_00564_),
    .B(_00375_),
    .Y(_00570_));
 sky130_fd_sc_hd__nand3_1 _06600_ (.A(_00569_),
    .B(_00570_),
    .C(_00562_),
    .Y(_00571_));
 sky130_fd_sc_hd__nand3_1 _06601_ (.A(_00374_),
    .B(_00568_),
    .C(_00571_),
    .Y(_00572_));
 sky130_fd_sc_hd__o21a_1 _06602_ (.A1(_00119_),
    .A2(_00118_),
    .B1(_00132_),
    .X(_00573_));
 sky130_fd_sc_hd__or2_1 _06603_ (.A(_00128_),
    .B(_00573_),
    .X(_00574_));
 sky130_fd_sc_hd__nand2_1 _06604_ (.A(_00573_),
    .B(_00128_),
    .Y(_00575_));
 sky130_fd_sc_hd__nand2_1 _06605_ (.A(_00574_),
    .B(_00575_),
    .Y(_00576_));
 sky130_fd_sc_hd__o21a_1 _06606_ (.A1(_00138_),
    .A2(_00141_),
    .B1(_00148_),
    .X(_00577_));
 sky130_fd_sc_hd__nor2_2 _06607_ (.A(_00576_),
    .B(_00577_),
    .Y(_00578_));
 sky130_fd_sc_hd__inv_2 _06608_ (.A(_00578_),
    .Y(_00579_));
 sky130_fd_sc_hd__nand2_1 _06609_ (.A(_00577_),
    .B(_00576_),
    .Y(_00580_));
 sky130_fd_sc_hd__nand2_2 _06610_ (.A(_00579_),
    .B(_00580_),
    .Y(_00581_));
 sky130_fd_sc_hd__inv_2 _06611_ (.A(_00581_),
    .Y(_00582_));
 sky130_fd_sc_hd__nand2_1 _06612_ (.A(_00568_),
    .B(_00571_),
    .Y(_00583_));
 sky130_fd_sc_hd__a21oi_1 _06613_ (.A1(_00372_),
    .A2(_00152_),
    .B1(_00373_),
    .Y(_00584_));
 sky130_fd_sc_hd__nand2_1 _06614_ (.A(_00583_),
    .B(_00584_),
    .Y(_00585_));
 sky130_fd_sc_hd__nand3_2 _06615_ (.A(_00572_),
    .B(_00582_),
    .C(_00585_),
    .Y(_00586_));
 sky130_fd_sc_hd__nand2_1 _06616_ (.A(_00583_),
    .B(_00374_),
    .Y(_00587_));
 sky130_fd_sc_hd__nand3_1 _06617_ (.A(_00584_),
    .B(_00568_),
    .C(_00571_),
    .Y(_00588_));
 sky130_fd_sc_hd__nand3_1 _06618_ (.A(_00587_),
    .B(_00588_),
    .C(_00581_),
    .Y(_00589_));
 sky130_fd_sc_hd__nand3_2 _06619_ (.A(_00371_),
    .B(_00586_),
    .C(_00589_),
    .Y(_00590_));
 sky130_fd_sc_hd__nand2_1 _06620_ (.A(_00586_),
    .B(_00589_),
    .Y(_00591_));
 sky130_fd_sc_hd__a21o_1 _06621_ (.A1(_00166_),
    .A2(_00163_),
    .B1(_00370_),
    .X(_00592_));
 sky130_fd_sc_hd__nand2_1 _06622_ (.A(_00591_),
    .B(_00592_),
    .Y(_00593_));
 sky130_fd_sc_hd__nand2_1 _06623_ (.A(_00590_),
    .B(_00593_),
    .Y(_00594_));
 sky130_fd_sc_hd__nand2_1 _06624_ (.A(_00594_),
    .B(_00160_),
    .Y(_00595_));
 sky130_fd_sc_hd__nand3_1 _06625_ (.A(_00590_),
    .B(_00593_),
    .C(_00159_),
    .Y(_00596_));
 sky130_fd_sc_hd__nand2_1 _06626_ (.A(_00595_),
    .B(_00596_),
    .Y(_00597_));
 sky130_fd_sc_hd__nand2_1 _06627_ (.A(_00172_),
    .B(_05148_),
    .Y(_00598_));
 sky130_fd_sc_hd__nor2_1 _06628_ (.A(_05148_),
    .B(_00172_),
    .Y(_00599_));
 sky130_fd_sc_hd__a21oi_2 _06629_ (.A1(_00598_),
    .A2(_00176_),
    .B1(_00599_),
    .Y(_00600_));
 sky130_fd_sc_hd__inv_2 _06630_ (.A(_00600_),
    .Y(_00601_));
 sky130_fd_sc_hd__nand2_2 _06631_ (.A(_00597_),
    .B(_00601_),
    .Y(_00602_));
 sky130_fd_sc_hd__nand3_1 _06632_ (.A(_00600_),
    .B(_00595_),
    .C(_00596_),
    .Y(_00603_));
 sky130_fd_sc_hd__nand3_2 _06633_ (.A(_00369_),
    .B(_00602_),
    .C(_00603_),
    .Y(_00604_));
 sky130_fd_sc_hd__nand2_1 _06634_ (.A(_00594_),
    .B(_00159_),
    .Y(_00605_));
 sky130_fd_sc_hd__nand3_1 _06635_ (.A(_00590_),
    .B(_00593_),
    .C(_00160_),
    .Y(_00606_));
 sky130_fd_sc_hd__nand2_1 _06636_ (.A(_00605_),
    .B(_00606_),
    .Y(_00607_));
 sky130_fd_sc_hd__nand2_1 _06637_ (.A(_00607_),
    .B(_00601_),
    .Y(_00608_));
 sky130_fd_sc_hd__nand3_1 _06638_ (.A(_00600_),
    .B(_00605_),
    .C(_00606_),
    .Y(_00609_));
 sky130_fd_sc_hd__nand3_2 _06639_ (.A(_00608_),
    .B(_00609_),
    .C(_00368_),
    .Y(_00610_));
 sky130_fd_sc_hd__nand2_1 _06640_ (.A(_00604_),
    .B(_00610_),
    .Y(_00611_));
 sky130_fd_sc_hd__nand2_1 _06641_ (.A(_00177_),
    .B(_00179_),
    .Y(_00612_));
 sky130_fd_sc_hd__inv_2 _06642_ (.A(_00362_),
    .Y(_00613_));
 sky130_fd_sc_hd__nand3_2 _06643_ (.A(_00613_),
    .B(_00365_),
    .C(_00364_),
    .Y(_00614_));
 sky130_fd_sc_hd__nand2_2 _06644_ (.A(_00612_),
    .B(_00614_),
    .Y(_00615_));
 sky130_fd_sc_hd__nand2_1 _06645_ (.A(_00615_),
    .B(_00368_),
    .Y(_00616_));
 sky130_fd_sc_hd__nand3_1 _06646_ (.A(_00355_),
    .B(_00291_),
    .C(_00292_),
    .Y(_00617_));
 sky130_fd_sc_hd__a21o_1 _06647_ (.A1(_00334_),
    .A2(_00342_),
    .B1(_00343_),
    .X(_00618_));
 sky130_fd_sc_hd__nand3_1 _06648_ (.A(_00618_),
    .B(_00301_),
    .C(_00302_),
    .Y(_00619_));
 sky130_fd_sc_hd__nand3_1 _06649_ (.A(_00619_),
    .B(_00353_),
    .C(_00345_),
    .Y(_00620_));
 sky130_fd_sc_hd__nand2_1 _06650_ (.A(_00620_),
    .B(_00619_),
    .Y(_00621_));
 sky130_fd_sc_hd__nand2_1 _06651_ (.A(_00293_),
    .B(_00621_),
    .Y(_00622_));
 sky130_fd_sc_hd__nand2_1 _06652_ (.A(_00617_),
    .B(_00622_),
    .Y(_00623_));
 sky130_fd_sc_hd__nand2_1 _06653_ (.A(_00623_),
    .B(_00286_),
    .Y(_00624_));
 sky130_fd_sc_hd__nand3_1 _06654_ (.A(_00285_),
    .B(_00617_),
    .C(_00622_),
    .Y(_00625_));
 sky130_fd_sc_hd__nand2_1 _06655_ (.A(_00624_),
    .B(_00625_),
    .Y(_00626_));
 sky130_fd_sc_hd__nand3_1 _06656_ (.A(_00273_),
    .B(_00276_),
    .C(_00278_),
    .Y(_00627_));
 sky130_fd_sc_hd__nand2_1 _06657_ (.A(_00280_),
    .B(_00627_),
    .Y(_00628_));
 sky130_fd_sc_hd__nand3_1 _06658_ (.A(_00234_),
    .B(_00235_),
    .C(_00240_),
    .Y(_00629_));
 sky130_fd_sc_hd__nand2_1 _06659_ (.A(_00242_),
    .B(_00629_),
    .Y(_00630_));
 sky130_fd_sc_hd__nand2_1 _06660_ (.A(_00208_),
    .B(_00205_),
    .Y(_00631_));
 sky130_fd_sc_hd__nand2_1 _06661_ (.A(_00206_),
    .B(_00207_),
    .Y(_00632_));
 sky130_fd_sc_hd__nand3_1 _06662_ (.A(_00631_),
    .B(_00632_),
    .C(_00210_),
    .Y(_00633_));
 sky130_fd_sc_hd__nand2_1 _06663_ (.A(_00633_),
    .B(_00213_),
    .Y(_00634_));
 sky130_fd_sc_hd__nand2_1 _06664_ (.A(_02049_),
    .B(_04260_),
    .Y(_00635_));
 sky130_fd_sc_hd__nand2_1 _06665_ (.A(_01873_),
    .B(_04293_),
    .Y(_00636_));
 sky130_fd_sc_hd__nand2_1 _06666_ (.A(_00635_),
    .B(_00636_),
    .Y(_00637_));
 sky130_fd_sc_hd__nand2_1 _06667_ (.A(_03160_),
    .B(_01565_),
    .Y(_00638_));
 sky130_fd_sc_hd__inv_2 _06668_ (.A(_00638_),
    .Y(_00639_));
 sky130_fd_sc_hd__nor2_1 _06669_ (.A(_00635_),
    .B(_00636_),
    .Y(_00640_));
 sky130_fd_sc_hd__a21oi_2 _06670_ (.A1(_00637_),
    .A2(_00639_),
    .B1(_00640_),
    .Y(_00641_));
 sky130_fd_sc_hd__nand2_1 _06671_ (.A(_00634_),
    .B(_00641_),
    .Y(_00642_));
 sky130_fd_sc_hd__nand2_1 _06672_ (.A(_05031_),
    .B(_00412_),
    .Y(_00643_));
 sky130_fd_sc_hd__inv_2 _06673_ (.A(_00643_),
    .Y(_00644_));
 sky130_fd_sc_hd__nand2_1 _06674_ (.A(_03182_),
    .B(_00204_),
    .Y(_00645_));
 sky130_fd_sc_hd__inv_2 _06675_ (.A(_00645_),
    .Y(_00646_));
 sky130_fd_sc_hd__nand2_1 _06676_ (.A(_00644_),
    .B(_00646_),
    .Y(_00647_));
 sky130_fd_sc_hd__nand2_1 _06677_ (.A(_05028_),
    .B(_00003_),
    .Y(_00648_));
 sky130_fd_sc_hd__inv_2 _06678_ (.A(_00648_),
    .Y(_00649_));
 sky130_fd_sc_hd__nand2_1 _06679_ (.A(_00643_),
    .B(_00645_),
    .Y(_00650_));
 sky130_fd_sc_hd__nand3_1 _06680_ (.A(_00647_),
    .B(_00649_),
    .C(_00650_),
    .Y(_00651_));
 sky130_fd_sc_hd__nand2_1 _06681_ (.A(_00651_),
    .B(_00647_),
    .Y(_00652_));
 sky130_fd_sc_hd__nor2_1 _06682_ (.A(_00641_),
    .B(_00634_),
    .Y(_00653_));
 sky130_fd_sc_hd__a21oi_2 _06683_ (.A1(_00642_),
    .A2(_00652_),
    .B1(_00653_),
    .Y(_00654_));
 sky130_fd_sc_hd__nand2_1 _06684_ (.A(_00630_),
    .B(_00654_),
    .Y(_00655_));
 sky130_fd_sc_hd__clkbuf_8 _06685_ (.A(_03820_),
    .X(_00656_));
 sky130_fd_sc_hd__nand2_1 _06686_ (.A(_00656_),
    .B(_05029_),
    .Y(_00657_));
 sky130_fd_sc_hd__nand2_1 _06687_ (.A(_04928_),
    .B(_05032_),
    .Y(_00658_));
 sky130_fd_sc_hd__nand2_1 _06688_ (.A(_00657_),
    .B(_00658_),
    .Y(_00659_));
 sky130_fd_sc_hd__nand2_1 _06689_ (.A(_03215_),
    .B(_04809_),
    .Y(_00660_));
 sky130_fd_sc_hd__inv_2 _06690_ (.A(_00660_),
    .Y(_00661_));
 sky130_fd_sc_hd__nor2_1 _06691_ (.A(_00657_),
    .B(_00658_),
    .Y(_00662_));
 sky130_fd_sc_hd__a21oi_2 _06692_ (.A1(_00659_),
    .A2(_00661_),
    .B1(_00662_),
    .Y(_00663_));
 sky130_fd_sc_hd__inv_2 _06693_ (.A(_00219_),
    .Y(_00664_));
 sky130_fd_sc_hd__nand2_1 _06694_ (.A(_00664_),
    .B(_00218_),
    .Y(_00665_));
 sky130_fd_sc_hd__inv_2 _06695_ (.A(_00218_),
    .Y(_00666_));
 sky130_fd_sc_hd__nand2_1 _06696_ (.A(_00666_),
    .B(_00219_),
    .Y(_00667_));
 sky130_fd_sc_hd__nand3_1 _06697_ (.A(_00665_),
    .B(_00667_),
    .C(_00221_),
    .Y(_00668_));
 sky130_fd_sc_hd__nand2_1 _06698_ (.A(_00666_),
    .B(_00664_),
    .Y(_00669_));
 sky130_fd_sc_hd__nand3_1 _06699_ (.A(_00669_),
    .B(_00222_),
    .C(_00220_),
    .Y(_00670_));
 sky130_fd_sc_hd__nand2_1 _06700_ (.A(_00668_),
    .B(_00670_),
    .Y(_00671_));
 sky130_fd_sc_hd__inv_2 _06701_ (.A(_00663_),
    .Y(_00672_));
 sky130_fd_sc_hd__nand2_1 _06702_ (.A(_00671_),
    .B(_00672_),
    .Y(_00673_));
 sky130_fd_sc_hd__nand3_1 _06703_ (.A(_00663_),
    .B(_00668_),
    .C(_00670_),
    .Y(_00674_));
 sky130_fd_sc_hd__nand2_1 _06704_ (.A(_00673_),
    .B(_00674_),
    .Y(_00675_));
 sky130_fd_sc_hd__inv_2 _06705_ (.A(_00256_),
    .Y(_00676_));
 sky130_fd_sc_hd__o21ai_1 _06706_ (.A1(_00259_),
    .A2(_00676_),
    .B1(_00257_),
    .Y(_00677_));
 sky130_fd_sc_hd__nand3b_1 _06707_ (.A_N(_00259_),
    .B(_00258_),
    .C(_00256_),
    .Y(_00678_));
 sky130_fd_sc_hd__nand2_1 _06708_ (.A(_00677_),
    .B(_00678_),
    .Y(_00679_));
 sky130_fd_sc_hd__inv_2 _06709_ (.A(_00679_),
    .Y(_00680_));
 sky130_fd_sc_hd__nand2_1 _06710_ (.A(_00675_),
    .B(_00680_),
    .Y(_00681_));
 sky130_fd_sc_hd__o21ai_1 _06711_ (.A1(_00663_),
    .A2(_00671_),
    .B1(_00681_),
    .Y(_00682_));
 sky130_fd_sc_hd__nor2_1 _06712_ (.A(_00654_),
    .B(_00630_),
    .Y(_00683_));
 sky130_fd_sc_hd__a21o_1 _06713_ (.A1(_00655_),
    .A2(_00682_),
    .B1(_00683_),
    .X(_00684_));
 sky130_fd_sc_hd__inv_2 _06714_ (.A(_00684_),
    .Y(_00685_));
 sky130_fd_sc_hd__nand2_1 _06715_ (.A(_00628_),
    .B(_00685_),
    .Y(_00686_));
 sky130_fd_sc_hd__nand3_1 _06716_ (.A(_00684_),
    .B(_00280_),
    .C(_00627_),
    .Y(_00687_));
 sky130_fd_sc_hd__nand2_1 _06717_ (.A(_00686_),
    .B(_00687_),
    .Y(_00688_));
 sky130_fd_sc_hd__a21o_1 _06718_ (.A1(_00262_),
    .A2(_00267_),
    .B1(_00266_),
    .X(_00689_));
 sky130_fd_sc_hd__o21ai_1 _06719_ (.A1(_00263_),
    .A2(_00264_),
    .B1(_00265_),
    .Y(_00690_));
 sky130_fd_sc_hd__or2b_1 _06720_ (.A(_00266_),
    .B_N(_00690_),
    .X(_00691_));
 sky130_fd_sc_hd__nand2_1 _06721_ (.A(_03809_),
    .B(_04911_),
    .Y(_00692_));
 sky130_fd_sc_hd__nand2_1 _06722_ (.A(_04962_),
    .B(_04828_),
    .Y(_00693_));
 sky130_fd_sc_hd__nand2_1 _06723_ (.A(_04964_),
    .B(_00522_),
    .Y(_00694_));
 sky130_fd_sc_hd__or2_1 _06724_ (.A(_00693_),
    .B(_00694_),
    .X(_00695_));
 sky130_fd_sc_hd__nand2_1 _06725_ (.A(_00693_),
    .B(_00694_),
    .Y(_00696_));
 sky130_fd_sc_hd__nand3b_1 _06726_ (.A_N(_00692_),
    .B(_00695_),
    .C(_00696_),
    .Y(_00697_));
 sky130_fd_sc_hd__and2_1 _06727_ (.A(_00697_),
    .B(_00695_),
    .X(_00698_));
 sky130_fd_sc_hd__nor2_1 _06728_ (.A(_00691_),
    .B(_00698_),
    .Y(_00699_));
 sky130_fd_sc_hd__nand3_2 _06729_ (.A(_00689_),
    .B(_00274_),
    .C(_00699_),
    .Y(_00700_));
 sky130_fd_sc_hd__nand2_1 _06730_ (.A(_00688_),
    .B(_00700_),
    .Y(_00701_));
 sky130_fd_sc_hd__inv_2 _06731_ (.A(_00700_),
    .Y(_00702_));
 sky130_fd_sc_hd__nand3_1 _06732_ (.A(_00686_),
    .B(_00687_),
    .C(_00702_),
    .Y(_00703_));
 sky130_fd_sc_hd__nand2_1 _06733_ (.A(_00701_),
    .B(_00703_),
    .Y(_00704_));
 sky130_fd_sc_hd__inv_2 _06734_ (.A(_00704_),
    .Y(_00705_));
 sky130_fd_sc_hd__nand2_1 _06735_ (.A(_00303_),
    .B(_00618_),
    .Y(_00706_));
 sky130_fd_sc_hd__nand3_1 _06736_ (.A(_00344_),
    .B(_00301_),
    .C(_00302_),
    .Y(_00707_));
 sky130_fd_sc_hd__nand3_1 _06737_ (.A(_00706_),
    .B(_00707_),
    .C(_00352_),
    .Y(_00708_));
 sky130_fd_sc_hd__nand2_1 _06738_ (.A(_00620_),
    .B(_00708_),
    .Y(_00709_));
 sky130_fd_sc_hd__nand3_1 _06739_ (.A(_00333_),
    .B(_00296_),
    .C(_00306_),
    .Y(_00710_));
 sky130_fd_sc_hd__inv_2 _06740_ (.A(_00322_),
    .Y(_00711_));
 sky130_fd_sc_hd__nand3_1 _06741_ (.A(_00711_),
    .B(_00314_),
    .C(_00312_),
    .Y(_00712_));
 sky130_fd_sc_hd__nand3_1 _06742_ (.A(_00712_),
    .B(_00323_),
    .C(_00331_),
    .Y(_00713_));
 sky130_fd_sc_hd__nand2_1 _06743_ (.A(_00713_),
    .B(_00712_),
    .Y(_00714_));
 sky130_fd_sc_hd__nand2_1 _06744_ (.A(_00307_),
    .B(_00714_),
    .Y(_00715_));
 sky130_fd_sc_hd__nand2_1 _06745_ (.A(_00710_),
    .B(_00715_),
    .Y(_00716_));
 sky130_fd_sc_hd__nand2_1 _06746_ (.A(_00716_),
    .B(_00342_),
    .Y(_00717_));
 sky130_fd_sc_hd__nand3_1 _06747_ (.A(_00710_),
    .B(_00715_),
    .C(_00341_),
    .Y(_00718_));
 sky130_fd_sc_hd__nand2_1 _06748_ (.A(_00717_),
    .B(_00718_),
    .Y(_00719_));
 sky130_fd_sc_hd__nand2_1 _06749_ (.A(_00315_),
    .B(_00711_),
    .Y(_00720_));
 sky130_fd_sc_hd__nand3_1 _06750_ (.A(_00322_),
    .B(_00312_),
    .C(_00314_),
    .Y(_00721_));
 sky130_fd_sc_hd__nand3_1 _06751_ (.A(_00720_),
    .B(_00721_),
    .C(_00330_),
    .Y(_00722_));
 sky130_fd_sc_hd__nand2_1 _06752_ (.A(_00713_),
    .B(_00722_),
    .Y(_00723_));
 sky130_fd_sc_hd__inv_4 _06753_ (.A(_00316_),
    .Y(_00724_));
 sky130_fd_sc_hd__nand2_1 _06754_ (.A(_00724_),
    .B(_00317_),
    .Y(_00725_));
 sky130_fd_sc_hd__inv_2 _06755_ (.A(_00317_),
    .Y(_00726_));
 sky130_fd_sc_hd__nand2_1 _06756_ (.A(_00726_),
    .B(_00316_),
    .Y(_00727_));
 sky130_fd_sc_hd__nand3_1 _06757_ (.A(_00725_),
    .B(_00727_),
    .C(_00319_),
    .Y(_00728_));
 sky130_fd_sc_hd__nand2_1 _06758_ (.A(_00724_),
    .B(_00726_),
    .Y(_00729_));
 sky130_fd_sc_hd__nand3_1 _06759_ (.A(_00729_),
    .B(_00320_),
    .C(_00318_),
    .Y(_00730_));
 sky130_fd_sc_hd__nand2_1 _06760_ (.A(_00728_),
    .B(_00730_),
    .Y(_00731_));
 sky130_fd_sc_hd__nand2_1 _06761_ (.A(_02544_),
    .B(_00751_),
    .Y(_00732_));
 sky130_fd_sc_hd__nand2_1 _06762_ (.A(_01147_),
    .B(_00795_),
    .Y(_00733_));
 sky130_fd_sc_hd__nand2_1 _06763_ (.A(_00732_),
    .B(_00733_),
    .Y(_00734_));
 sky130_fd_sc_hd__nand2_1 _06764_ (.A(_01873_),
    .B(_00861_),
    .Y(_00735_));
 sky130_fd_sc_hd__inv_2 _06765_ (.A(_00735_),
    .Y(_00736_));
 sky130_fd_sc_hd__nor2_1 _06766_ (.A(_00732_),
    .B(_00733_),
    .Y(_00737_));
 sky130_fd_sc_hd__a21oi_2 _06767_ (.A1(_00734_),
    .A2(_00736_),
    .B1(_00737_),
    .Y(_00738_));
 sky130_fd_sc_hd__nand2_1 _06768_ (.A(_00731_),
    .B(_00738_),
    .Y(_00739_));
 sky130_fd_sc_hd__inv_2 _06769_ (.A(_00635_),
    .Y(_00741_));
 sky130_fd_sc_hd__inv_2 _06770_ (.A(_00636_),
    .Y(_00742_));
 sky130_fd_sc_hd__nand2_1 _06771_ (.A(_00741_),
    .B(_00742_),
    .Y(_00743_));
 sky130_fd_sc_hd__nand2_1 _06772_ (.A(_00743_),
    .B(_00637_),
    .Y(_00744_));
 sky130_fd_sc_hd__nand2_1 _06773_ (.A(_00744_),
    .B(_00638_),
    .Y(_00745_));
 sky130_fd_sc_hd__nand3_1 _06774_ (.A(_00743_),
    .B(_00639_),
    .C(_00637_),
    .Y(_00746_));
 sky130_fd_sc_hd__nand2_1 _06775_ (.A(_00745_),
    .B(_00746_),
    .Y(_00747_));
 sky130_fd_sc_hd__inv_2 _06776_ (.A(_00747_),
    .Y(_00748_));
 sky130_fd_sc_hd__nor2_1 _06777_ (.A(_00738_),
    .B(_00731_),
    .Y(_00749_));
 sky130_fd_sc_hd__a21oi_1 _06778_ (.A1(_00739_),
    .A2(_00748_),
    .B1(_00749_),
    .Y(_00750_));
 sky130_fd_sc_hd__nand2_1 _06779_ (.A(_00723_),
    .B(_00750_),
    .Y(_00752_));
 sky130_fd_sc_hd__inv_2 _06780_ (.A(_00641_),
    .Y(_00753_));
 sky130_fd_sc_hd__nand2_1 _06781_ (.A(_00634_),
    .B(_00753_),
    .Y(_00754_));
 sky130_fd_sc_hd__nand3_1 _06782_ (.A(_00641_),
    .B(_00633_),
    .C(_00213_),
    .Y(_00755_));
 sky130_fd_sc_hd__nand2_1 _06783_ (.A(_00754_),
    .B(_00755_),
    .Y(_00756_));
 sky130_fd_sc_hd__nand2_1 _06784_ (.A(_00756_),
    .B(_00652_),
    .Y(_00757_));
 sky130_fd_sc_hd__nand3b_1 _06785_ (.A_N(_00652_),
    .B(_00754_),
    .C(_00755_),
    .Y(_00758_));
 sky130_fd_sc_hd__nand2_1 _06786_ (.A(_00757_),
    .B(_00758_),
    .Y(_00759_));
 sky130_fd_sc_hd__inv_2 _06787_ (.A(_00759_),
    .Y(_00760_));
 sky130_fd_sc_hd__nor2_1 _06788_ (.A(_00750_),
    .B(_00723_),
    .Y(_00761_));
 sky130_fd_sc_hd__a21oi_1 _06789_ (.A1(_00752_),
    .A2(_00760_),
    .B1(_00761_),
    .Y(_00763_));
 sky130_fd_sc_hd__nand2_1 _06790_ (.A(_00719_),
    .B(_00763_),
    .Y(_00764_));
 sky130_fd_sc_hd__nand3_1 _06791_ (.A(_00654_),
    .B(_00242_),
    .C(_00629_),
    .Y(_00765_));
 sky130_fd_sc_hd__inv_2 _06792_ (.A(_00654_),
    .Y(_00766_));
 sky130_fd_sc_hd__nand2_1 _06793_ (.A(_00766_),
    .B(_00630_),
    .Y(_00767_));
 sky130_fd_sc_hd__nand3b_1 _06794_ (.A_N(_00682_),
    .B(_00765_),
    .C(_00767_),
    .Y(_00768_));
 sky130_fd_sc_hd__nand2_1 _06795_ (.A(_00767_),
    .B(_00765_),
    .Y(_00769_));
 sky130_fd_sc_hd__nand2_1 _06796_ (.A(_00769_),
    .B(_00682_),
    .Y(_00770_));
 sky130_fd_sc_hd__nand2_1 _06797_ (.A(_00768_),
    .B(_00770_),
    .Y(_00771_));
 sky130_fd_sc_hd__inv_2 _06798_ (.A(_00771_),
    .Y(_00772_));
 sky130_fd_sc_hd__nor2_1 _06799_ (.A(_00763_),
    .B(_00719_),
    .Y(_00774_));
 sky130_fd_sc_hd__a21oi_1 _06800_ (.A1(_00764_),
    .A2(_00772_),
    .B1(_00774_),
    .Y(_00775_));
 sky130_fd_sc_hd__nand2_1 _06801_ (.A(_00709_),
    .B(_00775_),
    .Y(_00776_));
 sky130_fd_sc_hd__nor2_1 _06802_ (.A(_00775_),
    .B(_00709_),
    .Y(_00777_));
 sky130_fd_sc_hd__a21oi_1 _06803_ (.A1(_00705_),
    .A2(_00776_),
    .B1(_00777_),
    .Y(_00778_));
 sky130_fd_sc_hd__nand2_1 _06804_ (.A(_00626_),
    .B(_00778_),
    .Y(_00779_));
 sky130_fd_sc_hd__nand2_2 _06805_ (.A(_00703_),
    .B(_00687_),
    .Y(_00780_));
 sky130_fd_sc_hd__nor2_1 _06806_ (.A(_00778_),
    .B(_00626_),
    .Y(_00781_));
 sky130_fd_sc_hd__a21oi_2 _06807_ (.A1(_00779_),
    .A2(_00780_),
    .B1(_00781_),
    .Y(_00782_));
 sky130_fd_sc_hd__inv_2 _06808_ (.A(_00358_),
    .Y(_00783_));
 sky130_fd_sc_hd__nand2_1 _06809_ (.A(_00183_),
    .B(_00783_),
    .Y(_00785_));
 sky130_fd_sc_hd__nand3_1 _06810_ (.A(_00358_),
    .B(_00181_),
    .C(_00182_),
    .Y(_00786_));
 sky130_fd_sc_hd__nand2_1 _06811_ (.A(_00785_),
    .B(_00786_),
    .Y(_00787_));
 sky130_fd_sc_hd__nand2_1 _06812_ (.A(_00787_),
    .B(_00360_),
    .Y(_00788_));
 sky130_fd_sc_hd__nand3b_2 _06813_ (.A_N(_00360_),
    .B(_00785_),
    .C(_00786_),
    .Y(_00789_));
 sky130_fd_sc_hd__nand2_1 _06814_ (.A(_00788_),
    .B(_00789_),
    .Y(_00790_));
 sky130_fd_sc_hd__nor2_1 _06815_ (.A(_00782_),
    .B(_00790_),
    .Y(_00791_));
 sky130_fd_sc_hd__nand2_2 _06816_ (.A(_00366_),
    .B(_00362_),
    .Y(_00792_));
 sky130_fd_sc_hd__nand3_4 _06817_ (.A(_00614_),
    .B(_00791_),
    .C(_00792_),
    .Y(_00793_));
 sky130_fd_sc_hd__nand2_1 _06818_ (.A(_00616_),
    .B(_00793_),
    .Y(_00794_));
 sky130_fd_sc_hd__inv_2 _06819_ (.A(_00793_),
    .Y(_00796_));
 sky130_fd_sc_hd__nand3_2 _06820_ (.A(_00615_),
    .B(_00796_),
    .C(_00368_),
    .Y(_00797_));
 sky130_fd_sc_hd__nand2_1 _06821_ (.A(_00794_),
    .B(_00797_),
    .Y(_00798_));
 sky130_fd_sc_hd__nor2_1 _06822_ (.A(_00611_),
    .B(_00798_),
    .Y(_00799_));
 sky130_fd_sc_hd__nand3_1 _06823_ (.A(_00778_),
    .B(_00624_),
    .C(_00625_),
    .Y(_00800_));
 sky130_fd_sc_hd__a21o_1 _06824_ (.A1(_00705_),
    .A2(_00776_),
    .B1(_00777_),
    .X(_00801_));
 sky130_fd_sc_hd__nand2_1 _06825_ (.A(_00626_),
    .B(_00801_),
    .Y(_00802_));
 sky130_fd_sc_hd__nand2_1 _06826_ (.A(_00800_),
    .B(_00802_),
    .Y(_00803_));
 sky130_fd_sc_hd__nand2_2 _06827_ (.A(_00803_),
    .B(_00780_),
    .Y(_00804_));
 sky130_fd_sc_hd__inv_2 _06828_ (.A(_00780_),
    .Y(_00805_));
 sky130_fd_sc_hd__nand3_2 _06829_ (.A(_00800_),
    .B(_00802_),
    .C(_00805_),
    .Y(_00807_));
 sky130_fd_sc_hd__nand2_1 _06830_ (.A(_00804_),
    .B(_00807_),
    .Y(_00808_));
 sky130_fd_sc_hd__nand3_1 _06831_ (.A(_00775_),
    .B(_00620_),
    .C(_00708_),
    .Y(_00809_));
 sky130_fd_sc_hd__a21o_1 _06832_ (.A1(_00752_),
    .A2(_00760_),
    .B1(_00761_),
    .X(_00810_));
 sky130_fd_sc_hd__nand3_1 _06833_ (.A(_00810_),
    .B(_00717_),
    .C(_00718_),
    .Y(_00811_));
 sky130_fd_sc_hd__nand3_2 _06834_ (.A(_00811_),
    .B(_00764_),
    .C(_00772_),
    .Y(_00812_));
 sky130_fd_sc_hd__nand2_1 _06835_ (.A(_00812_),
    .B(_00811_),
    .Y(_00813_));
 sky130_fd_sc_hd__nand2_1 _06836_ (.A(_00813_),
    .B(_00709_),
    .Y(_00814_));
 sky130_fd_sc_hd__nand2_1 _06837_ (.A(_00809_),
    .B(_00814_),
    .Y(_00815_));
 sky130_fd_sc_hd__nand2_1 _06838_ (.A(_00815_),
    .B(_00705_),
    .Y(_00816_));
 sky130_fd_sc_hd__nand3_1 _06839_ (.A(_00809_),
    .B(_00814_),
    .C(_00704_),
    .Y(_00818_));
 sky130_fd_sc_hd__nand2_1 _06840_ (.A(_00816_),
    .B(_00818_),
    .Y(_00819_));
 sky130_fd_sc_hd__nand2_1 _06841_ (.A(_00719_),
    .B(_00810_),
    .Y(_00820_));
 sky130_fd_sc_hd__nand3_1 _06842_ (.A(_00763_),
    .B(_00717_),
    .C(_00718_),
    .Y(_00821_));
 sky130_fd_sc_hd__nand3_1 _06843_ (.A(_00820_),
    .B(_00821_),
    .C(_00771_),
    .Y(_00822_));
 sky130_fd_sc_hd__nand2_1 _06844_ (.A(_00812_),
    .B(_00822_),
    .Y(_00823_));
 sky130_fd_sc_hd__nand3_1 _06845_ (.A(_00750_),
    .B(_00713_),
    .C(_00722_),
    .Y(_00824_));
 sky130_fd_sc_hd__a21o_1 _06846_ (.A1(_00739_),
    .A2(_00748_),
    .B1(_00749_),
    .X(_00825_));
 sky130_fd_sc_hd__nand2_1 _06847_ (.A(_00825_),
    .B(_00723_),
    .Y(_00826_));
 sky130_fd_sc_hd__nand2_1 _06848_ (.A(_00824_),
    .B(_00826_),
    .Y(_00827_));
 sky130_fd_sc_hd__nand2_1 _06849_ (.A(_00827_),
    .B(_00760_),
    .Y(_00829_));
 sky130_fd_sc_hd__nand3_1 _06850_ (.A(_00824_),
    .B(_00826_),
    .C(_00759_),
    .Y(_00830_));
 sky130_fd_sc_hd__nand2_1 _06851_ (.A(_00829_),
    .B(_00830_),
    .Y(_00831_));
 sky130_fd_sc_hd__inv_2 _06852_ (.A(_00738_),
    .Y(_00832_));
 sky130_fd_sc_hd__nand2_1 _06853_ (.A(_00731_),
    .B(_00832_),
    .Y(_00833_));
 sky130_fd_sc_hd__nand3_1 _06854_ (.A(_00738_),
    .B(_00728_),
    .C(_00730_),
    .Y(_00834_));
 sky130_fd_sc_hd__nand2_1 _06855_ (.A(_00833_),
    .B(_00834_),
    .Y(_00835_));
 sky130_fd_sc_hd__nand2_1 _06856_ (.A(_00835_),
    .B(_00748_),
    .Y(_00836_));
 sky130_fd_sc_hd__nand3_1 _06857_ (.A(_00833_),
    .B(_00834_),
    .C(_00747_),
    .Y(_00837_));
 sky130_fd_sc_hd__nand2_1 _06858_ (.A(_00836_),
    .B(_00837_),
    .Y(_00838_));
 sky130_fd_sc_hd__inv_2 _06859_ (.A(_00732_),
    .Y(_00840_));
 sky130_fd_sc_hd__nand2_1 _06860_ (.A(_00840_),
    .B(_00733_),
    .Y(_00841_));
 sky130_fd_sc_hd__inv_2 _06861_ (.A(_00733_),
    .Y(_00842_));
 sky130_fd_sc_hd__nand2_1 _06862_ (.A(_00842_),
    .B(_00732_),
    .Y(_00843_));
 sky130_fd_sc_hd__nand3_1 _06863_ (.A(_00841_),
    .B(_00843_),
    .C(_00735_),
    .Y(_00844_));
 sky130_fd_sc_hd__nand2_1 _06864_ (.A(_00840_),
    .B(_00842_),
    .Y(_00845_));
 sky130_fd_sc_hd__nand3_1 _06865_ (.A(_00845_),
    .B(_00736_),
    .C(_00734_),
    .Y(_00846_));
 sky130_fd_sc_hd__nand2_1 _06866_ (.A(_00844_),
    .B(_00846_),
    .Y(_00847_));
 sky130_fd_sc_hd__nand2_2 _06867_ (.A(net4),
    .B(net44),
    .Y(_00848_));
 sky130_fd_sc_hd__nand2_1 _06868_ (.A(net5),
    .B(_00795_),
    .Y(_00849_));
 sky130_fd_sc_hd__nand2_1 _06869_ (.A(_00848_),
    .B(_00849_),
    .Y(_00851_));
 sky130_fd_sc_hd__nand2_1 _06870_ (.A(_02049_),
    .B(_00861_),
    .Y(_00852_));
 sky130_fd_sc_hd__inv_2 _06871_ (.A(_00852_),
    .Y(_00853_));
 sky130_fd_sc_hd__nor2_1 _06872_ (.A(_00848_),
    .B(_00849_),
    .Y(_00854_));
 sky130_fd_sc_hd__a21oi_2 _06873_ (.A1(_00851_),
    .A2(_00853_),
    .B1(_00854_),
    .Y(_00855_));
 sky130_fd_sc_hd__nand2_1 _06874_ (.A(_00847_),
    .B(_00855_),
    .Y(_00856_));
 sky130_fd_sc_hd__nand2_1 _06875_ (.A(_03160_),
    .B(_01048_),
    .Y(_00857_));
 sky130_fd_sc_hd__inv_2 _06876_ (.A(_00857_),
    .Y(_00858_));
 sky130_fd_sc_hd__nand2_1 _06877_ (.A(_02049_),
    .B(_01092_),
    .Y(_00859_));
 sky130_fd_sc_hd__inv_2 _06878_ (.A(_00859_),
    .Y(_00860_));
 sky130_fd_sc_hd__nand2_1 _06879_ (.A(_00858_),
    .B(_00860_),
    .Y(_00862_));
 sky130_fd_sc_hd__nand2_1 _06880_ (.A(_00857_),
    .B(_00859_),
    .Y(_00863_));
 sky130_fd_sc_hd__nand2_1 _06881_ (.A(_00862_),
    .B(_00863_),
    .Y(_00864_));
 sky130_fd_sc_hd__nand2_1 _06882_ (.A(_03094_),
    .B(_01158_),
    .Y(_00865_));
 sky130_fd_sc_hd__nand2_1 _06883_ (.A(_00864_),
    .B(_00865_),
    .Y(_00866_));
 sky130_fd_sc_hd__inv_2 _06884_ (.A(_00865_),
    .Y(_00867_));
 sky130_fd_sc_hd__nand3_1 _06885_ (.A(_00862_),
    .B(_00867_),
    .C(_00863_),
    .Y(_00868_));
 sky130_fd_sc_hd__nand2_1 _06886_ (.A(_00866_),
    .B(_00868_),
    .Y(_00869_));
 sky130_fd_sc_hd__inv_2 _06887_ (.A(_00869_),
    .Y(_00870_));
 sky130_fd_sc_hd__nor2_1 _06888_ (.A(_00855_),
    .B(_00847_),
    .Y(_00871_));
 sky130_fd_sc_hd__a21oi_1 _06889_ (.A1(_00856_),
    .A2(_00870_),
    .B1(_00871_),
    .Y(_00873_));
 sky130_fd_sc_hd__nand2_1 _06890_ (.A(_00838_),
    .B(_00873_),
    .Y(_00874_));
 sky130_fd_sc_hd__nand2_1 _06891_ (.A(_00644_),
    .B(_00645_),
    .Y(_00875_));
 sky130_fd_sc_hd__nand2_1 _06892_ (.A(_00646_),
    .B(_00643_),
    .Y(_00876_));
 sky130_fd_sc_hd__nand3_1 _06893_ (.A(_00875_),
    .B(_00876_),
    .C(_00648_),
    .Y(_00877_));
 sky130_fd_sc_hd__nand2_1 _06894_ (.A(_00877_),
    .B(_00651_),
    .Y(_00878_));
 sky130_fd_sc_hd__nor2_1 _06895_ (.A(_00857_),
    .B(_00859_),
    .Y(_00879_));
 sky130_fd_sc_hd__a21oi_2 _06896_ (.A1(_00863_),
    .A2(_00867_),
    .B1(_00879_),
    .Y(_00880_));
 sky130_fd_sc_hd__inv_2 _06897_ (.A(_00880_),
    .Y(_00881_));
 sky130_fd_sc_hd__nand2_1 _06898_ (.A(_00878_),
    .B(_00881_),
    .Y(_00882_));
 sky130_fd_sc_hd__nand3_1 _06899_ (.A(_00880_),
    .B(_00877_),
    .C(_00651_),
    .Y(_00884_));
 sky130_fd_sc_hd__nand2_1 _06900_ (.A(_00882_),
    .B(_00884_),
    .Y(_00885_));
 sky130_fd_sc_hd__nand2_1 _06901_ (.A(_04928_),
    .B(_00003_),
    .Y(_00886_));
 sky130_fd_sc_hd__nand2_1 _06902_ (.A(_05028_),
    .B(_00412_),
    .Y(_00887_));
 sky130_fd_sc_hd__inv_2 _06903_ (.A(_00887_),
    .Y(_00888_));
 sky130_fd_sc_hd__nand2_1 _06904_ (.A(_05031_),
    .B(_00204_),
    .Y(_00889_));
 sky130_fd_sc_hd__inv_2 _06905_ (.A(_00889_),
    .Y(_00890_));
 sky130_fd_sc_hd__nand2_1 _06906_ (.A(_00888_),
    .B(_00890_),
    .Y(_00891_));
 sky130_fd_sc_hd__nand2_1 _06907_ (.A(_00887_),
    .B(_00889_),
    .Y(_00892_));
 sky130_fd_sc_hd__nand3b_2 _06908_ (.A_N(_00886_),
    .B(_00891_),
    .C(_00892_),
    .Y(_00893_));
 sky130_fd_sc_hd__nand2_1 _06909_ (.A(_00893_),
    .B(_00891_),
    .Y(_00895_));
 sky130_fd_sc_hd__nand2_1 _06910_ (.A(_00885_),
    .B(_00895_),
    .Y(_00896_));
 sky130_fd_sc_hd__nand3b_1 _06911_ (.A_N(_00895_),
    .B(_00882_),
    .C(_00884_),
    .Y(_00897_));
 sky130_fd_sc_hd__nand2_1 _06912_ (.A(_00896_),
    .B(_00897_),
    .Y(_00898_));
 sky130_fd_sc_hd__inv_2 _06913_ (.A(_00898_),
    .Y(_00899_));
 sky130_fd_sc_hd__nor2_1 _06914_ (.A(_00873_),
    .B(_00838_),
    .Y(_00900_));
 sky130_fd_sc_hd__a21oi_2 _06915_ (.A1(_00874_),
    .A2(_00899_),
    .B1(_00900_),
    .Y(_00901_));
 sky130_fd_sc_hd__nand2_1 _06916_ (.A(_00831_),
    .B(_00901_),
    .Y(_00902_));
 sky130_fd_sc_hd__nand2_2 _06917_ (.A(_00254_),
    .B(_05029_),
    .Y(_00903_));
 sky130_fd_sc_hd__nand2_1 _06918_ (.A(_00656_),
    .B(_05032_),
    .Y(_00904_));
 sky130_fd_sc_hd__nand2_1 _06919_ (.A(_00903_),
    .B(_00904_),
    .Y(_00906_));
 sky130_fd_sc_hd__nand2_1 _06920_ (.A(_03215_),
    .B(_04819_),
    .Y(_00907_));
 sky130_fd_sc_hd__inv_2 _06921_ (.A(_00907_),
    .Y(_00908_));
 sky130_fd_sc_hd__nor2_1 _06922_ (.A(_00903_),
    .B(_00904_),
    .Y(_00909_));
 sky130_fd_sc_hd__a21oi_2 _06923_ (.A1(_00906_),
    .A2(_00908_),
    .B1(_00909_),
    .Y(_00910_));
 sky130_fd_sc_hd__inv_2 _06924_ (.A(_00658_),
    .Y(_00911_));
 sky130_fd_sc_hd__nand2_1 _06925_ (.A(_00911_),
    .B(_00657_),
    .Y(_00912_));
 sky130_fd_sc_hd__inv_2 _06926_ (.A(_00657_),
    .Y(_00913_));
 sky130_fd_sc_hd__nand2_1 _06927_ (.A(_00913_),
    .B(_00658_),
    .Y(_00914_));
 sky130_fd_sc_hd__nand3_1 _06928_ (.A(_00912_),
    .B(_00914_),
    .C(_00660_),
    .Y(_00915_));
 sky130_fd_sc_hd__nand2_1 _06929_ (.A(_00913_),
    .B(_00911_),
    .Y(_00917_));
 sky130_fd_sc_hd__nand3_1 _06930_ (.A(_00917_),
    .B(_00661_),
    .C(_00659_),
    .Y(_00918_));
 sky130_fd_sc_hd__nand2_1 _06931_ (.A(_00915_),
    .B(_00918_),
    .Y(_00919_));
 sky130_fd_sc_hd__inv_2 _06932_ (.A(_00910_),
    .Y(_00920_));
 sky130_fd_sc_hd__nand2_1 _06933_ (.A(_00919_),
    .B(_00920_),
    .Y(_00921_));
 sky130_fd_sc_hd__nand3_1 _06934_ (.A(_00910_),
    .B(_00915_),
    .C(_00918_),
    .Y(_00922_));
 sky130_fd_sc_hd__nand2_1 _06935_ (.A(_00921_),
    .B(_00922_),
    .Y(_00923_));
 sky130_fd_sc_hd__nand2_1 _06936_ (.A(_00695_),
    .B(_00696_),
    .Y(_00924_));
 sky130_fd_sc_hd__nand2_1 _06937_ (.A(_00924_),
    .B(_00692_),
    .Y(_00925_));
 sky130_fd_sc_hd__nand2_1 _06938_ (.A(_00925_),
    .B(_00697_),
    .Y(_00926_));
 sky130_fd_sc_hd__inv_2 _06939_ (.A(_00926_),
    .Y(_00928_));
 sky130_fd_sc_hd__nand2_1 _06940_ (.A(_00923_),
    .B(_00928_),
    .Y(_00929_));
 sky130_fd_sc_hd__o21ai_1 _06941_ (.A1(_00910_),
    .A2(_00919_),
    .B1(_00929_),
    .Y(_00930_));
 sky130_fd_sc_hd__nand2_1 _06942_ (.A(_00878_),
    .B(_00880_),
    .Y(_00931_));
 sky130_fd_sc_hd__nor2_1 _06943_ (.A(_00880_),
    .B(_00878_),
    .Y(_00932_));
 sky130_fd_sc_hd__a21oi_2 _06944_ (.A1(_00931_),
    .A2(_00895_),
    .B1(_00932_),
    .Y(_00933_));
 sky130_fd_sc_hd__inv_2 _06945_ (.A(_00933_),
    .Y(_00934_));
 sky130_fd_sc_hd__nand3_1 _06946_ (.A(_00673_),
    .B(_00674_),
    .C(_00679_),
    .Y(_00935_));
 sky130_fd_sc_hd__nand2_1 _06947_ (.A(_00681_),
    .B(_00935_),
    .Y(_00936_));
 sky130_fd_sc_hd__nand2_1 _06948_ (.A(_00934_),
    .B(_00936_),
    .Y(_00937_));
 sky130_fd_sc_hd__nand3_1 _06949_ (.A(_00933_),
    .B(_00681_),
    .C(_00935_),
    .Y(_00939_));
 sky130_fd_sc_hd__nand3b_1 _06950_ (.A_N(_00930_),
    .B(_00937_),
    .C(_00939_),
    .Y(_00940_));
 sky130_fd_sc_hd__nand2_1 _06951_ (.A(_00937_),
    .B(_00939_),
    .Y(_00941_));
 sky130_fd_sc_hd__nand2_1 _06952_ (.A(_00941_),
    .B(_00930_),
    .Y(_00942_));
 sky130_fd_sc_hd__nand2_1 _06953_ (.A(_00940_),
    .B(_00942_),
    .Y(_00943_));
 sky130_fd_sc_hd__inv_2 _06954_ (.A(_00943_),
    .Y(_00944_));
 sky130_fd_sc_hd__nor2_1 _06955_ (.A(_00901_),
    .B(_00831_),
    .Y(_00945_));
 sky130_fd_sc_hd__a21oi_2 _06956_ (.A1(_00902_),
    .A2(_00944_),
    .B1(_00945_),
    .Y(_00946_));
 sky130_fd_sc_hd__nand2_1 _06957_ (.A(_00823_),
    .B(_00946_),
    .Y(_00947_));
 sky130_fd_sc_hd__nand2_1 _06958_ (.A(_00936_),
    .B(_00933_),
    .Y(_00948_));
 sky130_fd_sc_hd__nor2_1 _06959_ (.A(_00933_),
    .B(_00936_),
    .Y(_00950_));
 sky130_fd_sc_hd__a21oi_1 _06960_ (.A1(_00948_),
    .A2(_00930_),
    .B1(_00950_),
    .Y(_00951_));
 sky130_fd_sc_hd__inv_2 _06961_ (.A(_00951_),
    .Y(_00952_));
 sky130_fd_sc_hd__nand2_1 _06962_ (.A(_00689_),
    .B(_00274_),
    .Y(_00953_));
 sky130_fd_sc_hd__inv_2 _06963_ (.A(_00699_),
    .Y(_00954_));
 sky130_fd_sc_hd__nand2_1 _06964_ (.A(_00953_),
    .B(_00954_),
    .Y(_00955_));
 sky130_fd_sc_hd__nand2_1 _06965_ (.A(_00955_),
    .B(_00700_),
    .Y(_00956_));
 sky130_fd_sc_hd__inv_2 _06966_ (.A(_00956_),
    .Y(_00957_));
 sky130_fd_sc_hd__nand2_1 _06967_ (.A(_00952_),
    .B(_00957_),
    .Y(_00958_));
 sky130_fd_sc_hd__nand2_1 _06968_ (.A(_00951_),
    .B(_00956_),
    .Y(_00959_));
 sky130_fd_sc_hd__nand2_1 _06969_ (.A(_00958_),
    .B(_00959_),
    .Y(_00961_));
 sky130_fd_sc_hd__nand2_1 _06970_ (.A(_04812_),
    .B(_04992_),
    .Y(_00962_));
 sky130_fd_sc_hd__nand2_1 _06971_ (.A(_03809_),
    .B(_04895_),
    .Y(_00963_));
 sky130_fd_sc_hd__nand2_1 _06972_ (.A(_04962_),
    .B(_04911_),
    .Y(_00964_));
 sky130_fd_sc_hd__inv_2 _06973_ (.A(_00964_),
    .Y(_00965_));
 sky130_fd_sc_hd__nand2_1 _06974_ (.A(_04964_),
    .B(_04828_),
    .Y(_00966_));
 sky130_fd_sc_hd__inv_2 _06975_ (.A(_00966_),
    .Y(_00967_));
 sky130_fd_sc_hd__nand2_1 _06976_ (.A(_00965_),
    .B(_00967_),
    .Y(_00968_));
 sky130_fd_sc_hd__nand2_1 _06977_ (.A(_00964_),
    .B(_00966_),
    .Y(_00969_));
 sky130_fd_sc_hd__nand3b_1 _06978_ (.A_N(_00963_),
    .B(_00968_),
    .C(_00969_),
    .Y(_00970_));
 sky130_fd_sc_hd__and2_1 _06979_ (.A(_00970_),
    .B(_00968_),
    .X(_00972_));
 sky130_fd_sc_hd__nor2_1 _06980_ (.A(_00962_),
    .B(_00972_),
    .Y(_00973_));
 sky130_fd_sc_hd__inv_2 _06981_ (.A(_00973_),
    .Y(_00974_));
 sky130_fd_sc_hd__nand2_1 _06982_ (.A(_00698_),
    .B(_00691_),
    .Y(_00975_));
 sky130_fd_sc_hd__nand2_1 _06983_ (.A(_00954_),
    .B(_00975_),
    .Y(_00976_));
 sky130_fd_sc_hd__or2_1 _06984_ (.A(_00974_),
    .B(_00976_),
    .X(_00977_));
 sky130_fd_sc_hd__nand2_1 _06985_ (.A(_00961_),
    .B(_00977_),
    .Y(_00978_));
 sky130_fd_sc_hd__nand3b_1 _06986_ (.A_N(_00977_),
    .B(_00958_),
    .C(_00959_),
    .Y(_00979_));
 sky130_fd_sc_hd__nand2_1 _06987_ (.A(_00978_),
    .B(_00979_),
    .Y(_00980_));
 sky130_fd_sc_hd__inv_2 _06988_ (.A(_00980_),
    .Y(_00981_));
 sky130_fd_sc_hd__nor2_1 _06989_ (.A(_00946_),
    .B(_00823_),
    .Y(_00983_));
 sky130_fd_sc_hd__a21oi_2 _06990_ (.A1(_00947_),
    .A2(_00981_),
    .B1(_00983_),
    .Y(_00984_));
 sky130_fd_sc_hd__nand2_1 _06991_ (.A(_00819_),
    .B(_00984_),
    .Y(_00985_));
 sky130_fd_sc_hd__nand2_2 _06992_ (.A(_00979_),
    .B(_00958_),
    .Y(_00986_));
 sky130_fd_sc_hd__nor2_1 _06993_ (.A(_00984_),
    .B(_00819_),
    .Y(_00987_));
 sky130_fd_sc_hd__a21oi_2 _06994_ (.A1(_00985_),
    .A2(_00986_),
    .B1(_00987_),
    .Y(_00988_));
 sky130_fd_sc_hd__inv_2 _06995_ (.A(_00988_),
    .Y(_00989_));
 sky130_fd_sc_hd__nand2_1 _06996_ (.A(_00808_),
    .B(_00989_),
    .Y(_00990_));
 sky130_fd_sc_hd__nand3_1 _06997_ (.A(_00988_),
    .B(_00804_),
    .C(_00807_),
    .Y(_00991_));
 sky130_fd_sc_hd__nand2_1 _06998_ (.A(_00990_),
    .B(_00991_),
    .Y(_00992_));
 sky130_fd_sc_hd__nand3_1 _06999_ (.A(_00946_),
    .B(_00812_),
    .C(_00822_),
    .Y(_00994_));
 sky130_fd_sc_hd__inv_2 _07000_ (.A(_00946_),
    .Y(_00995_));
 sky130_fd_sc_hd__nand2_1 _07001_ (.A(_00995_),
    .B(_00823_),
    .Y(_00996_));
 sky130_fd_sc_hd__nand2_1 _07002_ (.A(_00994_),
    .B(_00996_),
    .Y(_00997_));
 sky130_fd_sc_hd__nand2_1 _07003_ (.A(_00997_),
    .B(_00981_),
    .Y(_00998_));
 sky130_fd_sc_hd__nand3_1 _07004_ (.A(_00994_),
    .B(_00996_),
    .C(_00980_),
    .Y(_00999_));
 sky130_fd_sc_hd__nand2_1 _07005_ (.A(_00998_),
    .B(_00999_),
    .Y(_01000_));
 sky130_fd_sc_hd__inv_2 _07006_ (.A(_00901_),
    .Y(_01001_));
 sky130_fd_sc_hd__nand2_1 _07007_ (.A(_00831_),
    .B(_01001_),
    .Y(_01002_));
 sky130_fd_sc_hd__nand3_1 _07008_ (.A(_00901_),
    .B(_00829_),
    .C(_00830_),
    .Y(_01003_));
 sky130_fd_sc_hd__nand2_1 _07009_ (.A(_01002_),
    .B(_01003_),
    .Y(_01005_));
 sky130_fd_sc_hd__nand2_1 _07010_ (.A(_01005_),
    .B(_00944_),
    .Y(_01006_));
 sky130_fd_sc_hd__nand3_1 _07011_ (.A(_01002_),
    .B(_01003_),
    .C(_00943_),
    .Y(_01007_));
 sky130_fd_sc_hd__nand2_1 _07012_ (.A(_01006_),
    .B(_01007_),
    .Y(_01008_));
 sky130_fd_sc_hd__nand3_1 _07013_ (.A(_00873_),
    .B(_00836_),
    .C(_00837_),
    .Y(_01009_));
 sky130_fd_sc_hd__inv_2 _07014_ (.A(_00855_),
    .Y(_01010_));
 sky130_fd_sc_hd__nand3_1 _07015_ (.A(_01010_),
    .B(_00846_),
    .C(_00844_),
    .Y(_01011_));
 sky130_fd_sc_hd__nand3_1 _07016_ (.A(_01011_),
    .B(_00856_),
    .C(_00870_),
    .Y(_01012_));
 sky130_fd_sc_hd__nand2_1 _07017_ (.A(_01012_),
    .B(_01011_),
    .Y(_01013_));
 sky130_fd_sc_hd__nand2_1 _07018_ (.A(_00838_),
    .B(_01013_),
    .Y(_01014_));
 sky130_fd_sc_hd__nand2_1 _07019_ (.A(_01009_),
    .B(_01014_),
    .Y(_01016_));
 sky130_fd_sc_hd__nand2_1 _07020_ (.A(_01016_),
    .B(_00899_),
    .Y(_01017_));
 sky130_fd_sc_hd__nand3_1 _07021_ (.A(_01009_),
    .B(_01014_),
    .C(_00898_),
    .Y(_01018_));
 sky130_fd_sc_hd__nand2_1 _07022_ (.A(_01017_),
    .B(_01018_),
    .Y(_01019_));
 sky130_fd_sc_hd__nand2_1 _07023_ (.A(_00847_),
    .B(_01010_),
    .Y(_01020_));
 sky130_fd_sc_hd__nand3_1 _07024_ (.A(_00855_),
    .B(_00844_),
    .C(_00846_),
    .Y(_01021_));
 sky130_fd_sc_hd__nand3_1 _07025_ (.A(_01020_),
    .B(_01021_),
    .C(_00869_),
    .Y(_01022_));
 sky130_fd_sc_hd__nand2_1 _07026_ (.A(_01012_),
    .B(_01022_),
    .Y(_01023_));
 sky130_fd_sc_hd__inv_2 _07027_ (.A(_00848_),
    .Y(_01024_));
 sky130_fd_sc_hd__nand2_1 _07028_ (.A(_01024_),
    .B(_00849_),
    .Y(_01025_));
 sky130_fd_sc_hd__inv_2 _07029_ (.A(_00849_),
    .Y(_01027_));
 sky130_fd_sc_hd__nand2_1 _07030_ (.A(_01027_),
    .B(_00848_),
    .Y(_01028_));
 sky130_fd_sc_hd__nand3_1 _07031_ (.A(_01025_),
    .B(_01028_),
    .C(_00852_),
    .Y(_01029_));
 sky130_fd_sc_hd__nand2_1 _07032_ (.A(_01024_),
    .B(_01027_),
    .Y(_01030_));
 sky130_fd_sc_hd__nand3_1 _07033_ (.A(_01030_),
    .B(_00853_),
    .C(_00851_),
    .Y(_01031_));
 sky130_fd_sc_hd__nand2_1 _07034_ (.A(_01029_),
    .B(_01031_),
    .Y(_01032_));
 sky130_fd_sc_hd__nand2_1 _07035_ (.A(_02049_),
    .B(_00751_),
    .Y(_01033_));
 sky130_fd_sc_hd__nand2_1 _07036_ (.A(_01873_),
    .B(_00795_),
    .Y(_01034_));
 sky130_fd_sc_hd__nand2_1 _07037_ (.A(_01033_),
    .B(_01034_),
    .Y(_01035_));
 sky130_fd_sc_hd__nand2_1 _07038_ (.A(_03160_),
    .B(_00861_),
    .Y(_01036_));
 sky130_fd_sc_hd__inv_2 _07039_ (.A(_01036_),
    .Y(_01038_));
 sky130_fd_sc_hd__nor2_1 _07040_ (.A(_01033_),
    .B(_01034_),
    .Y(_01039_));
 sky130_fd_sc_hd__a21oi_1 _07041_ (.A1(_01035_),
    .A2(_01038_),
    .B1(_01039_),
    .Y(_01040_));
 sky130_fd_sc_hd__nand2_1 _07042_ (.A(_01032_),
    .B(_01040_),
    .Y(_01041_));
 sky130_fd_sc_hd__nand2_2 _07043_ (.A(_03094_),
    .B(_01048_),
    .Y(_01042_));
 sky130_fd_sc_hd__inv_2 _07044_ (.A(_01042_),
    .Y(_01043_));
 sky130_fd_sc_hd__nand2_1 _07045_ (.A(_02753_),
    .B(_01092_),
    .Y(_01044_));
 sky130_fd_sc_hd__nand2_1 _07046_ (.A(_01043_),
    .B(_01044_),
    .Y(_01045_));
 sky130_fd_sc_hd__inv_2 _07047_ (.A(_01044_),
    .Y(_01046_));
 sky130_fd_sc_hd__nand2_1 _07048_ (.A(_01046_),
    .B(_01042_),
    .Y(_01047_));
 sky130_fd_sc_hd__nand2_1 _07049_ (.A(_03226_),
    .B(_01158_),
    .Y(_01049_));
 sky130_fd_sc_hd__nand3_1 _07050_ (.A(_01045_),
    .B(_01047_),
    .C(_01049_),
    .Y(_01050_));
 sky130_fd_sc_hd__nand2_1 _07051_ (.A(_01043_),
    .B(_01046_),
    .Y(_01051_));
 sky130_fd_sc_hd__inv_2 _07052_ (.A(_01049_),
    .Y(_01052_));
 sky130_fd_sc_hd__nand2_1 _07053_ (.A(_01042_),
    .B(_01044_),
    .Y(_01053_));
 sky130_fd_sc_hd__nand3_1 _07054_ (.A(_01051_),
    .B(_01052_),
    .C(_01053_),
    .Y(_01054_));
 sky130_fd_sc_hd__nand2_1 _07055_ (.A(_01050_),
    .B(_01054_),
    .Y(_01055_));
 sky130_fd_sc_hd__inv_2 _07056_ (.A(_01055_),
    .Y(_01056_));
 sky130_fd_sc_hd__nor2_1 _07057_ (.A(_01040_),
    .B(_01032_),
    .Y(_01057_));
 sky130_fd_sc_hd__a21oi_1 _07058_ (.A1(_01041_),
    .A2(_01056_),
    .B1(_01057_),
    .Y(_01058_));
 sky130_fd_sc_hd__nand2_1 _07059_ (.A(_01023_),
    .B(_01058_),
    .Y(_01060_));
 sky130_fd_sc_hd__nor2_1 _07060_ (.A(_01042_),
    .B(_01044_),
    .Y(_01061_));
 sky130_fd_sc_hd__a21oi_2 _07061_ (.A1(_01053_),
    .A2(_01052_),
    .B1(_01061_),
    .Y(_01062_));
 sky130_fd_sc_hd__inv_2 _07062_ (.A(_01062_),
    .Y(_01063_));
 sky130_fd_sc_hd__nand2_1 _07063_ (.A(_00891_),
    .B(_00892_),
    .Y(_01064_));
 sky130_fd_sc_hd__nand2_1 _07064_ (.A(_01064_),
    .B(_00886_),
    .Y(_01065_));
 sky130_fd_sc_hd__nand3_1 _07065_ (.A(_01063_),
    .B(_00893_),
    .C(_01065_),
    .Y(_01066_));
 sky130_fd_sc_hd__nand2_1 _07066_ (.A(_01065_),
    .B(_00893_),
    .Y(_01067_));
 sky130_fd_sc_hd__nand2_1 _07067_ (.A(_01067_),
    .B(_01062_),
    .Y(_01068_));
 sky130_fd_sc_hd__nand2_1 _07068_ (.A(_04928_),
    .B(_01774_),
    .Y(_01069_));
 sky130_fd_sc_hd__inv_2 _07069_ (.A(_01069_),
    .Y(_01071_));
 sky130_fd_sc_hd__nand2_1 _07070_ (.A(_03314_),
    .B(_01807_),
    .Y(_01072_));
 sky130_fd_sc_hd__inv_2 _07071_ (.A(_01072_),
    .Y(_01073_));
 sky130_fd_sc_hd__nand2_1 _07072_ (.A(_01071_),
    .B(_01073_),
    .Y(_01074_));
 sky130_fd_sc_hd__nand2_1 _07073_ (.A(_00656_),
    .B(_01884_),
    .Y(_01075_));
 sky130_fd_sc_hd__inv_2 _07074_ (.A(_01075_),
    .Y(_01076_));
 sky130_fd_sc_hd__nand2_1 _07075_ (.A(_01069_),
    .B(_01072_),
    .Y(_01077_));
 sky130_fd_sc_hd__nand3_1 _07076_ (.A(_01074_),
    .B(_01076_),
    .C(_01077_),
    .Y(_01078_));
 sky130_fd_sc_hd__nand2_1 _07077_ (.A(_01078_),
    .B(_01074_),
    .Y(_01079_));
 sky130_fd_sc_hd__nand3_1 _07078_ (.A(_01066_),
    .B(_01068_),
    .C(_01079_),
    .Y(_01080_));
 sky130_fd_sc_hd__nand2_1 _07079_ (.A(_01067_),
    .B(_01063_),
    .Y(_01082_));
 sky130_fd_sc_hd__nand3_1 _07080_ (.A(_01065_),
    .B(_00893_),
    .C(_01062_),
    .Y(_01083_));
 sky130_fd_sc_hd__inv_2 _07081_ (.A(_01079_),
    .Y(_01084_));
 sky130_fd_sc_hd__nand3_1 _07082_ (.A(_01082_),
    .B(_01083_),
    .C(_01084_),
    .Y(_01085_));
 sky130_fd_sc_hd__nand2_1 _07083_ (.A(_01080_),
    .B(_01085_),
    .Y(_01086_));
 sky130_fd_sc_hd__inv_2 _07084_ (.A(_01086_),
    .Y(_01087_));
 sky130_fd_sc_hd__nor2_1 _07085_ (.A(_01058_),
    .B(_01023_),
    .Y(_01088_));
 sky130_fd_sc_hd__a21oi_1 _07086_ (.A1(_01060_),
    .A2(_01087_),
    .B1(_01088_),
    .Y(_01089_));
 sky130_fd_sc_hd__nand2_1 _07087_ (.A(_01019_),
    .B(_01089_),
    .Y(_01090_));
 sky130_fd_sc_hd__nor2_1 _07088_ (.A(_01062_),
    .B(_01067_),
    .Y(_01091_));
 sky130_fd_sc_hd__a21oi_1 _07089_ (.A1(_01068_),
    .A2(_01079_),
    .B1(_01091_),
    .Y(_01093_));
 sky130_fd_sc_hd__nand3_1 _07090_ (.A(_00921_),
    .B(_00926_),
    .C(_00922_),
    .Y(_01094_));
 sky130_fd_sc_hd__nand3_1 _07091_ (.A(_01093_),
    .B(_00929_),
    .C(_01094_),
    .Y(_01095_));
 sky130_fd_sc_hd__nand2_1 _07092_ (.A(_01080_),
    .B(_01066_),
    .Y(_01096_));
 sky130_fd_sc_hd__nand2_1 _07093_ (.A(_00929_),
    .B(_01094_),
    .Y(_01097_));
 sky130_fd_sc_hd__nand2_1 _07094_ (.A(_01096_),
    .B(_01097_),
    .Y(_01098_));
 sky130_fd_sc_hd__nand2_1 _07095_ (.A(_01095_),
    .B(_01098_),
    .Y(_01099_));
 sky130_fd_sc_hd__nand2_1 _07096_ (.A(_00968_),
    .B(_00969_),
    .Y(_01100_));
 sky130_fd_sc_hd__nand2_1 _07097_ (.A(_01100_),
    .B(_00963_),
    .Y(_01101_));
 sky130_fd_sc_hd__nand2_1 _07098_ (.A(_01101_),
    .B(_00970_),
    .Y(_01102_));
 sky130_fd_sc_hd__nand2_1 _07099_ (.A(_00522_),
    .B(_05029_),
    .Y(_01104_));
 sky130_fd_sc_hd__nand2_1 _07100_ (.A(_00254_),
    .B(_05032_),
    .Y(_01105_));
 sky130_fd_sc_hd__nand2_1 _07101_ (.A(_01104_),
    .B(_01105_),
    .Y(_01106_));
 sky130_fd_sc_hd__nand2_1 _07102_ (.A(_03215_),
    .B(_04828_),
    .Y(_01107_));
 sky130_fd_sc_hd__inv_2 _07103_ (.A(_01107_),
    .Y(_01108_));
 sky130_fd_sc_hd__nor2_1 _07104_ (.A(_01104_),
    .B(_01105_),
    .Y(_01109_));
 sky130_fd_sc_hd__a21o_1 _07105_ (.A1(_01106_),
    .A2(_01108_),
    .B1(_01109_),
    .X(_01110_));
 sky130_fd_sc_hd__inv_2 _07106_ (.A(_00903_),
    .Y(_01111_));
 sky130_fd_sc_hd__inv_2 _07107_ (.A(_00904_),
    .Y(_01112_));
 sky130_fd_sc_hd__nand2_1 _07108_ (.A(_01111_),
    .B(_01112_),
    .Y(_01113_));
 sky130_fd_sc_hd__nand3_1 _07109_ (.A(_01113_),
    .B(_00908_),
    .C(_00906_),
    .Y(_01115_));
 sky130_fd_sc_hd__nand2_1 _07110_ (.A(_01111_),
    .B(_00904_),
    .Y(_01116_));
 sky130_fd_sc_hd__nand2_1 _07111_ (.A(_01112_),
    .B(_00903_),
    .Y(_01117_));
 sky130_fd_sc_hd__nand3_1 _07112_ (.A(_01116_),
    .B(_01117_),
    .C(_00907_),
    .Y(_01118_));
 sky130_fd_sc_hd__nand3_1 _07113_ (.A(_01110_),
    .B(_01115_),
    .C(_01118_),
    .Y(_01119_));
 sky130_fd_sc_hd__nand2_1 _07114_ (.A(_01118_),
    .B(_01115_),
    .Y(_01120_));
 sky130_fd_sc_hd__a21oi_1 _07115_ (.A1(_01106_),
    .A2(_01108_),
    .B1(_01109_),
    .Y(_01121_));
 sky130_fd_sc_hd__nand2_1 _07116_ (.A(_01120_),
    .B(_01121_),
    .Y(_01122_));
 sky130_fd_sc_hd__nand3b_1 _07117_ (.A_N(_01102_),
    .B(_01119_),
    .C(_01122_),
    .Y(_01123_));
 sky130_fd_sc_hd__nand2_1 _07118_ (.A(_01123_),
    .B(_01119_),
    .Y(_01124_));
 sky130_fd_sc_hd__nand2_1 _07119_ (.A(_01099_),
    .B(_01124_),
    .Y(_01126_));
 sky130_fd_sc_hd__nand3b_1 _07120_ (.A_N(_01124_),
    .B(_01095_),
    .C(_01098_),
    .Y(_01127_));
 sky130_fd_sc_hd__nand2_1 _07121_ (.A(_01126_),
    .B(_01127_),
    .Y(_01128_));
 sky130_fd_sc_hd__inv_2 _07122_ (.A(_01128_),
    .Y(_01129_));
 sky130_fd_sc_hd__nor2_1 _07123_ (.A(_01089_),
    .B(_01019_),
    .Y(_01130_));
 sky130_fd_sc_hd__a21oi_1 _07124_ (.A1(_01090_),
    .A2(_01129_),
    .B1(_01130_),
    .Y(_01131_));
 sky130_fd_sc_hd__nand2_1 _07125_ (.A(_01008_),
    .B(_01131_),
    .Y(_01132_));
 sky130_fd_sc_hd__nand2_1 _07126_ (.A(_00976_),
    .B(_00974_),
    .Y(_01133_));
 sky130_fd_sc_hd__nand2_2 _07127_ (.A(_00977_),
    .B(_01133_),
    .Y(_01134_));
 sky130_fd_sc_hd__o21a_1 _07128_ (.A1(_01097_),
    .A2(_01093_),
    .B1(_01126_),
    .X(_01135_));
 sky130_fd_sc_hd__xor2_2 _07129_ (.A(_01134_),
    .B(_01135_),
    .X(_01137_));
 sky130_fd_sc_hd__nor2_1 _07130_ (.A(_01131_),
    .B(_01008_),
    .Y(_01138_));
 sky130_fd_sc_hd__a21oi_2 _07131_ (.A1(_01132_),
    .A2(_01137_),
    .B1(_01138_),
    .Y(_01139_));
 sky130_fd_sc_hd__nand2_1 _07132_ (.A(_01000_),
    .B(_01139_),
    .Y(_01140_));
 sky130_fd_sc_hd__nor2_2 _07133_ (.A(_01134_),
    .B(_01135_),
    .Y(_01141_));
 sky130_fd_sc_hd__nor2_1 _07134_ (.A(_01139_),
    .B(_01000_),
    .Y(_01142_));
 sky130_fd_sc_hd__a21oi_1 _07135_ (.A1(_01140_),
    .A2(_01141_),
    .B1(_01142_),
    .Y(_01143_));
 sky130_fd_sc_hd__inv_2 _07136_ (.A(_00984_),
    .Y(_01144_));
 sky130_fd_sc_hd__nand2_1 _07137_ (.A(_00819_),
    .B(_01144_),
    .Y(_01145_));
 sky130_fd_sc_hd__nand3_1 _07138_ (.A(_00984_),
    .B(_00816_),
    .C(_00818_),
    .Y(_01146_));
 sky130_fd_sc_hd__nand2_1 _07139_ (.A(_01145_),
    .B(_01146_),
    .Y(_01148_));
 sky130_fd_sc_hd__nand2_1 _07140_ (.A(_01148_),
    .B(_00986_),
    .Y(_01149_));
 sky130_fd_sc_hd__inv_2 _07141_ (.A(_00986_),
    .Y(_01150_));
 sky130_fd_sc_hd__nand3_1 _07142_ (.A(_01145_),
    .B(_01146_),
    .C(_01150_),
    .Y(_01151_));
 sky130_fd_sc_hd__nand2_1 _07143_ (.A(_01149_),
    .B(_01151_),
    .Y(_01152_));
 sky130_fd_sc_hd__nor2_1 _07144_ (.A(_01143_),
    .B(_01152_),
    .Y(_01153_));
 sky130_fd_sc_hd__nand2_1 _07145_ (.A(_00992_),
    .B(_01153_),
    .Y(_01154_));
 sky130_fd_sc_hd__nand3_1 _07146_ (.A(_00989_),
    .B(_00804_),
    .C(_00807_),
    .Y(_01155_));
 sky130_fd_sc_hd__nand3b_4 _07147_ (.A_N(_00782_),
    .B(_00788_),
    .C(_00789_),
    .Y(_01156_));
 sky130_fd_sc_hd__nand2_2 _07148_ (.A(_00790_),
    .B(_00782_),
    .Y(_01157_));
 sky130_fd_sc_hd__nand3b_2 _07149_ (.A_N(_01155_),
    .B(_01156_),
    .C(_01157_),
    .Y(_01159_));
 sky130_fd_sc_hd__nand2_1 _07150_ (.A(_01156_),
    .B(_01157_),
    .Y(_01160_));
 sky130_fd_sc_hd__nand2_1 _07151_ (.A(_01160_),
    .B(_01155_),
    .Y(_01161_));
 sky130_fd_sc_hd__nand3b_2 _07152_ (.A_N(_01154_),
    .B(_01159_),
    .C(_01161_),
    .Y(_01162_));
 sky130_fd_sc_hd__nand2_1 _07153_ (.A(_00614_),
    .B(_00792_),
    .Y(_01163_));
 sky130_fd_sc_hd__nand2_2 _07154_ (.A(_01163_),
    .B(_01156_),
    .Y(_01164_));
 sky130_fd_sc_hd__inv_2 _07155_ (.A(_01159_),
    .Y(_01165_));
 sky130_fd_sc_hd__a21oi_1 _07156_ (.A1(_01164_),
    .A2(_00793_),
    .B1(_01165_),
    .Y(_01166_));
 sky130_fd_sc_hd__nand3_1 _07157_ (.A(_01165_),
    .B(_00793_),
    .C(_01164_),
    .Y(_01167_));
 sky130_fd_sc_hd__o21ai_1 _07158_ (.A1(_01162_),
    .A2(_01166_),
    .B1(_01167_),
    .Y(_01168_));
 sky130_fd_sc_hd__nand2_1 _07159_ (.A(_00799_),
    .B(_01168_),
    .Y(_01170_));
 sky130_fd_sc_hd__inv_2 _07160_ (.A(_00797_),
    .Y(_01171_));
 sky130_fd_sc_hd__a21boi_1 _07161_ (.A1(_01171_),
    .A2(_00610_),
    .B1_N(_00604_),
    .Y(_01172_));
 sky130_fd_sc_hd__nand2_1 _07162_ (.A(_01170_),
    .B(_01172_),
    .Y(_01173_));
 sky130_fd_sc_hd__nand2_1 _07163_ (.A(_03226_),
    .B(_01048_),
    .Y(_01174_));
 sky130_fd_sc_hd__nand2_1 _07164_ (.A(_03094_),
    .B(_01092_),
    .Y(_01175_));
 sky130_fd_sc_hd__nor2_1 _07165_ (.A(_01174_),
    .B(_01175_),
    .Y(_01176_));
 sky130_fd_sc_hd__nand2_1 _07166_ (.A(_05028_),
    .B(_01158_),
    .Y(_01177_));
 sky130_fd_sc_hd__inv_2 _07167_ (.A(_01177_),
    .Y(_01178_));
 sky130_fd_sc_hd__nand2_1 _07168_ (.A(_01174_),
    .B(_01175_),
    .Y(_01179_));
 sky130_fd_sc_hd__nand3b_1 _07169_ (.A_N(_01176_),
    .B(_01178_),
    .C(_01179_),
    .Y(_01181_));
 sky130_fd_sc_hd__or2b_1 _07170_ (.A(_01174_),
    .B_N(_01175_),
    .X(_01182_));
 sky130_fd_sc_hd__or2b_1 _07171_ (.A(_01175_),
    .B_N(_01174_),
    .X(_01183_));
 sky130_fd_sc_hd__nand3_1 _07172_ (.A(_01182_),
    .B(_01183_),
    .C(_01177_),
    .Y(_01184_));
 sky130_fd_sc_hd__nand2_1 _07173_ (.A(_01181_),
    .B(_01184_),
    .Y(_01185_));
 sky130_fd_sc_hd__inv_2 _07174_ (.A(_01185_),
    .Y(_01186_));
 sky130_fd_sc_hd__inv_2 _07175_ (.A(_01033_),
    .Y(_01187_));
 sky130_fd_sc_hd__nand2_1 _07176_ (.A(_01187_),
    .B(_01034_),
    .Y(_01188_));
 sky130_fd_sc_hd__inv_2 _07177_ (.A(_01034_),
    .Y(_01189_));
 sky130_fd_sc_hd__nand2_1 _07178_ (.A(_01189_),
    .B(_01033_),
    .Y(_01190_));
 sky130_fd_sc_hd__nand3_1 _07179_ (.A(_01188_),
    .B(_01190_),
    .C(_01036_),
    .Y(_01192_));
 sky130_fd_sc_hd__nand2_1 _07180_ (.A(_01187_),
    .B(_01189_),
    .Y(_01193_));
 sky130_fd_sc_hd__nand3_1 _07181_ (.A(_01193_),
    .B(_01038_),
    .C(_01035_),
    .Y(_01194_));
 sky130_fd_sc_hd__nand2_2 _07182_ (.A(_01192_),
    .B(_01194_),
    .Y(_01195_));
 sky130_fd_sc_hd__nand2_1 _07183_ (.A(_03160_),
    .B(_00751_),
    .Y(_01196_));
 sky130_fd_sc_hd__nand2_1 _07184_ (.A(_02049_),
    .B(_02379_),
    .Y(_01197_));
 sky130_fd_sc_hd__nand2_2 _07185_ (.A(_01196_),
    .B(_01197_),
    .Y(_01198_));
 sky130_fd_sc_hd__nand2_1 _07186_ (.A(_03182_),
    .B(_00861_),
    .Y(_01199_));
 sky130_fd_sc_hd__inv_2 _07187_ (.A(_01199_),
    .Y(_01200_));
 sky130_fd_sc_hd__nor2_1 _07188_ (.A(_01196_),
    .B(_01197_),
    .Y(_01201_));
 sky130_fd_sc_hd__a21oi_4 _07189_ (.A1(_01198_),
    .A2(_01200_),
    .B1(_01201_),
    .Y(_01203_));
 sky130_fd_sc_hd__nand2_1 _07190_ (.A(_01195_),
    .B(_01203_),
    .Y(_01204_));
 sky130_fd_sc_hd__nor2_1 _07191_ (.A(_01203_),
    .B(_01195_),
    .Y(_01205_));
 sky130_fd_sc_hd__a21oi_2 _07192_ (.A1(_01186_),
    .A2(_01204_),
    .B1(_01205_),
    .Y(_01206_));
 sky130_fd_sc_hd__a21o_1 _07193_ (.A1(_01035_),
    .A2(_01038_),
    .B1(_01039_),
    .X(_01207_));
 sky130_fd_sc_hd__nand3_1 _07194_ (.A(_01207_),
    .B(_01031_),
    .C(_01029_),
    .Y(_01208_));
 sky130_fd_sc_hd__nand3_1 _07195_ (.A(_01208_),
    .B(_01041_),
    .C(_01056_),
    .Y(_01209_));
 sky130_fd_sc_hd__nand2_1 _07196_ (.A(_01032_),
    .B(_01207_),
    .Y(_01210_));
 sky130_fd_sc_hd__nand3_1 _07197_ (.A(_01040_),
    .B(_01029_),
    .C(_01031_),
    .Y(_01211_));
 sky130_fd_sc_hd__nand3_1 _07198_ (.A(_01210_),
    .B(_01211_),
    .C(_01055_),
    .Y(_01212_));
 sky130_fd_sc_hd__nand2_2 _07199_ (.A(_01209_),
    .B(_01212_),
    .Y(_01214_));
 sky130_fd_sc_hd__nor2_1 _07200_ (.A(_01206_),
    .B(_01214_),
    .Y(_01215_));
 sky130_fd_sc_hd__nand2_1 _07201_ (.A(_01214_),
    .B(_01206_),
    .Y(_01216_));
 sky130_fd_sc_hd__inv_2 _07202_ (.A(_01216_),
    .Y(_01217_));
 sky130_fd_sc_hd__nor2_1 _07203_ (.A(_01215_),
    .B(_01217_),
    .Y(_01218_));
 sky130_fd_sc_hd__a21o_1 _07204_ (.A1(_01179_),
    .A2(_01178_),
    .B1(_01176_),
    .X(_01219_));
 sky130_fd_sc_hd__nand2_1 _07205_ (.A(_01071_),
    .B(_01072_),
    .Y(_01220_));
 sky130_fd_sc_hd__nand2_1 _07206_ (.A(_01073_),
    .B(_01069_),
    .Y(_01221_));
 sky130_fd_sc_hd__nand3_1 _07207_ (.A(_01220_),
    .B(_01221_),
    .C(_01075_),
    .Y(_01222_));
 sky130_fd_sc_hd__nand3_1 _07208_ (.A(_01219_),
    .B(_01078_),
    .C(_01222_),
    .Y(_01223_));
 sky130_fd_sc_hd__nand2_1 _07209_ (.A(_01222_),
    .B(_01078_),
    .Y(_01225_));
 sky130_fd_sc_hd__a21oi_1 _07210_ (.A1(_01179_),
    .A2(_01178_),
    .B1(_01176_),
    .Y(_01226_));
 sky130_fd_sc_hd__nand2_1 _07211_ (.A(_01225_),
    .B(_01226_),
    .Y(_01227_));
 sky130_fd_sc_hd__nand2_1 _07212_ (.A(_01223_),
    .B(_01227_),
    .Y(_01228_));
 sky130_fd_sc_hd__nand2_1 _07213_ (.A(_03820_),
    .B(_01774_),
    .Y(_01229_));
 sky130_fd_sc_hd__nand2_1 _07214_ (.A(_03402_),
    .B(_01807_),
    .Y(_01230_));
 sky130_fd_sc_hd__nand2_1 _07215_ (.A(_01229_),
    .B(_01230_),
    .Y(_01231_));
 sky130_fd_sc_hd__nand2_1 _07216_ (.A(_04809_),
    .B(_01884_),
    .Y(_01232_));
 sky130_fd_sc_hd__inv_2 _07217_ (.A(_01232_),
    .Y(_01233_));
 sky130_fd_sc_hd__nor2_1 _07218_ (.A(_01229_),
    .B(_01230_),
    .Y(_01234_));
 sky130_fd_sc_hd__a21oi_1 _07219_ (.A1(_01231_),
    .A2(_01233_),
    .B1(_01234_),
    .Y(_01236_));
 sky130_fd_sc_hd__nand2_1 _07220_ (.A(_01228_),
    .B(_01236_),
    .Y(_01237_));
 sky130_fd_sc_hd__inv_2 _07221_ (.A(_01236_),
    .Y(_01238_));
 sky130_fd_sc_hd__nand3_1 _07222_ (.A(_01223_),
    .B(_01227_),
    .C(_01238_),
    .Y(_01239_));
 sky130_fd_sc_hd__nand2_1 _07223_ (.A(_01237_),
    .B(_01239_),
    .Y(_01240_));
 sky130_fd_sc_hd__inv_2 _07224_ (.A(_01240_),
    .Y(_01241_));
 sky130_fd_sc_hd__nand2_1 _07225_ (.A(_01218_),
    .B(_01241_),
    .Y(_01242_));
 sky130_fd_sc_hd__nand2b_1 _07226_ (.A_N(_01214_),
    .B(_01206_),
    .Y(_01243_));
 sky130_fd_sc_hd__inv_2 _07227_ (.A(_01206_),
    .Y(_01244_));
 sky130_fd_sc_hd__nand2_1 _07228_ (.A(_01244_),
    .B(_01214_),
    .Y(_01245_));
 sky130_fd_sc_hd__nand3_1 _07229_ (.A(_01243_),
    .B(_01245_),
    .C(_01240_),
    .Y(_01247_));
 sky130_fd_sc_hd__nand2_1 _07230_ (.A(_01242_),
    .B(_01247_),
    .Y(_01248_));
 sky130_fd_sc_hd__inv_2 _07231_ (.A(_01195_),
    .Y(_01249_));
 sky130_fd_sc_hd__inv_2 _07232_ (.A(_01203_),
    .Y(_01250_));
 sky130_fd_sc_hd__nand2_1 _07233_ (.A(_01249_),
    .B(_01250_),
    .Y(_01251_));
 sky130_fd_sc_hd__nand3_1 _07234_ (.A(_01251_),
    .B(_01186_),
    .C(_01204_),
    .Y(_01252_));
 sky130_fd_sc_hd__nand2_1 _07235_ (.A(_01249_),
    .B(_01203_),
    .Y(_01253_));
 sky130_fd_sc_hd__nand2_1 _07236_ (.A(_01195_),
    .B(_01250_),
    .Y(_01254_));
 sky130_fd_sc_hd__nand3_1 _07237_ (.A(_01253_),
    .B(_01185_),
    .C(_01254_),
    .Y(_01255_));
 sky130_fd_sc_hd__nand2_1 _07238_ (.A(_01252_),
    .B(_01255_),
    .Y(_01256_));
 sky130_fd_sc_hd__inv_2 _07239_ (.A(_01198_),
    .Y(_01258_));
 sky130_fd_sc_hd__o21ai_1 _07240_ (.A1(_01201_),
    .A2(_01258_),
    .B1(_01199_),
    .Y(_01259_));
 sky130_fd_sc_hd__nand3b_1 _07241_ (.A_N(_01201_),
    .B(_01200_),
    .C(_01198_),
    .Y(_01260_));
 sky130_fd_sc_hd__nand2_1 _07242_ (.A(_01259_),
    .B(_01260_),
    .Y(_01261_));
 sky130_fd_sc_hd__nand2_1 _07243_ (.A(_03182_),
    .B(_00751_),
    .Y(_01262_));
 sky130_fd_sc_hd__nand2_1 _07244_ (.A(_03160_),
    .B(_00795_),
    .Y(_01263_));
 sky130_fd_sc_hd__nand2_1 _07245_ (.A(_01262_),
    .B(_01263_),
    .Y(_01264_));
 sky130_fd_sc_hd__nand2_1 _07246_ (.A(_05031_),
    .B(_00861_),
    .Y(_01265_));
 sky130_fd_sc_hd__inv_2 _07247_ (.A(_01265_),
    .Y(_01266_));
 sky130_fd_sc_hd__nor2_1 _07248_ (.A(_01262_),
    .B(_01263_),
    .Y(_01267_));
 sky130_fd_sc_hd__a21oi_2 _07249_ (.A1(_01264_),
    .A2(_01266_),
    .B1(_01267_),
    .Y(_01269_));
 sky130_fd_sc_hd__nand2_1 _07250_ (.A(_01261_),
    .B(_01269_),
    .Y(_01270_));
 sky130_fd_sc_hd__nand2_1 _07251_ (.A(_05028_),
    .B(_04260_),
    .Y(_01271_));
 sky130_fd_sc_hd__nand2_1 _07252_ (.A(_05031_),
    .B(_01092_),
    .Y(_01272_));
 sky130_fd_sc_hd__nor2_1 _07253_ (.A(_01271_),
    .B(_01272_),
    .Y(_01273_));
 sky130_fd_sc_hd__nand2_1 _07254_ (.A(_01271_),
    .B(_01272_),
    .Y(_01274_));
 sky130_fd_sc_hd__inv_2 _07255_ (.A(_01274_),
    .Y(_01275_));
 sky130_fd_sc_hd__nand2_1 _07256_ (.A(_04928_),
    .B(_01158_),
    .Y(_01276_));
 sky130_fd_sc_hd__o21ai_1 _07257_ (.A1(_01273_),
    .A2(_01275_),
    .B1(_01276_),
    .Y(_01277_));
 sky130_fd_sc_hd__inv_2 _07258_ (.A(_01276_),
    .Y(_01278_));
 sky130_fd_sc_hd__nand3b_1 _07259_ (.A_N(_01273_),
    .B(_01278_),
    .C(_01274_),
    .Y(_01280_));
 sky130_fd_sc_hd__nand2_1 _07260_ (.A(_01277_),
    .B(_01280_),
    .Y(_01281_));
 sky130_fd_sc_hd__inv_2 _07261_ (.A(_01281_),
    .Y(_01282_));
 sky130_fd_sc_hd__nor2_1 _07262_ (.A(_01269_),
    .B(_01261_),
    .Y(_01283_));
 sky130_fd_sc_hd__a21oi_2 _07263_ (.A1(_01270_),
    .A2(_01282_),
    .B1(_01283_),
    .Y(_01284_));
 sky130_fd_sc_hd__nand2_1 _07264_ (.A(_01256_),
    .B(_01284_),
    .Y(_01285_));
 sky130_fd_sc_hd__nand2_1 _07265_ (.A(_00254_),
    .B(_00412_),
    .Y(_01286_));
 sky130_fd_sc_hd__nand2_1 _07266_ (.A(_00656_),
    .B(_00204_),
    .Y(_01287_));
 sky130_fd_sc_hd__nand2_1 _07267_ (.A(_01286_),
    .B(_01287_),
    .Y(_01288_));
 sky130_fd_sc_hd__nand2_1 _07268_ (.A(_00522_),
    .B(_00003_),
    .Y(_01289_));
 sky130_fd_sc_hd__inv_2 _07269_ (.A(_01289_),
    .Y(_01291_));
 sky130_fd_sc_hd__nor2_1 _07270_ (.A(_01286_),
    .B(_01287_),
    .Y(_01292_));
 sky130_fd_sc_hd__a21o_1 _07271_ (.A1(_01288_),
    .A2(_01291_),
    .B1(_01292_),
    .X(_01293_));
 sky130_fd_sc_hd__inv_2 _07272_ (.A(_01231_),
    .Y(_01294_));
 sky130_fd_sc_hd__o21ai_1 _07273_ (.A1(_01234_),
    .A2(_01294_),
    .B1(_01232_),
    .Y(_01295_));
 sky130_fd_sc_hd__nor2_1 _07274_ (.A(_01234_),
    .B(_01294_),
    .Y(_01296_));
 sky130_fd_sc_hd__nand2_1 _07275_ (.A(_01296_),
    .B(_01233_),
    .Y(_01297_));
 sky130_fd_sc_hd__nand2_1 _07276_ (.A(_01295_),
    .B(_01297_),
    .Y(_01298_));
 sky130_fd_sc_hd__a21oi_2 _07277_ (.A1(_01274_),
    .A2(_01278_),
    .B1(_01273_),
    .Y(_01299_));
 sky130_fd_sc_hd__inv_2 _07278_ (.A(_01299_),
    .Y(_01300_));
 sky130_fd_sc_hd__nand2_1 _07279_ (.A(_01298_),
    .B(_01300_),
    .Y(_01302_));
 sky130_fd_sc_hd__nand3_1 _07280_ (.A(_01295_),
    .B(_01297_),
    .C(_01299_),
    .Y(_01303_));
 sky130_fd_sc_hd__nand3b_1 _07281_ (.A_N(_01293_),
    .B(_01302_),
    .C(_01303_),
    .Y(_01304_));
 sky130_fd_sc_hd__nand2_1 _07282_ (.A(_01298_),
    .B(_01299_),
    .Y(_01305_));
 sky130_fd_sc_hd__nand3_1 _07283_ (.A(_01295_),
    .B(_01300_),
    .C(_01297_),
    .Y(_01306_));
 sky130_fd_sc_hd__nand3_1 _07284_ (.A(_01305_),
    .B(_01306_),
    .C(_01293_),
    .Y(_01307_));
 sky130_fd_sc_hd__nand2_1 _07285_ (.A(_01304_),
    .B(_01307_),
    .Y(_01308_));
 sky130_fd_sc_hd__inv_2 _07286_ (.A(_01308_),
    .Y(_01309_));
 sky130_fd_sc_hd__nor2_1 _07287_ (.A(_01284_),
    .B(_01256_),
    .Y(_01310_));
 sky130_fd_sc_hd__a21oi_1 _07288_ (.A1(_01285_),
    .A2(_01309_),
    .B1(_01310_),
    .Y(_01311_));
 sky130_fd_sc_hd__nand2_1 _07289_ (.A(_01248_),
    .B(_01311_),
    .Y(_01313_));
 sky130_fd_sc_hd__inv_2 _07290_ (.A(_01106_),
    .Y(_01314_));
 sky130_fd_sc_hd__o21ai_1 _07291_ (.A1(_01109_),
    .A2(_01314_),
    .B1(_01107_),
    .Y(_01315_));
 sky130_fd_sc_hd__nand3b_1 _07292_ (.A_N(_01109_),
    .B(_01108_),
    .C(_01106_),
    .Y(_01316_));
 sky130_fd_sc_hd__nand2_1 _07293_ (.A(_01315_),
    .B(_01316_),
    .Y(_01317_));
 sky130_fd_sc_hd__nand2_1 _07294_ (.A(_04827_),
    .B(_05029_),
    .Y(_01318_));
 sky130_fd_sc_hd__nand2_1 _07295_ (.A(_00522_),
    .B(_05032_),
    .Y(_01319_));
 sky130_fd_sc_hd__nand2_1 _07296_ (.A(_01318_),
    .B(_01319_),
    .Y(_01320_));
 sky130_fd_sc_hd__nand2_1 _07297_ (.A(_03215_),
    .B(_04911_),
    .Y(_01321_));
 sky130_fd_sc_hd__inv_2 _07298_ (.A(_01321_),
    .Y(_01322_));
 sky130_fd_sc_hd__nor2_1 _07299_ (.A(_01318_),
    .B(_01319_),
    .Y(_01324_));
 sky130_fd_sc_hd__a21oi_2 _07300_ (.A1(_01320_),
    .A2(_01322_),
    .B1(_01324_),
    .Y(_01325_));
 sky130_fd_sc_hd__inv_2 _07301_ (.A(_01325_),
    .Y(_01326_));
 sky130_fd_sc_hd__nand2_1 _07302_ (.A(_01317_),
    .B(_01326_),
    .Y(_01327_));
 sky130_fd_sc_hd__nand3_1 _07303_ (.A(_01315_),
    .B(_01316_),
    .C(_01325_),
    .Y(_01328_));
 sky130_fd_sc_hd__nand2_1 _07304_ (.A(_01327_),
    .B(_01328_),
    .Y(_01329_));
 sky130_fd_sc_hd__clkinv_4 _07305_ (.A(net36),
    .Y(_01330_));
 sky130_fd_sc_hd__nand2_1 _07306_ (.A(_04962_),
    .B(_04895_),
    .Y(_01331_));
 sky130_fd_sc_hd__nor3_1 _07307_ (.A(_01330_),
    .B(_00264_),
    .C(_01331_),
    .Y(_01332_));
 sky130_fd_sc_hd__inv_2 _07308_ (.A(_01332_),
    .Y(_01333_));
 sky130_fd_sc_hd__o21ai_1 _07309_ (.A1(_01330_),
    .A2(_00264_),
    .B1(_01331_),
    .Y(_01335_));
 sky130_fd_sc_hd__nand2_1 _07310_ (.A(_01333_),
    .B(_01335_),
    .Y(_01336_));
 sky130_fd_sc_hd__inv_2 _07311_ (.A(_01336_),
    .Y(_01337_));
 sky130_fd_sc_hd__nand2_1 _07312_ (.A(_01329_),
    .B(_01337_),
    .Y(_01338_));
 sky130_fd_sc_hd__nand3_1 _07313_ (.A(_01327_),
    .B(_01328_),
    .C(_01336_),
    .Y(_01339_));
 sky130_fd_sc_hd__nand2_1 _07314_ (.A(_01338_),
    .B(_01339_),
    .Y(_01340_));
 sky130_fd_sc_hd__nor2_1 _07315_ (.A(_01299_),
    .B(_01298_),
    .Y(_01341_));
 sky130_fd_sc_hd__a21oi_2 _07316_ (.A1(_01305_),
    .A2(_01293_),
    .B1(_01341_),
    .Y(_01342_));
 sky130_fd_sc_hd__inv_2 _07317_ (.A(_01342_),
    .Y(_01343_));
 sky130_fd_sc_hd__nand2_1 _07318_ (.A(_01340_),
    .B(_01343_),
    .Y(_01344_));
 sky130_fd_sc_hd__nand3_1 _07319_ (.A(_01342_),
    .B(_01338_),
    .C(_01339_),
    .Y(_01346_));
 sky130_fd_sc_hd__nand2_1 _07320_ (.A(_01344_),
    .B(_01346_),
    .Y(_01347_));
 sky130_fd_sc_hd__inv_2 _07321_ (.A(_01324_),
    .Y(_01348_));
 sky130_fd_sc_hd__a21o_1 _07322_ (.A1(_01348_),
    .A2(_01320_),
    .B1(_01322_),
    .X(_01349_));
 sky130_fd_sc_hd__nand3_1 _07323_ (.A(_01348_),
    .B(_01322_),
    .C(_01320_),
    .Y(_01350_));
 sky130_fd_sc_hd__nand2_1 _07324_ (.A(_01349_),
    .B(_01350_),
    .Y(_01351_));
 sky130_fd_sc_hd__nand2_1 _07325_ (.A(_04911_),
    .B(_05029_),
    .Y(_01352_));
 sky130_fd_sc_hd__nand2_1 _07326_ (.A(_04828_),
    .B(_05032_),
    .Y(_01353_));
 sky130_fd_sc_hd__nand2_1 _07327_ (.A(_01352_),
    .B(_01353_),
    .Y(_01354_));
 sky130_fd_sc_hd__nand2_1 _07328_ (.A(_03215_),
    .B(_04895_),
    .Y(_01355_));
 sky130_fd_sc_hd__inv_2 _07329_ (.A(_01355_),
    .Y(_01357_));
 sky130_fd_sc_hd__nor2_1 _07330_ (.A(_01352_),
    .B(_01353_),
    .Y(_01358_));
 sky130_fd_sc_hd__a21oi_2 _07331_ (.A1(_01354_),
    .A2(_01357_),
    .B1(_01358_),
    .Y(_01359_));
 sky130_fd_sc_hd__nand2_1 _07332_ (.A(_01351_),
    .B(_01359_),
    .Y(_01360_));
 sky130_fd_sc_hd__nand2_1 _07333_ (.A(_04964_),
    .B(_04895_),
    .Y(_01361_));
 sky130_fd_sc_hd__inv_2 _07334_ (.A(_01361_),
    .Y(_01362_));
 sky130_fd_sc_hd__nor2_1 _07335_ (.A(_01359_),
    .B(_01351_),
    .Y(_01363_));
 sky130_fd_sc_hd__a21oi_1 _07336_ (.A1(_01360_),
    .A2(_01362_),
    .B1(_01363_),
    .Y(_01364_));
 sky130_fd_sc_hd__inv_2 _07337_ (.A(_01364_),
    .Y(_01365_));
 sky130_fd_sc_hd__nand2_1 _07338_ (.A(_01347_),
    .B(_01365_),
    .Y(_01366_));
 sky130_fd_sc_hd__nand3_1 _07339_ (.A(_01344_),
    .B(_01346_),
    .C(_01364_),
    .Y(_01368_));
 sky130_fd_sc_hd__nand2_1 _07340_ (.A(_01366_),
    .B(_01368_),
    .Y(_01369_));
 sky130_fd_sc_hd__inv_2 _07341_ (.A(_01369_),
    .Y(_01370_));
 sky130_fd_sc_hd__nor2_1 _07342_ (.A(_01311_),
    .B(_01248_),
    .Y(_01371_));
 sky130_fd_sc_hd__a21oi_1 _07343_ (.A1(_01313_),
    .A2(_01370_),
    .B1(_01371_),
    .Y(_01372_));
 sky130_fd_sc_hd__a21oi_1 _07344_ (.A1(_01216_),
    .A2(_01241_),
    .B1(_01215_),
    .Y(_01373_));
 sky130_fd_sc_hd__nand3_1 _07345_ (.A(_01058_),
    .B(_01012_),
    .C(_01022_),
    .Y(_01374_));
 sky130_fd_sc_hd__nand2_1 _07346_ (.A(_01209_),
    .B(_01208_),
    .Y(_01375_));
 sky130_fd_sc_hd__nand2_1 _07347_ (.A(_01023_),
    .B(_01375_),
    .Y(_01376_));
 sky130_fd_sc_hd__nand2_1 _07348_ (.A(_01374_),
    .B(_01376_),
    .Y(_01377_));
 sky130_fd_sc_hd__nand2_1 _07349_ (.A(_01377_),
    .B(_01087_),
    .Y(_01379_));
 sky130_fd_sc_hd__nand3_1 _07350_ (.A(_01374_),
    .B(_01376_),
    .C(_01086_),
    .Y(_01380_));
 sky130_fd_sc_hd__nand3_1 _07351_ (.A(_01373_),
    .B(_01379_),
    .C(_01380_),
    .Y(_01381_));
 sky130_fd_sc_hd__nand2_1 _07352_ (.A(_01379_),
    .B(_01380_),
    .Y(_01382_));
 sky130_fd_sc_hd__a21o_1 _07353_ (.A1(_01216_),
    .A2(_01241_),
    .B1(_01215_),
    .X(_01383_));
 sky130_fd_sc_hd__nand2_1 _07354_ (.A(_01382_),
    .B(_01383_),
    .Y(_01384_));
 sky130_fd_sc_hd__nand2_1 _07355_ (.A(_01381_),
    .B(_01384_),
    .Y(_01385_));
 sky130_fd_sc_hd__nand2_1 _07356_ (.A(_01119_),
    .B(_01122_),
    .Y(_01386_));
 sky130_fd_sc_hd__nand2_1 _07357_ (.A(_01386_),
    .B(_01102_),
    .Y(_01387_));
 sky130_fd_sc_hd__nand2_1 _07358_ (.A(_01387_),
    .B(_01123_),
    .Y(_01388_));
 sky130_fd_sc_hd__nor2_1 _07359_ (.A(_01226_),
    .B(_01225_),
    .Y(_01390_));
 sky130_fd_sc_hd__a21oi_2 _07360_ (.A1(_01227_),
    .A2(_01238_),
    .B1(_01390_),
    .Y(_01391_));
 sky130_fd_sc_hd__inv_2 _07361_ (.A(_01391_),
    .Y(_01392_));
 sky130_fd_sc_hd__nand2_1 _07362_ (.A(_01388_),
    .B(_01392_),
    .Y(_01393_));
 sky130_fd_sc_hd__nand3_1 _07363_ (.A(_01391_),
    .B(_01387_),
    .C(_01123_),
    .Y(_01394_));
 sky130_fd_sc_hd__nand2_1 _07364_ (.A(_01393_),
    .B(_01394_),
    .Y(_01395_));
 sky130_fd_sc_hd__nand2_1 _07365_ (.A(_01317_),
    .B(_01325_),
    .Y(_01396_));
 sky130_fd_sc_hd__nor2_1 _07366_ (.A(_01325_),
    .B(_01317_),
    .Y(_01397_));
 sky130_fd_sc_hd__a21oi_1 _07367_ (.A1(_01396_),
    .A2(_01337_),
    .B1(_01397_),
    .Y(_01398_));
 sky130_fd_sc_hd__inv_2 _07368_ (.A(_01398_),
    .Y(_01399_));
 sky130_fd_sc_hd__nand2_1 _07369_ (.A(_01395_),
    .B(_01399_),
    .Y(_01401_));
 sky130_fd_sc_hd__nand3_1 _07370_ (.A(_01393_),
    .B(_01394_),
    .C(_01398_),
    .Y(_01402_));
 sky130_fd_sc_hd__nand2_1 _07371_ (.A(_01401_),
    .B(_01402_),
    .Y(_01403_));
 sky130_fd_sc_hd__inv_2 _07372_ (.A(_01403_),
    .Y(_01404_));
 sky130_fd_sc_hd__nand2_1 _07373_ (.A(_01385_),
    .B(_01404_),
    .Y(_01405_));
 sky130_fd_sc_hd__nand3_1 _07374_ (.A(_01381_),
    .B(_01384_),
    .C(_01403_),
    .Y(_01406_));
 sky130_fd_sc_hd__nand2_1 _07375_ (.A(_01405_),
    .B(_01406_),
    .Y(_01407_));
 sky130_fd_sc_hd__nand2_1 _07376_ (.A(_01372_),
    .B(_01407_),
    .Y(_01408_));
 sky130_fd_sc_hd__or2_1 _07377_ (.A(_01342_),
    .B(_01340_),
    .X(_01409_));
 sky130_fd_sc_hd__and2_1 _07378_ (.A(_01366_),
    .B(_01409_),
    .X(_01410_));
 sky130_fd_sc_hd__nor2_2 _07379_ (.A(_01333_),
    .B(_01410_),
    .Y(_01412_));
 sky130_fd_sc_hd__nand2_1 _07380_ (.A(_01410_),
    .B(_01333_),
    .Y(_01413_));
 sky130_fd_sc_hd__nor2b_1 _07381_ (.A(_01412_),
    .B_N(_01413_),
    .Y(_01414_));
 sky130_fd_sc_hd__nor2_1 _07382_ (.A(_01407_),
    .B(_01372_),
    .Y(_01415_));
 sky130_fd_sc_hd__a21oi_2 _07383_ (.A1(_01408_),
    .A2(_01414_),
    .B1(_01415_),
    .Y(_01416_));
 sky130_fd_sc_hd__inv_2 _07384_ (.A(_01416_),
    .Y(_01417_));
 sky130_fd_sc_hd__nand2_1 _07385_ (.A(_01382_),
    .B(_01373_),
    .Y(_01418_));
 sky130_fd_sc_hd__nor2_1 _07386_ (.A(_01373_),
    .B(_01382_),
    .Y(_01419_));
 sky130_fd_sc_hd__a21oi_1 _07387_ (.A1(_01418_),
    .A2(_01404_),
    .B1(_01419_),
    .Y(_01420_));
 sky130_fd_sc_hd__a21o_1 _07388_ (.A1(_01060_),
    .A2(_01087_),
    .B1(_01088_),
    .X(_01421_));
 sky130_fd_sc_hd__nand3_1 _07389_ (.A(_01421_),
    .B(_01017_),
    .C(_01018_),
    .Y(_01423_));
 sky130_fd_sc_hd__nand3_2 _07390_ (.A(_01423_),
    .B(_01129_),
    .C(_01090_),
    .Y(_01424_));
 sky130_fd_sc_hd__nand2_1 _07391_ (.A(_01019_),
    .B(_01421_),
    .Y(_01425_));
 sky130_fd_sc_hd__nand3_1 _07392_ (.A(_01089_),
    .B(_01017_),
    .C(_01018_),
    .Y(_01426_));
 sky130_fd_sc_hd__nand3_1 _07393_ (.A(_01425_),
    .B(_01426_),
    .C(_01128_),
    .Y(_01427_));
 sky130_fd_sc_hd__nand3_1 _07394_ (.A(_01420_),
    .B(_01424_),
    .C(_01427_),
    .Y(_01428_));
 sky130_fd_sc_hd__nand2_1 _07395_ (.A(_01424_),
    .B(_01427_),
    .Y(_01429_));
 sky130_fd_sc_hd__a21o_1 _07396_ (.A1(_01418_),
    .A2(_01404_),
    .B1(_01419_),
    .X(_01430_));
 sky130_fd_sc_hd__nand2_1 _07397_ (.A(_01429_),
    .B(_01430_),
    .Y(_01431_));
 sky130_fd_sc_hd__nand2_1 _07398_ (.A(_01428_),
    .B(_01431_),
    .Y(_01432_));
 sky130_fd_sc_hd__nand2_1 _07399_ (.A(_00972_),
    .B(_00962_),
    .Y(_01434_));
 sky130_fd_sc_hd__nand2_2 _07400_ (.A(_00974_),
    .B(_01434_),
    .Y(_01435_));
 sky130_fd_sc_hd__o21a_1 _07401_ (.A1(_01388_),
    .A2(_01391_),
    .B1(_01401_),
    .X(_01436_));
 sky130_fd_sc_hd__xor2_2 _07402_ (.A(_01435_),
    .B(_01436_),
    .X(_01437_));
 sky130_fd_sc_hd__nand2_1 _07403_ (.A(_01432_),
    .B(_01437_),
    .Y(_01438_));
 sky130_fd_sc_hd__nand3b_1 _07404_ (.A_N(_01437_),
    .B(_01428_),
    .C(_01431_),
    .Y(_01439_));
 sky130_fd_sc_hd__nand2_1 _07405_ (.A(_01438_),
    .B(_01439_),
    .Y(_01440_));
 sky130_fd_sc_hd__nand2_1 _07406_ (.A(_01417_),
    .B(_01440_),
    .Y(_01441_));
 sky130_fd_sc_hd__nand3_1 _07407_ (.A(_01416_),
    .B(_01438_),
    .C(_01439_),
    .Y(_01442_));
 sky130_fd_sc_hd__nand2_1 _07408_ (.A(_01441_),
    .B(_01442_),
    .Y(_01443_));
 sky130_fd_sc_hd__nand2_1 _07409_ (.A(_01443_),
    .B(_01412_),
    .Y(_01445_));
 sky130_fd_sc_hd__inv_2 _07410_ (.A(_01412_),
    .Y(_01446_));
 sky130_fd_sc_hd__nand3_1 _07411_ (.A(_01441_),
    .B(_01442_),
    .C(_01446_),
    .Y(_01447_));
 sky130_fd_sc_hd__nand2_1 _07412_ (.A(_01445_),
    .B(_01447_),
    .Y(_01448_));
 sky130_fd_sc_hd__a21o_1 _07413_ (.A1(_01285_),
    .A2(_01309_),
    .B1(_01310_),
    .X(_01449_));
 sky130_fd_sc_hd__nand3_1 _07414_ (.A(_01449_),
    .B(_01242_),
    .C(_01247_),
    .Y(_01450_));
 sky130_fd_sc_hd__nand3_1 _07415_ (.A(_01450_),
    .B(_01313_),
    .C(_01370_),
    .Y(_01451_));
 sky130_fd_sc_hd__nand2_1 _07416_ (.A(_01248_),
    .B(_01449_),
    .Y(_01452_));
 sky130_fd_sc_hd__nand3_1 _07417_ (.A(_01311_),
    .B(_01242_),
    .C(_01247_),
    .Y(_01453_));
 sky130_fd_sc_hd__nand3_1 _07418_ (.A(_01452_),
    .B(_01453_),
    .C(_01369_),
    .Y(_01454_));
 sky130_fd_sc_hd__nand2_1 _07419_ (.A(_01451_),
    .B(_01454_),
    .Y(_01456_));
 sky130_fd_sc_hd__inv_2 _07420_ (.A(_01456_),
    .Y(_01457_));
 sky130_fd_sc_hd__inv_2 _07421_ (.A(_01288_),
    .Y(_01458_));
 sky130_fd_sc_hd__o21ai_1 _07422_ (.A1(_01292_),
    .A2(_01458_),
    .B1(_01289_),
    .Y(_01459_));
 sky130_fd_sc_hd__nand3b_1 _07423_ (.A_N(_01292_),
    .B(_01291_),
    .C(_01288_),
    .Y(_01460_));
 sky130_fd_sc_hd__nand2_1 _07424_ (.A(_01459_),
    .B(_01460_),
    .Y(_01461_));
 sky130_fd_sc_hd__nand2_1 _07425_ (.A(_03402_),
    .B(_01048_),
    .Y(_01462_));
 sky130_fd_sc_hd__nand2_1 _07426_ (.A(_03314_),
    .B(_01092_),
    .Y(_01463_));
 sky130_fd_sc_hd__nand2_1 _07427_ (.A(_01462_),
    .B(_01463_),
    .Y(_01464_));
 sky130_fd_sc_hd__nand2_1 _07428_ (.A(_00656_),
    .B(_01565_),
    .Y(_01465_));
 sky130_fd_sc_hd__inv_2 _07429_ (.A(_01465_),
    .Y(_01467_));
 sky130_fd_sc_hd__nor2_1 _07430_ (.A(_01462_),
    .B(_01463_),
    .Y(_01468_));
 sky130_fd_sc_hd__a21oi_2 _07431_ (.A1(_01464_),
    .A2(_01467_),
    .B1(_01468_),
    .Y(_01469_));
 sky130_fd_sc_hd__nand2_1 _07432_ (.A(_01461_),
    .B(_01469_),
    .Y(_01470_));
 sky130_fd_sc_hd__nand2_1 _07433_ (.A(_00522_),
    .B(_00412_),
    .Y(_01471_));
 sky130_fd_sc_hd__inv_2 _07434_ (.A(_01471_),
    .Y(_01472_));
 sky130_fd_sc_hd__nand2_1 _07435_ (.A(_00254_),
    .B(_00204_),
    .Y(_01473_));
 sky130_fd_sc_hd__inv_2 _07436_ (.A(_01473_),
    .Y(_01474_));
 sky130_fd_sc_hd__nand2_1 _07437_ (.A(_01472_),
    .B(_01474_),
    .Y(_01475_));
 sky130_fd_sc_hd__nand2_1 _07438_ (.A(_04828_),
    .B(_00003_),
    .Y(_01476_));
 sky130_fd_sc_hd__inv_2 _07439_ (.A(_01476_),
    .Y(_01478_));
 sky130_fd_sc_hd__nand2_1 _07440_ (.A(_01471_),
    .B(_01473_),
    .Y(_01479_));
 sky130_fd_sc_hd__nand3_1 _07441_ (.A(_01475_),
    .B(_01478_),
    .C(_01479_),
    .Y(_01480_));
 sky130_fd_sc_hd__nand2_1 _07442_ (.A(_01480_),
    .B(_01475_),
    .Y(_01481_));
 sky130_fd_sc_hd__nor2_1 _07443_ (.A(_01469_),
    .B(_01461_),
    .Y(_01482_));
 sky130_fd_sc_hd__a21oi_1 _07444_ (.A1(_01470_),
    .A2(_01481_),
    .B1(_01482_),
    .Y(_01483_));
 sky130_fd_sc_hd__inv_2 _07445_ (.A(_01483_),
    .Y(_01484_));
 sky130_fd_sc_hd__inv_2 _07446_ (.A(_01359_),
    .Y(_01485_));
 sky130_fd_sc_hd__nand2_1 _07447_ (.A(_01351_),
    .B(_01485_),
    .Y(_01486_));
 sky130_fd_sc_hd__nand3_1 _07448_ (.A(_01349_),
    .B(_01359_),
    .C(_01350_),
    .Y(_01487_));
 sky130_fd_sc_hd__nand2_1 _07449_ (.A(_01486_),
    .B(_01487_),
    .Y(_01489_));
 sky130_fd_sc_hd__nand2_1 _07450_ (.A(_01489_),
    .B(_01362_),
    .Y(_01490_));
 sky130_fd_sc_hd__nand3_1 _07451_ (.A(_01486_),
    .B(_01361_),
    .C(_01487_),
    .Y(_01491_));
 sky130_fd_sc_hd__nand3_1 _07452_ (.A(_01484_),
    .B(_01490_),
    .C(_01491_),
    .Y(_01492_));
 sky130_fd_sc_hd__nand2_1 _07453_ (.A(_01490_),
    .B(_01491_),
    .Y(_01493_));
 sky130_fd_sc_hd__nand2_1 _07454_ (.A(_01493_),
    .B(_01483_),
    .Y(_01494_));
 sky130_fd_sc_hd__nand2_1 _07455_ (.A(_01492_),
    .B(_01494_),
    .Y(_01495_));
 sky130_fd_sc_hd__and4_1 _07456_ (.A(_04991_),
    .B(_04895_),
    .C(_05032_),
    .D(_05029_),
    .X(_01496_));
 sky130_fd_sc_hd__inv_2 _07457_ (.A(_01496_),
    .Y(_01497_));
 sky130_fd_sc_hd__nor2b_1 _07458_ (.A(_01358_),
    .B_N(_01354_),
    .Y(_01498_));
 sky130_fd_sc_hd__xor2_1 _07459_ (.A(_01355_),
    .B(_01498_),
    .X(_01500_));
 sky130_fd_sc_hd__nor2_1 _07460_ (.A(_01497_),
    .B(_01500_),
    .Y(_01501_));
 sky130_fd_sc_hd__inv_2 _07461_ (.A(_01501_),
    .Y(_01502_));
 sky130_fd_sc_hd__nand2_1 _07462_ (.A(_01495_),
    .B(_01502_),
    .Y(_01503_));
 sky130_fd_sc_hd__nand3_1 _07463_ (.A(_01492_),
    .B(_01494_),
    .C(_01501_),
    .Y(_01504_));
 sky130_fd_sc_hd__nand2_1 _07464_ (.A(_01503_),
    .B(_01504_),
    .Y(_01505_));
 sky130_fd_sc_hd__inv_2 _07465_ (.A(_01505_),
    .Y(_01506_));
 sky130_fd_sc_hd__nand3_1 _07466_ (.A(_01284_),
    .B(_01252_),
    .C(_01255_),
    .Y(_01507_));
 sky130_fd_sc_hd__inv_2 _07467_ (.A(_01284_),
    .Y(_01508_));
 sky130_fd_sc_hd__nand2_1 _07468_ (.A(_01508_),
    .B(_01256_),
    .Y(_01509_));
 sky130_fd_sc_hd__nand2_1 _07469_ (.A(_01507_),
    .B(_01509_),
    .Y(_01511_));
 sky130_fd_sc_hd__nand2_1 _07470_ (.A(_01511_),
    .B(_01309_),
    .Y(_01512_));
 sky130_fd_sc_hd__nand3_1 _07471_ (.A(_01507_),
    .B(_01509_),
    .C(_01308_),
    .Y(_01513_));
 sky130_fd_sc_hd__nand2_1 _07472_ (.A(_01512_),
    .B(_01513_),
    .Y(_01514_));
 sky130_fd_sc_hd__inv_2 _07473_ (.A(_01269_),
    .Y(_01515_));
 sky130_fd_sc_hd__nand2_1 _07474_ (.A(_01261_),
    .B(_01515_),
    .Y(_01516_));
 sky130_fd_sc_hd__nand3_1 _07475_ (.A(_01259_),
    .B(_01260_),
    .C(_01269_),
    .Y(_01517_));
 sky130_fd_sc_hd__nand2_1 _07476_ (.A(_01516_),
    .B(_01517_),
    .Y(_01518_));
 sky130_fd_sc_hd__nand2_1 _07477_ (.A(_01518_),
    .B(_01282_),
    .Y(_01519_));
 sky130_fd_sc_hd__nand3_1 _07478_ (.A(_01516_),
    .B(_01517_),
    .C(_01281_),
    .Y(_01520_));
 sky130_fd_sc_hd__nand2_1 _07479_ (.A(_01519_),
    .B(_01520_),
    .Y(_01522_));
 sky130_fd_sc_hd__inv_2 _07480_ (.A(_01468_),
    .Y(_01523_));
 sky130_fd_sc_hd__nand2_1 _07481_ (.A(_01523_),
    .B(_01464_),
    .Y(_01524_));
 sky130_fd_sc_hd__nand2_1 _07482_ (.A(_01524_),
    .B(_01465_),
    .Y(_01525_));
 sky130_fd_sc_hd__nand3_1 _07483_ (.A(_01523_),
    .B(_01467_),
    .C(_01464_),
    .Y(_01526_));
 sky130_fd_sc_hd__nand2_1 _07484_ (.A(_01525_),
    .B(_01526_),
    .Y(_01527_));
 sky130_fd_sc_hd__inv_2 _07485_ (.A(_01527_),
    .Y(_01528_));
 sky130_fd_sc_hd__inv_2 _07486_ (.A(_01267_),
    .Y(_01529_));
 sky130_fd_sc_hd__nand2_1 _07487_ (.A(_01529_),
    .B(_01264_),
    .Y(_01530_));
 sky130_fd_sc_hd__nand2_1 _07488_ (.A(_01530_),
    .B(_01265_),
    .Y(_01531_));
 sky130_fd_sc_hd__nand3_1 _07489_ (.A(_01529_),
    .B(_01266_),
    .C(_01264_),
    .Y(_01533_));
 sky130_fd_sc_hd__nand2_1 _07490_ (.A(_01531_),
    .B(_01533_),
    .Y(_01534_));
 sky130_fd_sc_hd__clkbuf_8 _07491_ (.A(_00861_),
    .X(_01535_));
 sky130_fd_sc_hd__nand2_1 _07492_ (.A(_05028_),
    .B(_01535_),
    .Y(_01536_));
 sky130_fd_sc_hd__nand2_1 _07493_ (.A(_05031_),
    .B(_00751_),
    .Y(_01537_));
 sky130_fd_sc_hd__nand2_1 _07494_ (.A(_03182_),
    .B(_00795_),
    .Y(_01538_));
 sky130_fd_sc_hd__nand2_1 _07495_ (.A(_01537_),
    .B(_01538_),
    .Y(_01539_));
 sky130_fd_sc_hd__inv_2 _07496_ (.A(_01539_),
    .Y(_01540_));
 sky130_fd_sc_hd__inv_2 _07497_ (.A(_01537_),
    .Y(_01541_));
 sky130_fd_sc_hd__inv_2 _07498_ (.A(_01538_),
    .Y(_01542_));
 sky130_fd_sc_hd__nand2_1 _07499_ (.A(_01541_),
    .B(_01542_),
    .Y(_01544_));
 sky130_fd_sc_hd__o21a_1 _07500_ (.A1(_01536_),
    .A2(_01540_),
    .B1(_01544_),
    .X(_01545_));
 sky130_fd_sc_hd__nand2_1 _07501_ (.A(_01534_),
    .B(_01545_),
    .Y(_01546_));
 sky130_fd_sc_hd__o21ai_1 _07502_ (.A1(_01536_),
    .A2(_01540_),
    .B1(_01544_),
    .Y(_01547_));
 sky130_fd_sc_hd__nand3_1 _07503_ (.A(_01547_),
    .B(_01531_),
    .C(_01533_),
    .Y(_01548_));
 sky130_fd_sc_hd__a21boi_1 _07504_ (.A1(_01528_),
    .A2(_01546_),
    .B1_N(_01548_),
    .Y(_01549_));
 sky130_fd_sc_hd__nand2_1 _07505_ (.A(_01522_),
    .B(_01549_),
    .Y(_01550_));
 sky130_fd_sc_hd__inv_2 _07506_ (.A(_01469_),
    .Y(_01551_));
 sky130_fd_sc_hd__nand2_1 _07507_ (.A(_01461_),
    .B(_01551_),
    .Y(_01552_));
 sky130_fd_sc_hd__nand3_1 _07508_ (.A(_01459_),
    .B(_01460_),
    .C(_01469_),
    .Y(_01553_));
 sky130_fd_sc_hd__nand2_1 _07509_ (.A(_01552_),
    .B(_01553_),
    .Y(_01555_));
 sky130_fd_sc_hd__nand2_1 _07510_ (.A(_01555_),
    .B(_01481_),
    .Y(_01556_));
 sky130_fd_sc_hd__nand3b_1 _07511_ (.A_N(_01481_),
    .B(_01552_),
    .C(_01553_),
    .Y(_01557_));
 sky130_fd_sc_hd__nand2_1 _07512_ (.A(_01556_),
    .B(_01557_),
    .Y(_01558_));
 sky130_fd_sc_hd__inv_2 _07513_ (.A(_01558_),
    .Y(_01559_));
 sky130_fd_sc_hd__nor2_1 _07514_ (.A(_01549_),
    .B(_01522_),
    .Y(_01560_));
 sky130_fd_sc_hd__a21oi_2 _07515_ (.A1(_01550_),
    .A2(_01559_),
    .B1(_01560_),
    .Y(_01561_));
 sky130_fd_sc_hd__nand2_1 _07516_ (.A(_01514_),
    .B(_01561_),
    .Y(_01562_));
 sky130_fd_sc_hd__nor2_1 _07517_ (.A(_01561_),
    .B(_01514_),
    .Y(_01563_));
 sky130_fd_sc_hd__a21o_1 _07518_ (.A1(_01506_),
    .A2(_01562_),
    .B1(_01563_),
    .X(_01564_));
 sky130_fd_sc_hd__nand2_1 _07519_ (.A(_01457_),
    .B(_01564_),
    .Y(_01566_));
 sky130_fd_sc_hd__nand2_1 _07520_ (.A(_01504_),
    .B(_01492_),
    .Y(_01567_));
 sky130_fd_sc_hd__a21oi_1 _07521_ (.A1(_01506_),
    .A2(_01562_),
    .B1(_01563_),
    .Y(_01568_));
 sky130_fd_sc_hd__nand2_1 _07522_ (.A(_01568_),
    .B(_01456_),
    .Y(_01569_));
 sky130_fd_sc_hd__nand3_1 _07523_ (.A(_01566_),
    .B(_01567_),
    .C(_01569_),
    .Y(_01570_));
 sky130_fd_sc_hd__nand2_1 _07524_ (.A(_01570_),
    .B(_01566_),
    .Y(_01571_));
 sky130_fd_sc_hd__inv_2 _07525_ (.A(_01415_),
    .Y(_01572_));
 sky130_fd_sc_hd__nand3_1 _07526_ (.A(_01572_),
    .B(_01414_),
    .C(_01408_),
    .Y(_01573_));
 sky130_fd_sc_hd__nand2_1 _07527_ (.A(_01572_),
    .B(_01408_),
    .Y(_01574_));
 sky130_fd_sc_hd__nand2_1 _07528_ (.A(_01446_),
    .B(_01413_),
    .Y(_01575_));
 sky130_fd_sc_hd__nand2_1 _07529_ (.A(_01574_),
    .B(_01575_),
    .Y(_01577_));
 sky130_fd_sc_hd__nand3_2 _07530_ (.A(_01571_),
    .B(_01573_),
    .C(_01577_),
    .Y(_01578_));
 sky130_fd_sc_hd__nand2_1 _07531_ (.A(_01448_),
    .B(_01578_),
    .Y(_01579_));
 sky130_fd_sc_hd__inv_2 _07532_ (.A(_01561_),
    .Y(_01580_));
 sky130_fd_sc_hd__nand2_1 _07533_ (.A(_01514_),
    .B(_01580_),
    .Y(_01581_));
 sky130_fd_sc_hd__nand3_1 _07534_ (.A(_01561_),
    .B(_01512_),
    .C(_01513_),
    .Y(_01582_));
 sky130_fd_sc_hd__nand2_1 _07535_ (.A(_01581_),
    .B(_01582_),
    .Y(_01583_));
 sky130_fd_sc_hd__nand2_1 _07536_ (.A(_01583_),
    .B(_01506_),
    .Y(_01584_));
 sky130_fd_sc_hd__nand3_1 _07537_ (.A(_01581_),
    .B(_01582_),
    .C(_01505_),
    .Y(_01585_));
 sky130_fd_sc_hd__nand2_1 _07538_ (.A(_01584_),
    .B(_01585_),
    .Y(_01586_));
 sky130_fd_sc_hd__nand3_1 _07539_ (.A(_01549_),
    .B(_01519_),
    .C(_01520_),
    .Y(_01588_));
 sky130_fd_sc_hd__nand3_1 _07540_ (.A(_01546_),
    .B(_01548_),
    .C(_01528_),
    .Y(_01589_));
 sky130_fd_sc_hd__nand2_1 _07541_ (.A(_01589_),
    .B(_01548_),
    .Y(_01590_));
 sky130_fd_sc_hd__nand2_1 _07542_ (.A(_01522_),
    .B(_01590_),
    .Y(_01591_));
 sky130_fd_sc_hd__nand2_1 _07543_ (.A(_01588_),
    .B(_01591_),
    .Y(_01592_));
 sky130_fd_sc_hd__nand2_1 _07544_ (.A(_01592_),
    .B(_01559_),
    .Y(_01593_));
 sky130_fd_sc_hd__nand3_1 _07545_ (.A(_01588_),
    .B(_01591_),
    .C(_01558_),
    .Y(_01594_));
 sky130_fd_sc_hd__nand2_1 _07546_ (.A(_01593_),
    .B(_01594_),
    .Y(_01595_));
 sky130_fd_sc_hd__inv_2 _07547_ (.A(_03226_),
    .Y(_01596_));
 sky130_fd_sc_hd__clkinv_4 _07548_ (.A(_00795_),
    .Y(_01597_));
 sky130_fd_sc_hd__nand2_1 _07549_ (.A(_03314_),
    .B(net44),
    .Y(_01599_));
 sky130_fd_sc_hd__o21ai_2 _07550_ (.A1(_01596_),
    .A2(_01597_),
    .B1(_01599_),
    .Y(_01600_));
 sky130_fd_sc_hd__nand2_1 _07551_ (.A(_04928_),
    .B(net55),
    .Y(_01601_));
 sky130_fd_sc_hd__inv_2 _07552_ (.A(_01601_),
    .Y(_01602_));
 sky130_fd_sc_hd__inv_2 _07553_ (.A(_01599_),
    .Y(_01603_));
 sky130_fd_sc_hd__nand3_1 _07554_ (.A(_01603_),
    .B(_05031_),
    .C(_00795_),
    .Y(_01604_));
 sky130_fd_sc_hd__a21boi_1 _07555_ (.A1(_01600_),
    .A2(_01602_),
    .B1_N(_01604_),
    .Y(_01605_));
 sky130_fd_sc_hd__nand3_1 _07556_ (.A(_01544_),
    .B(_01539_),
    .C(_01536_),
    .Y(_01606_));
 sky130_fd_sc_hd__a21o_1 _07557_ (.A1(_01544_),
    .A2(_01539_),
    .B1(_01536_),
    .X(_01607_));
 sky130_fd_sc_hd__nand3_2 _07558_ (.A(_01605_),
    .B(_01606_),
    .C(_01607_),
    .Y(_01608_));
 sky130_fd_sc_hd__nand2_1 _07559_ (.A(_00254_),
    .B(_01565_),
    .Y(_01610_));
 sky130_fd_sc_hd__nand2_1 _07560_ (.A(_00656_),
    .B(_04260_),
    .Y(_01611_));
 sky130_fd_sc_hd__nand2_1 _07561_ (.A(_04928_),
    .B(_04293_),
    .Y(_01612_));
 sky130_fd_sc_hd__nor2_1 _07562_ (.A(_01611_),
    .B(_01612_),
    .Y(_01613_));
 sky130_fd_sc_hd__nand2_1 _07563_ (.A(_01611_),
    .B(_01612_),
    .Y(_01614_));
 sky130_fd_sc_hd__nand2b_1 _07564_ (.A_N(_01613_),
    .B(_01614_),
    .Y(_01615_));
 sky130_fd_sc_hd__xor2_1 _07565_ (.A(_01610_),
    .B(_01615_),
    .X(_01616_));
 sky130_fd_sc_hd__nand2_1 _07566_ (.A(_01607_),
    .B(_01606_),
    .Y(_01617_));
 sky130_fd_sc_hd__nand3_1 _07567_ (.A(_01604_),
    .B(_01600_),
    .C(_01602_),
    .Y(_01618_));
 sky130_fd_sc_hd__nand2_1 _07568_ (.A(_01618_),
    .B(_01604_),
    .Y(_01619_));
 sky130_fd_sc_hd__nand2_2 _07569_ (.A(_01617_),
    .B(_01619_),
    .Y(_01621_));
 sky130_fd_sc_hd__a21boi_1 _07570_ (.A1(_01608_),
    .A2(_01616_),
    .B1_N(_01621_),
    .Y(_01622_));
 sky130_fd_sc_hd__nand2_1 _07571_ (.A(_01546_),
    .B(_01548_),
    .Y(_01623_));
 sky130_fd_sc_hd__nand2_1 _07572_ (.A(_01623_),
    .B(_01527_),
    .Y(_01624_));
 sky130_fd_sc_hd__nand2_2 _07573_ (.A(_01624_),
    .B(_01589_),
    .Y(_01625_));
 sky130_fd_sc_hd__nand2_1 _07574_ (.A(_01622_),
    .B(_01625_),
    .Y(_01626_));
 sky130_fd_sc_hd__a21o_1 _07575_ (.A1(_01475_),
    .A2(_01479_),
    .B1(_01478_),
    .X(_01627_));
 sky130_fd_sc_hd__nand2_1 _07576_ (.A(_01627_),
    .B(_01480_),
    .Y(_01628_));
 sky130_fd_sc_hd__inv_2 _07577_ (.A(_01610_),
    .Y(_01629_));
 sky130_fd_sc_hd__a21oi_1 _07578_ (.A1(_01614_),
    .A2(_01629_),
    .B1(_01613_),
    .Y(_01630_));
 sky130_fd_sc_hd__nand2_1 _07579_ (.A(_01628_),
    .B(_01630_),
    .Y(_01632_));
 sky130_fd_sc_hd__nand3b_1 _07580_ (.A_N(_01630_),
    .B(_01627_),
    .C(_01480_),
    .Y(_01633_));
 sky130_fd_sc_hd__nand2_1 _07581_ (.A(_01632_),
    .B(_01633_),
    .Y(_01634_));
 sky130_fd_sc_hd__nand2_1 _07582_ (.A(_04991_),
    .B(_00003_),
    .Y(_01635_));
 sky130_fd_sc_hd__nand2_1 _07583_ (.A(_04827_),
    .B(_01774_),
    .Y(_01636_));
 sky130_fd_sc_hd__nand2_1 _07584_ (.A(_00522_),
    .B(_00204_),
    .Y(_01637_));
 sky130_fd_sc_hd__or2_1 _07585_ (.A(_01636_),
    .B(_01637_),
    .X(_01638_));
 sky130_fd_sc_hd__nand2_1 _07586_ (.A(_01636_),
    .B(_01637_),
    .Y(_01639_));
 sky130_fd_sc_hd__nand2_1 _07587_ (.A(_01638_),
    .B(_01639_),
    .Y(_01640_));
 sky130_fd_sc_hd__or2_1 _07588_ (.A(_01635_),
    .B(_01640_),
    .X(_01641_));
 sky130_fd_sc_hd__nand2_1 _07589_ (.A(_01641_),
    .B(_01638_),
    .Y(_01643_));
 sky130_fd_sc_hd__inv_2 _07590_ (.A(_01643_),
    .Y(_01644_));
 sky130_fd_sc_hd__nand2_1 _07591_ (.A(_01634_),
    .B(_01644_),
    .Y(_01645_));
 sky130_fd_sc_hd__nand3_1 _07592_ (.A(_01643_),
    .B(_01632_),
    .C(_01633_),
    .Y(_01646_));
 sky130_fd_sc_hd__nand2_1 _07593_ (.A(_01645_),
    .B(_01646_),
    .Y(_01647_));
 sky130_fd_sc_hd__inv_2 _07594_ (.A(_01647_),
    .Y(_01648_));
 sky130_fd_sc_hd__nor2_1 _07595_ (.A(_01625_),
    .B(_01622_),
    .Y(_01649_));
 sky130_fd_sc_hd__a21oi_1 _07596_ (.A1(_01626_),
    .A2(_01648_),
    .B1(_01649_),
    .Y(_01650_));
 sky130_fd_sc_hd__nand2_1 _07597_ (.A(_01595_),
    .B(_01650_),
    .Y(_01651_));
 sky130_fd_sc_hd__nand2_1 _07598_ (.A(_01500_),
    .B(_01497_),
    .Y(_01652_));
 sky130_fd_sc_hd__nand2_1 _07599_ (.A(_01502_),
    .B(_01652_),
    .Y(_01654_));
 sky130_fd_sc_hd__and2_1 _07600_ (.A(_01646_),
    .B(_01633_),
    .X(_01655_));
 sky130_fd_sc_hd__nor2_1 _07601_ (.A(_01654_),
    .B(_01655_),
    .Y(_01656_));
 sky130_fd_sc_hd__nand2_1 _07602_ (.A(_01655_),
    .B(_01654_),
    .Y(_01657_));
 sky130_fd_sc_hd__nor2b_1 _07603_ (.A(_01656_),
    .B_N(_01657_),
    .Y(_01658_));
 sky130_fd_sc_hd__nor2_1 _07604_ (.A(_01650_),
    .B(_01595_),
    .Y(_01659_));
 sky130_fd_sc_hd__a21oi_1 _07605_ (.A1(_01651_),
    .A2(_01658_),
    .B1(_01659_),
    .Y(_01660_));
 sky130_fd_sc_hd__nand2_1 _07606_ (.A(_01586_),
    .B(_01660_),
    .Y(_01661_));
 sky130_fd_sc_hd__nor2_1 _07607_ (.A(_01660_),
    .B(_01586_),
    .Y(_01662_));
 sky130_fd_sc_hd__a21oi_1 _07608_ (.A1(_01661_),
    .A2(_01656_),
    .B1(_01662_),
    .Y(_01663_));
 sky130_fd_sc_hd__nand2_1 _07609_ (.A(_01457_),
    .B(_01568_),
    .Y(_01665_));
 sky130_fd_sc_hd__nand2_1 _07610_ (.A(_01564_),
    .B(_01456_),
    .Y(_01666_));
 sky130_fd_sc_hd__nand3b_1 _07611_ (.A_N(_01567_),
    .B(_01665_),
    .C(_01666_),
    .Y(_01667_));
 sky130_fd_sc_hd__nand2_1 _07612_ (.A(_01667_),
    .B(_01570_),
    .Y(_01668_));
 sky130_fd_sc_hd__nor2_1 _07613_ (.A(_01663_),
    .B(_01668_),
    .Y(_01669_));
 sky130_fd_sc_hd__nand2_1 _07614_ (.A(_01577_),
    .B(_01573_),
    .Y(_01670_));
 sky130_fd_sc_hd__a21boi_1 _07615_ (.A1(_01567_),
    .A2(_01569_),
    .B1_N(_01566_),
    .Y(_01671_));
 sky130_fd_sc_hd__nand2_1 _07616_ (.A(_01670_),
    .B(_01671_),
    .Y(_01672_));
 sky130_fd_sc_hd__nand3_2 _07617_ (.A(_01578_),
    .B(_01669_),
    .C(_01672_),
    .Y(_01673_));
 sky130_fd_sc_hd__inv_2 _07618_ (.A(_01673_),
    .Y(_01674_));
 sky130_fd_sc_hd__inv_2 _07619_ (.A(_01578_),
    .Y(_01676_));
 sky130_fd_sc_hd__nand3_2 _07620_ (.A(_01445_),
    .B(_01447_),
    .C(_01676_),
    .Y(_01677_));
 sky130_fd_sc_hd__nand3_2 _07621_ (.A(_01579_),
    .B(_01674_),
    .C(_01677_),
    .Y(_01678_));
 sky130_fd_sc_hd__inv_2 _07622_ (.A(_01678_),
    .Y(_01679_));
 sky130_fd_sc_hd__nand3_1 _07623_ (.A(_01131_),
    .B(_01006_),
    .C(_01007_),
    .Y(_01680_));
 sky130_fd_sc_hd__nand2_1 _07624_ (.A(_01424_),
    .B(_01423_),
    .Y(_01681_));
 sky130_fd_sc_hd__nand2_1 _07625_ (.A(_01008_),
    .B(_01681_),
    .Y(_01682_));
 sky130_fd_sc_hd__nand2_1 _07626_ (.A(_01680_),
    .B(_01682_),
    .Y(_01683_));
 sky130_fd_sc_hd__nand2_1 _07627_ (.A(_01683_),
    .B(_01137_),
    .Y(_01684_));
 sky130_fd_sc_hd__nand3b_1 _07628_ (.A_N(_01137_),
    .B(_01680_),
    .C(_01682_),
    .Y(_01685_));
 sky130_fd_sc_hd__nand2_1 _07629_ (.A(_01684_),
    .B(_01685_),
    .Y(_01687_));
 sky130_fd_sc_hd__nand2_1 _07630_ (.A(_01429_),
    .B(_01420_),
    .Y(_01688_));
 sky130_fd_sc_hd__nor2_1 _07631_ (.A(_01420_),
    .B(_01429_),
    .Y(_01689_));
 sky130_fd_sc_hd__a21oi_2 _07632_ (.A1(_01688_),
    .A2(_01437_),
    .B1(_01689_),
    .Y(_01690_));
 sky130_fd_sc_hd__inv_2 _07633_ (.A(_01690_),
    .Y(_01691_));
 sky130_fd_sc_hd__nand2_1 _07634_ (.A(_01687_),
    .B(_01691_),
    .Y(_01692_));
 sky130_fd_sc_hd__nand3_1 _07635_ (.A(_01690_),
    .B(_01684_),
    .C(_01685_),
    .Y(_01693_));
 sky130_fd_sc_hd__nand2_1 _07636_ (.A(_01692_),
    .B(_01693_),
    .Y(_01694_));
 sky130_fd_sc_hd__nor2_1 _07637_ (.A(_01435_),
    .B(_01436_),
    .Y(_01695_));
 sky130_fd_sc_hd__inv_2 _07638_ (.A(_01695_),
    .Y(_01696_));
 sky130_fd_sc_hd__nand2_1 _07639_ (.A(_01694_),
    .B(_01696_),
    .Y(_01698_));
 sky130_fd_sc_hd__nand3_1 _07640_ (.A(_01692_),
    .B(_01693_),
    .C(_01695_),
    .Y(_01699_));
 sky130_fd_sc_hd__nand2_1 _07641_ (.A(_01698_),
    .B(_01699_),
    .Y(_01700_));
 sky130_fd_sc_hd__nand2_1 _07642_ (.A(_01440_),
    .B(_01416_),
    .Y(_01701_));
 sky130_fd_sc_hd__nor2_1 _07643_ (.A(_01416_),
    .B(_01440_),
    .Y(_01702_));
 sky130_fd_sc_hd__a21o_1 _07644_ (.A1(_01701_),
    .A2(_01412_),
    .B1(_01702_),
    .X(_01703_));
 sky130_fd_sc_hd__nand2_2 _07645_ (.A(_01700_),
    .B(_01703_),
    .Y(_01704_));
 sky130_fd_sc_hd__a21oi_1 _07646_ (.A1(_01701_),
    .A2(_01412_),
    .B1(_01702_),
    .Y(_01705_));
 sky130_fd_sc_hd__nand3_1 _07647_ (.A(_01705_),
    .B(_01698_),
    .C(_01699_),
    .Y(_01706_));
 sky130_fd_sc_hd__nand2_1 _07648_ (.A(_01704_),
    .B(_01706_),
    .Y(_01707_));
 sky130_fd_sc_hd__nand2_1 _07649_ (.A(_01707_),
    .B(_01677_),
    .Y(_01709_));
 sky130_fd_sc_hd__inv_2 _07650_ (.A(_01677_),
    .Y(_01710_));
 sky130_fd_sc_hd__nand3_2 _07651_ (.A(_01710_),
    .B(_01704_),
    .C(_01706_),
    .Y(_01711_));
 sky130_fd_sc_hd__nand3_1 _07652_ (.A(_01679_),
    .B(_01709_),
    .C(_01711_),
    .Y(_01712_));
 sky130_fd_sc_hd__inv_2 _07653_ (.A(_01711_),
    .Y(_01713_));
 sky130_fd_sc_hd__nand2_1 _07654_ (.A(_01687_),
    .B(_01690_),
    .Y(_01714_));
 sky130_fd_sc_hd__nor2_1 _07655_ (.A(_01690_),
    .B(_01687_),
    .Y(_01715_));
 sky130_fd_sc_hd__a21o_1 _07656_ (.A1(_01714_),
    .A2(_01695_),
    .B1(_01715_),
    .X(_01716_));
 sky130_fd_sc_hd__inv_2 _07657_ (.A(_01139_),
    .Y(_01717_));
 sky130_fd_sc_hd__nand2_1 _07658_ (.A(_01000_),
    .B(_01717_),
    .Y(_01718_));
 sky130_fd_sc_hd__nand3_1 _07659_ (.A(_01139_),
    .B(_00998_),
    .C(_00999_),
    .Y(_01720_));
 sky130_fd_sc_hd__nand2_1 _07660_ (.A(_01718_),
    .B(_01720_),
    .Y(_01721_));
 sky130_fd_sc_hd__inv_2 _07661_ (.A(_01141_),
    .Y(_01722_));
 sky130_fd_sc_hd__nand2_1 _07662_ (.A(_01721_),
    .B(_01722_),
    .Y(_01723_));
 sky130_fd_sc_hd__nand3_1 _07663_ (.A(_01718_),
    .B(_01720_),
    .C(_01141_),
    .Y(_01724_));
 sky130_fd_sc_hd__nand2_1 _07664_ (.A(_01723_),
    .B(_01724_),
    .Y(_01725_));
 sky130_fd_sc_hd__nand2_1 _07665_ (.A(_01716_),
    .B(_01725_),
    .Y(_01726_));
 sky130_fd_sc_hd__nand2_1 _07666_ (.A(_01721_),
    .B(_01141_),
    .Y(_01727_));
 sky130_fd_sc_hd__nand3_1 _07667_ (.A(_01718_),
    .B(_01720_),
    .C(_01722_),
    .Y(_01728_));
 sky130_fd_sc_hd__nand2_1 _07668_ (.A(_01727_),
    .B(_01728_),
    .Y(_01729_));
 sky130_fd_sc_hd__a21oi_1 _07669_ (.A1(_01714_),
    .A2(_01695_),
    .B1(_01715_),
    .Y(_01731_));
 sky130_fd_sc_hd__nand2_1 _07670_ (.A(_01729_),
    .B(_01731_),
    .Y(_01732_));
 sky130_fd_sc_hd__nand2_1 _07671_ (.A(_01726_),
    .B(_01732_),
    .Y(_01733_));
 sky130_fd_sc_hd__inv_2 _07672_ (.A(_01704_),
    .Y(_01734_));
 sky130_fd_sc_hd__nand2_1 _07673_ (.A(_01733_),
    .B(_01734_),
    .Y(_01735_));
 sky130_fd_sc_hd__nand3_1 _07674_ (.A(_01726_),
    .B(_01704_),
    .C(_01732_),
    .Y(_01736_));
 sky130_fd_sc_hd__nand2_1 _07675_ (.A(_01735_),
    .B(_01736_),
    .Y(_01737_));
 sky130_fd_sc_hd__nor2_1 _07676_ (.A(_01713_),
    .B(_01737_),
    .Y(_01738_));
 sky130_fd_sc_hd__nand2_1 _07677_ (.A(_01737_),
    .B(_01713_),
    .Y(_01739_));
 sky130_fd_sc_hd__o21ai_1 _07678_ (.A1(_01712_),
    .A2(_01738_),
    .B1(_01739_),
    .Y(_01740_));
 sky130_fd_sc_hd__nand2_1 _07679_ (.A(_01148_),
    .B(_01150_),
    .Y(_01742_));
 sky130_fd_sc_hd__nand3_1 _07680_ (.A(_01145_),
    .B(_01146_),
    .C(_00986_),
    .Y(_01743_));
 sky130_fd_sc_hd__nand2_1 _07681_ (.A(_01742_),
    .B(_01743_),
    .Y(_01744_));
 sky130_fd_sc_hd__a21o_1 _07682_ (.A1(_01140_),
    .A2(_01141_),
    .B1(_01142_),
    .X(_01745_));
 sky130_fd_sc_hd__nand2_1 _07683_ (.A(_01744_),
    .B(_01745_),
    .Y(_01746_));
 sky130_fd_sc_hd__nand2_1 _07684_ (.A(_01152_),
    .B(_01143_),
    .Y(_01747_));
 sky130_fd_sc_hd__nand2_1 _07685_ (.A(_01746_),
    .B(_01747_),
    .Y(_01748_));
 sky130_fd_sc_hd__nor2_1 _07686_ (.A(_01726_),
    .B(_01748_),
    .Y(_01749_));
 sky130_fd_sc_hd__nand3_1 _07687_ (.A(_00990_),
    .B(_01746_),
    .C(_00991_),
    .Y(_01750_));
 sky130_fd_sc_hd__nand3_1 _07688_ (.A(_01749_),
    .B(_01154_),
    .C(_01750_),
    .Y(_01751_));
 sky130_fd_sc_hd__nand2_1 _07689_ (.A(_00992_),
    .B(_01746_),
    .Y(_01753_));
 sky130_fd_sc_hd__nand3_1 _07690_ (.A(_01153_),
    .B(_00990_),
    .C(_00991_),
    .Y(_01754_));
 sky130_fd_sc_hd__nor2_1 _07691_ (.A(_01731_),
    .B(_01729_),
    .Y(_01755_));
 sky130_fd_sc_hd__nand3_1 _07692_ (.A(_01755_),
    .B(_01746_),
    .C(_01747_),
    .Y(_01756_));
 sky130_fd_sc_hd__nand3_1 _07693_ (.A(_01753_),
    .B(_01754_),
    .C(_01756_),
    .Y(_01757_));
 sky130_fd_sc_hd__nand2_1 _07694_ (.A(_01751_),
    .B(_01757_),
    .Y(_01758_));
 sky130_fd_sc_hd__nand2_1 _07695_ (.A(_01748_),
    .B(_01726_),
    .Y(_01759_));
 sky130_fd_sc_hd__nand2_1 _07696_ (.A(_01759_),
    .B(_01756_),
    .Y(_01760_));
 sky130_fd_sc_hd__nor2_1 _07697_ (.A(_01704_),
    .B(_01733_),
    .Y(_01761_));
 sky130_fd_sc_hd__inv_2 _07698_ (.A(_01761_),
    .Y(_01762_));
 sky130_fd_sc_hd__nand2_1 _07699_ (.A(_01760_),
    .B(_01762_),
    .Y(_01764_));
 sky130_fd_sc_hd__nand3_1 _07700_ (.A(_01761_),
    .B(_01756_),
    .C(_01759_),
    .Y(_01765_));
 sky130_fd_sc_hd__nand2_1 _07701_ (.A(_01764_),
    .B(_01765_),
    .Y(_01766_));
 sky130_fd_sc_hd__nor2_1 _07702_ (.A(_01758_),
    .B(_01766_),
    .Y(_01767_));
 sky130_fd_sc_hd__inv_2 _07703_ (.A(_01757_),
    .Y(_01768_));
 sky130_fd_sc_hd__o21ai_1 _07704_ (.A1(_01765_),
    .A2(_01768_),
    .B1(_01751_),
    .Y(_01769_));
 sky130_fd_sc_hd__a21oi_1 _07705_ (.A1(_01740_),
    .A2(_01767_),
    .B1(_01769_),
    .Y(_01770_));
 sky130_fd_sc_hd__nand2_1 _07706_ (.A(_01159_),
    .B(_01161_),
    .Y(_01771_));
 sky130_fd_sc_hd__nand2_1 _07707_ (.A(_01771_),
    .B(_01154_),
    .Y(_01772_));
 sky130_fd_sc_hd__nand2_1 _07708_ (.A(_01772_),
    .B(_01162_),
    .Y(_01773_));
 sky130_fd_sc_hd__nand2_1 _07709_ (.A(_01164_),
    .B(_00793_),
    .Y(_01775_));
 sky130_fd_sc_hd__nand2_1 _07710_ (.A(_01775_),
    .B(_01159_),
    .Y(_01776_));
 sky130_fd_sc_hd__nand2_1 _07711_ (.A(_01167_),
    .B(_01776_),
    .Y(_01777_));
 sky130_fd_sc_hd__nor2_1 _07712_ (.A(_01773_),
    .B(_01777_),
    .Y(_01778_));
 sky130_fd_sc_hd__nand2_1 _07713_ (.A(_00799_),
    .B(_01778_),
    .Y(_01779_));
 sky130_fd_sc_hd__nor2_1 _07714_ (.A(_01770_),
    .B(_01779_),
    .Y(_01780_));
 sky130_fd_sc_hd__nor2_1 _07715_ (.A(_01173_),
    .B(_01780_),
    .Y(_01781_));
 sky130_fd_sc_hd__inv_2 _07716_ (.A(_01779_),
    .Y(_01782_));
 sky130_fd_sc_hd__nand3_1 _07717_ (.A(_01650_),
    .B(_01593_),
    .C(_01594_),
    .Y(_01783_));
 sky130_fd_sc_hd__a21o_1 _07718_ (.A1(_01626_),
    .A2(_01648_),
    .B1(_01649_),
    .X(_01784_));
 sky130_fd_sc_hd__nand2_1 _07719_ (.A(_01784_),
    .B(_01595_),
    .Y(_01786_));
 sky130_fd_sc_hd__nand2_1 _07720_ (.A(_01783_),
    .B(_01786_),
    .Y(_01787_));
 sky130_fd_sc_hd__nand2_1 _07721_ (.A(_01787_),
    .B(_01658_),
    .Y(_01788_));
 sky130_fd_sc_hd__nand3b_1 _07722_ (.A_N(_01658_),
    .B(_01783_),
    .C(_01786_),
    .Y(_01789_));
 sky130_fd_sc_hd__nand2_1 _07723_ (.A(_01788_),
    .B(_01789_),
    .Y(_01790_));
 sky130_fd_sc_hd__inv_2 _07724_ (.A(_01625_),
    .Y(_01791_));
 sky130_fd_sc_hd__nand2_1 _07725_ (.A(_01791_),
    .B(_01622_),
    .Y(_01792_));
 sky130_fd_sc_hd__nand3_1 _07726_ (.A(_01608_),
    .B(_01621_),
    .C(_01616_),
    .Y(_01793_));
 sky130_fd_sc_hd__nand2_1 _07727_ (.A(_01793_),
    .B(_01621_),
    .Y(_01794_));
 sky130_fd_sc_hd__nand2_1 _07728_ (.A(_01794_),
    .B(_01625_),
    .Y(_01795_));
 sky130_fd_sc_hd__nand2_1 _07729_ (.A(_01792_),
    .B(_01795_),
    .Y(_01797_));
 sky130_fd_sc_hd__nand2_1 _07730_ (.A(_01797_),
    .B(_01648_),
    .Y(_01798_));
 sky130_fd_sc_hd__nand3_1 _07731_ (.A(_01792_),
    .B(_01795_),
    .C(_01647_),
    .Y(_01799_));
 sky130_fd_sc_hd__nand2_1 _07732_ (.A(_01798_),
    .B(_01799_),
    .Y(_01800_));
 sky130_fd_sc_hd__nand2_1 _07733_ (.A(_01604_),
    .B(_01600_),
    .Y(_01801_));
 sky130_fd_sc_hd__nand2_1 _07734_ (.A(_01801_),
    .B(_01601_),
    .Y(_01802_));
 sky130_fd_sc_hd__nand2_1 _07735_ (.A(_01802_),
    .B(_01618_),
    .Y(_01803_));
 sky130_fd_sc_hd__nand2_1 _07736_ (.A(_03402_),
    .B(net44),
    .Y(_01804_));
 sky130_fd_sc_hd__nand2_1 _07737_ (.A(_03314_),
    .B(net33),
    .Y(_01805_));
 sky130_fd_sc_hd__nand2_1 _07738_ (.A(_01804_),
    .B(_01805_),
    .Y(_01806_));
 sky130_fd_sc_hd__nand2_1 _07739_ (.A(_03820_),
    .B(net55),
    .Y(_01808_));
 sky130_fd_sc_hd__inv_2 _07740_ (.A(_01808_),
    .Y(_01809_));
 sky130_fd_sc_hd__nor2_1 _07741_ (.A(_01804_),
    .B(_01805_),
    .Y(_01810_));
 sky130_fd_sc_hd__a21oi_1 _07742_ (.A1(_01806_),
    .A2(_01809_),
    .B1(_01810_),
    .Y(_01811_));
 sky130_fd_sc_hd__nand2_1 _07743_ (.A(_01803_),
    .B(_01811_),
    .Y(_01812_));
 sky130_fd_sc_hd__nand3b_1 _07744_ (.A_N(_01811_),
    .B(_01802_),
    .C(_01618_),
    .Y(_01813_));
 sky130_fd_sc_hd__nand2_1 _07745_ (.A(_04809_),
    .B(_01048_),
    .Y(_01814_));
 sky130_fd_sc_hd__nand2_1 _07746_ (.A(_03820_),
    .B(_01092_),
    .Y(_01815_));
 sky130_fd_sc_hd__nor2_1 _07747_ (.A(_01814_),
    .B(_01815_),
    .Y(_01816_));
 sky130_fd_sc_hd__inv_2 _07748_ (.A(_01816_),
    .Y(_01817_));
 sky130_fd_sc_hd__nand2_1 _07749_ (.A(_01814_),
    .B(_01815_),
    .Y(_01819_));
 sky130_fd_sc_hd__nand2_1 _07750_ (.A(_01817_),
    .B(_01819_),
    .Y(_01820_));
 sky130_fd_sc_hd__nand2_1 _07751_ (.A(_04819_),
    .B(_01158_),
    .Y(_01821_));
 sky130_fd_sc_hd__nand2_1 _07752_ (.A(_01820_),
    .B(_01821_),
    .Y(_01822_));
 sky130_fd_sc_hd__inv_2 _07753_ (.A(_01821_),
    .Y(_01823_));
 sky130_fd_sc_hd__nand3_1 _07754_ (.A(_01817_),
    .B(_01823_),
    .C(_01819_),
    .Y(_01824_));
 sky130_fd_sc_hd__nand2_1 _07755_ (.A(_01822_),
    .B(_01824_),
    .Y(_01825_));
 sky130_fd_sc_hd__inv_2 _07756_ (.A(_01825_),
    .Y(_01826_));
 sky130_fd_sc_hd__nand3_1 _07757_ (.A(_01812_),
    .B(_01813_),
    .C(_01826_),
    .Y(_01827_));
 sky130_fd_sc_hd__nand2_1 _07758_ (.A(_01827_),
    .B(_01813_),
    .Y(_01828_));
 sky130_fd_sc_hd__inv_2 _07759_ (.A(_01828_),
    .Y(_01830_));
 sky130_fd_sc_hd__nand2_1 _07760_ (.A(_01608_),
    .B(_01621_),
    .Y(_01831_));
 sky130_fd_sc_hd__xor2_1 _07761_ (.A(_01629_),
    .B(_01615_),
    .X(_01832_));
 sky130_fd_sc_hd__nand2_1 _07762_ (.A(_01831_),
    .B(_01832_),
    .Y(_01833_));
 sky130_fd_sc_hd__nand2_1 _07763_ (.A(_01833_),
    .B(_01793_),
    .Y(_01834_));
 sky130_fd_sc_hd__nand2_1 _07764_ (.A(_01830_),
    .B(_01834_),
    .Y(_01835_));
 sky130_fd_sc_hd__nand2_1 _07765_ (.A(_01640_),
    .B(_01635_),
    .Y(_01836_));
 sky130_fd_sc_hd__nand2_1 _07766_ (.A(_01641_),
    .B(_01836_),
    .Y(_01837_));
 sky130_fd_sc_hd__nand2_1 _07767_ (.A(_01824_),
    .B(_01817_),
    .Y(_01838_));
 sky130_fd_sc_hd__inv_2 _07768_ (.A(_01838_),
    .Y(_01839_));
 sky130_fd_sc_hd__nand2_1 _07769_ (.A(_01837_),
    .B(_01839_),
    .Y(_01841_));
 sky130_fd_sc_hd__nand3_2 _07770_ (.A(_01641_),
    .B(_01838_),
    .C(_01836_),
    .Y(_01842_));
 sky130_fd_sc_hd__nand2_1 _07771_ (.A(_01841_),
    .B(_01842_),
    .Y(_01843_));
 sky130_fd_sc_hd__nand2_1 _07772_ (.A(_04895_),
    .B(_00003_),
    .Y(_01844_));
 sky130_fd_sc_hd__nand2_1 _07773_ (.A(_04911_),
    .B(_00412_),
    .Y(_01845_));
 sky130_fd_sc_hd__nand2_1 _07774_ (.A(_04827_),
    .B(_00204_),
    .Y(_01846_));
 sky130_fd_sc_hd__or2_1 _07775_ (.A(_01845_),
    .B(_01846_),
    .X(_01847_));
 sky130_fd_sc_hd__nand2_1 _07776_ (.A(_01845_),
    .B(_01846_),
    .Y(_01848_));
 sky130_fd_sc_hd__nand2_1 _07777_ (.A(_01847_),
    .B(_01848_),
    .Y(_01849_));
 sky130_fd_sc_hd__or2_1 _07778_ (.A(_01844_),
    .B(_01849_),
    .X(_01850_));
 sky130_fd_sc_hd__nand2_1 _07779_ (.A(_01850_),
    .B(_01847_),
    .Y(_01852_));
 sky130_fd_sc_hd__nand2_1 _07780_ (.A(_01843_),
    .B(_01852_),
    .Y(_01853_));
 sky130_fd_sc_hd__inv_2 _07781_ (.A(_01852_),
    .Y(_01854_));
 sky130_fd_sc_hd__nand3_1 _07782_ (.A(_01841_),
    .B(_01854_),
    .C(_01842_),
    .Y(_01855_));
 sky130_fd_sc_hd__nand2_1 _07783_ (.A(_01853_),
    .B(_01855_),
    .Y(_01856_));
 sky130_fd_sc_hd__nor2_1 _07784_ (.A(_01834_),
    .B(_01830_),
    .Y(_01857_));
 sky130_fd_sc_hd__a21oi_1 _07785_ (.A1(_01835_),
    .A2(_01856_),
    .B1(_01857_),
    .Y(_01858_));
 sky130_fd_sc_hd__nand2_1 _07786_ (.A(_01800_),
    .B(_01858_),
    .Y(_01859_));
 sky130_fd_sc_hd__a22o_1 _07787_ (.A1(_04991_),
    .A2(_05032_),
    .B1(_04992_),
    .B2(_05029_),
    .X(_01860_));
 sky130_fd_sc_hd__nand2_1 _07788_ (.A(_01497_),
    .B(_01860_),
    .Y(_01861_));
 sky130_fd_sc_hd__nand3_1 _07789_ (.A(_01841_),
    .B(_01842_),
    .C(_01852_),
    .Y(_01863_));
 sky130_fd_sc_hd__and2_1 _07790_ (.A(_01863_),
    .B(_01842_),
    .X(_01864_));
 sky130_fd_sc_hd__nor2_2 _07791_ (.A(_01861_),
    .B(_01864_),
    .Y(_01865_));
 sky130_fd_sc_hd__nand2_1 _07792_ (.A(_01864_),
    .B(_01861_),
    .Y(_01866_));
 sky130_fd_sc_hd__nor2b_1 _07793_ (.A(_01865_),
    .B_N(_01866_),
    .Y(_01867_));
 sky130_fd_sc_hd__nor2_1 _07794_ (.A(_01858_),
    .B(_01800_),
    .Y(_01868_));
 sky130_fd_sc_hd__a21oi_2 _07795_ (.A1(_01859_),
    .A2(_01867_),
    .B1(_01868_),
    .Y(_01869_));
 sky130_fd_sc_hd__nand2_1 _07796_ (.A(_01790_),
    .B(_01869_),
    .Y(_01870_));
 sky130_fd_sc_hd__nor2_1 _07797_ (.A(_01869_),
    .B(_01790_),
    .Y(_01871_));
 sky130_fd_sc_hd__a21o_1 _07798_ (.A1(_01870_),
    .A2(_01865_),
    .B1(_01871_),
    .X(_01872_));
 sky130_fd_sc_hd__nand3_1 _07799_ (.A(_01660_),
    .B(_01584_),
    .C(_01585_),
    .Y(_01874_));
 sky130_fd_sc_hd__a21o_1 _07800_ (.A1(_01651_),
    .A2(_01658_),
    .B1(_01659_),
    .X(_01875_));
 sky130_fd_sc_hd__nand2_1 _07801_ (.A(_01586_),
    .B(_01875_),
    .Y(_01876_));
 sky130_fd_sc_hd__nand2_1 _07802_ (.A(_01874_),
    .B(_01876_),
    .Y(_01877_));
 sky130_fd_sc_hd__nand2_1 _07803_ (.A(_01877_),
    .B(_01656_),
    .Y(_01878_));
 sky130_fd_sc_hd__nand3b_1 _07804_ (.A_N(_01656_),
    .B(_01874_),
    .C(_01876_),
    .Y(_01879_));
 sky130_fd_sc_hd__nand3_2 _07805_ (.A(_01872_),
    .B(_01878_),
    .C(_01879_),
    .Y(_01880_));
 sky130_fd_sc_hd__nand2_1 _07806_ (.A(_01843_),
    .B(_01854_),
    .Y(_01881_));
 sky130_fd_sc_hd__nand2_1 _07807_ (.A(_01881_),
    .B(_01863_),
    .Y(_01882_));
 sky130_fd_sc_hd__nand2_1 _07808_ (.A(_01831_),
    .B(_01616_),
    .Y(_01883_));
 sky130_fd_sc_hd__nand3_1 _07809_ (.A(_01608_),
    .B(_01621_),
    .C(_01832_),
    .Y(_01885_));
 sky130_fd_sc_hd__nand2_1 _07810_ (.A(_01883_),
    .B(_01885_),
    .Y(_01886_));
 sky130_fd_sc_hd__nor2_1 _07811_ (.A(_01828_),
    .B(_01886_),
    .Y(_01887_));
 sky130_fd_sc_hd__nand2_1 _07812_ (.A(_01886_),
    .B(_01828_),
    .Y(_01888_));
 sky130_fd_sc_hd__o21ai_1 _07813_ (.A1(_01882_),
    .A2(_01887_),
    .B1(_01888_),
    .Y(_01889_));
 sky130_fd_sc_hd__nand3_1 _07814_ (.A(_01889_),
    .B(_01798_),
    .C(_01799_),
    .Y(_01890_));
 sky130_fd_sc_hd__nand3_1 _07815_ (.A(_01890_),
    .B(_01867_),
    .C(_01859_),
    .Y(_01891_));
 sky130_fd_sc_hd__nand3_1 _07816_ (.A(_01858_),
    .B(_01798_),
    .C(_01799_),
    .Y(_01892_));
 sky130_fd_sc_hd__nand2_1 _07817_ (.A(_01800_),
    .B(_01889_),
    .Y(_01893_));
 sky130_fd_sc_hd__nand2b_1 _07818_ (.A_N(_01865_),
    .B(_01866_),
    .Y(_01894_));
 sky130_fd_sc_hd__nand3_1 _07819_ (.A(_01892_),
    .B(_01893_),
    .C(_01894_),
    .Y(_01896_));
 sky130_fd_sc_hd__nand2_1 _07820_ (.A(_01891_),
    .B(_01896_),
    .Y(_01897_));
 sky130_fd_sc_hd__nand2_1 _07821_ (.A(_01812_),
    .B(_01813_),
    .Y(_01898_));
 sky130_fd_sc_hd__nand2_1 _07822_ (.A(_01898_),
    .B(_01825_),
    .Y(_01899_));
 sky130_fd_sc_hd__nand2_1 _07823_ (.A(_01899_),
    .B(_01827_),
    .Y(_01900_));
 sky130_fd_sc_hd__nand2b_1 _07824_ (.A_N(_01810_),
    .B(_01806_),
    .Y(_01901_));
 sky130_fd_sc_hd__or2b_1 _07825_ (.A(_01901_),
    .B_N(_01808_),
    .X(_01902_));
 sky130_fd_sc_hd__nand2_1 _07826_ (.A(_01901_),
    .B(_01809_),
    .Y(_01903_));
 sky130_fd_sc_hd__nand2_1 _07827_ (.A(_01902_),
    .B(_01903_),
    .Y(_01904_));
 sky130_fd_sc_hd__nand2_1 _07828_ (.A(_00656_),
    .B(_00751_),
    .Y(_01905_));
 sky130_fd_sc_hd__nand2_1 _07829_ (.A(_04928_),
    .B(_00795_),
    .Y(_01907_));
 sky130_fd_sc_hd__nand2_1 _07830_ (.A(_01905_),
    .B(_01907_),
    .Y(_01908_));
 sky130_fd_sc_hd__nand2_1 _07831_ (.A(_04809_),
    .B(_00861_),
    .Y(_01909_));
 sky130_fd_sc_hd__inv_2 _07832_ (.A(_01909_),
    .Y(_01910_));
 sky130_fd_sc_hd__nor2_1 _07833_ (.A(_01905_),
    .B(_01907_),
    .Y(_01911_));
 sky130_fd_sc_hd__a21oi_1 _07834_ (.A1(_01908_),
    .A2(_01910_),
    .B1(_01911_),
    .Y(_01912_));
 sky130_fd_sc_hd__inv_2 _07835_ (.A(_01912_),
    .Y(_01913_));
 sky130_fd_sc_hd__nand2_1 _07836_ (.A(_01904_),
    .B(_01913_),
    .Y(_01914_));
 sky130_fd_sc_hd__nand2_1 _07837_ (.A(_04827_),
    .B(_01565_),
    .Y(_01915_));
 sky130_fd_sc_hd__nand2_1 _07838_ (.A(_04819_),
    .B(_01048_),
    .Y(_01916_));
 sky130_fd_sc_hd__nand2_1 _07839_ (.A(_00254_),
    .B(_01092_),
    .Y(_01918_));
 sky130_fd_sc_hd__nor2_1 _07840_ (.A(_01916_),
    .B(_01918_),
    .Y(_01919_));
 sky130_fd_sc_hd__nand2_1 _07841_ (.A(_01916_),
    .B(_01918_),
    .Y(_01920_));
 sky130_fd_sc_hd__nor2b_1 _07842_ (.A(_01919_),
    .B_N(_01920_),
    .Y(_01921_));
 sky130_fd_sc_hd__or2_1 _07843_ (.A(_01915_),
    .B(_01921_),
    .X(_01922_));
 sky130_fd_sc_hd__nand2_1 _07844_ (.A(_01921_),
    .B(_01915_),
    .Y(_01923_));
 sky130_fd_sc_hd__nand2_1 _07845_ (.A(_01922_),
    .B(_01923_),
    .Y(_01924_));
 sky130_fd_sc_hd__nand3_1 _07846_ (.A(_01902_),
    .B(_01912_),
    .C(_01903_),
    .Y(_01925_));
 sky130_fd_sc_hd__nand3_1 _07847_ (.A(_01914_),
    .B(_01924_),
    .C(_01925_),
    .Y(_01926_));
 sky130_fd_sc_hd__nand3_1 _07848_ (.A(_01900_),
    .B(_01926_),
    .C(_01914_),
    .Y(_01927_));
 sky130_fd_sc_hd__nand2_1 _07849_ (.A(_01849_),
    .B(_01844_),
    .Y(_01929_));
 sky130_fd_sc_hd__nand2_1 _07850_ (.A(_01850_),
    .B(_01929_),
    .Y(_01930_));
 sky130_fd_sc_hd__inv_2 _07851_ (.A(_01915_),
    .Y(_01931_));
 sky130_fd_sc_hd__a21oi_1 _07852_ (.A1(_01920_),
    .A2(_01931_),
    .B1(_01919_),
    .Y(_01932_));
 sky130_fd_sc_hd__nand2_1 _07853_ (.A(_01930_),
    .B(_01932_),
    .Y(_01933_));
 sky130_fd_sc_hd__inv_2 _07854_ (.A(_01932_),
    .Y(_01934_));
 sky130_fd_sc_hd__nand3_1 _07855_ (.A(_01850_),
    .B(_01929_),
    .C(_01934_),
    .Y(_01935_));
 sky130_fd_sc_hd__nand2_1 _07856_ (.A(_01933_),
    .B(_01935_),
    .Y(_01936_));
 sky130_fd_sc_hd__inv_2 _07857_ (.A(_01807_),
    .Y(_01937_));
 sky130_fd_sc_hd__nand2_1 _07858_ (.A(_04895_),
    .B(_00412_),
    .Y(_01938_));
 sky130_fd_sc_hd__nor3_1 _07859_ (.A(_00264_),
    .B(_01937_),
    .C(_01938_),
    .Y(_01940_));
 sky130_fd_sc_hd__nand2_1 _07860_ (.A(_01936_),
    .B(_01940_),
    .Y(_01941_));
 sky130_fd_sc_hd__inv_2 _07861_ (.A(_01940_),
    .Y(_01942_));
 sky130_fd_sc_hd__nand3_1 _07862_ (.A(_01933_),
    .B(_01942_),
    .C(_01935_),
    .Y(_01943_));
 sky130_fd_sc_hd__nand2_1 _07863_ (.A(_01941_),
    .B(_01943_),
    .Y(_01944_));
 sky130_fd_sc_hd__nand2_1 _07864_ (.A(_01926_),
    .B(_01914_),
    .Y(_01945_));
 sky130_fd_sc_hd__inv_2 _07865_ (.A(_01900_),
    .Y(_01946_));
 sky130_fd_sc_hd__nand2_2 _07866_ (.A(_01945_),
    .B(_01946_),
    .Y(_01947_));
 sky130_fd_sc_hd__inv_2 _07867_ (.A(_01947_),
    .Y(_01948_));
 sky130_fd_sc_hd__a21oi_1 _07868_ (.A1(_01927_),
    .A2(_01944_),
    .B1(_01948_),
    .Y(_01949_));
 sky130_fd_sc_hd__nand2_1 _07869_ (.A(_01835_),
    .B(_01888_),
    .Y(_01951_));
 sky130_fd_sc_hd__nand2_1 _07870_ (.A(_01951_),
    .B(_01882_),
    .Y(_01952_));
 sky130_fd_sc_hd__nand3_1 _07871_ (.A(_01835_),
    .B(_01888_),
    .C(_01856_),
    .Y(_01953_));
 sky130_fd_sc_hd__nand2_1 _07872_ (.A(_01952_),
    .B(_01953_),
    .Y(_01954_));
 sky130_fd_sc_hd__nand2_1 _07873_ (.A(_01949_),
    .B(_01954_),
    .Y(_01955_));
 sky130_fd_sc_hd__inv_2 _07874_ (.A(_04992_),
    .Y(_01956_));
 sky130_fd_sc_hd__clkinv_4 _07875_ (.A(_03028_),
    .Y(_01957_));
 sky130_fd_sc_hd__a21boi_1 _07876_ (.A1(_01933_),
    .A2(_01940_),
    .B1_N(_01935_),
    .Y(_01958_));
 sky130_fd_sc_hd__nor3_2 _07877_ (.A(_01956_),
    .B(_01957_),
    .C(_01958_),
    .Y(_01959_));
 sky130_fd_sc_hd__o21ai_1 _07878_ (.A1(_01956_),
    .A2(_01957_),
    .B1(_01958_),
    .Y(_01960_));
 sky130_fd_sc_hd__nor2b_1 _07879_ (.A(_01959_),
    .B_N(_01960_),
    .Y(_01962_));
 sky130_fd_sc_hd__nor2_1 _07880_ (.A(_01954_),
    .B(_01949_),
    .Y(_01963_));
 sky130_fd_sc_hd__a21oi_1 _07881_ (.A1(_01955_),
    .A2(_01962_),
    .B1(_01963_),
    .Y(_01964_));
 sky130_fd_sc_hd__nand2_1 _07882_ (.A(_01897_),
    .B(_01964_),
    .Y(_01965_));
 sky130_fd_sc_hd__nor2_1 _07883_ (.A(_01964_),
    .B(_01897_),
    .Y(_01966_));
 sky130_fd_sc_hd__a21oi_1 _07884_ (.A1(_01965_),
    .A2(_01959_),
    .B1(_01966_),
    .Y(_01967_));
 sky130_fd_sc_hd__inv_2 _07885_ (.A(_01869_),
    .Y(_01968_));
 sky130_fd_sc_hd__nand2_1 _07886_ (.A(_01968_),
    .B(_01790_),
    .Y(_01969_));
 sky130_fd_sc_hd__nand3_1 _07887_ (.A(_01869_),
    .B(_01788_),
    .C(_01789_),
    .Y(_01970_));
 sky130_fd_sc_hd__nand2_1 _07888_ (.A(_01969_),
    .B(_01970_),
    .Y(_01971_));
 sky130_fd_sc_hd__nand2_1 _07889_ (.A(_01971_),
    .B(_01865_),
    .Y(_01973_));
 sky130_fd_sc_hd__nand3b_1 _07890_ (.A_N(_01865_),
    .B(_01969_),
    .C(_01970_),
    .Y(_01974_));
 sky130_fd_sc_hd__nand2_1 _07891_ (.A(_01973_),
    .B(_01974_),
    .Y(_01975_));
 sky130_fd_sc_hd__nor2_1 _07892_ (.A(_01967_),
    .B(_01975_),
    .Y(_01976_));
 sky130_fd_sc_hd__nand2_1 _07893_ (.A(_01878_),
    .B(_01879_),
    .Y(_01977_));
 sky130_fd_sc_hd__a21oi_1 _07894_ (.A1(_01870_),
    .A2(_01865_),
    .B1(_01871_),
    .Y(_01978_));
 sky130_fd_sc_hd__nand2_1 _07895_ (.A(_01977_),
    .B(_01978_),
    .Y(_01979_));
 sky130_fd_sc_hd__nand3_2 _07896_ (.A(_01880_),
    .B(_01976_),
    .C(_01979_),
    .Y(_01980_));
 sky130_fd_sc_hd__a21o_1 _07897_ (.A1(_01661_),
    .A2(_01656_),
    .B1(_01662_),
    .X(_01981_));
 sky130_fd_sc_hd__nand3_1 _07898_ (.A(_01981_),
    .B(_01570_),
    .C(_01667_),
    .Y(_01982_));
 sky130_fd_sc_hd__nand2_1 _07899_ (.A(_01668_),
    .B(_01663_),
    .Y(_01984_));
 sky130_fd_sc_hd__nand2_1 _07900_ (.A(_01982_),
    .B(_01984_),
    .Y(_01985_));
 sky130_fd_sc_hd__nand2_1 _07901_ (.A(_01985_),
    .B(_01880_),
    .Y(_01986_));
 sky130_fd_sc_hd__nor2_1 _07902_ (.A(_01978_),
    .B(_01977_),
    .Y(_01987_));
 sky130_fd_sc_hd__nand3_1 _07903_ (.A(_01982_),
    .B(_01987_),
    .C(_01984_),
    .Y(_01988_));
 sky130_fd_sc_hd__nand2_1 _07904_ (.A(_01986_),
    .B(_01988_),
    .Y(_01989_));
 sky130_fd_sc_hd__nor2_1 _07905_ (.A(_01980_),
    .B(_01989_),
    .Y(_01990_));
 sky130_fd_sc_hd__nand2_1 _07906_ (.A(_01578_),
    .B(_01672_),
    .Y(_01991_));
 sky130_fd_sc_hd__nand2_1 _07907_ (.A(_01991_),
    .B(_01982_),
    .Y(_01992_));
 sky130_fd_sc_hd__nand2_1 _07908_ (.A(_01992_),
    .B(_01673_),
    .Y(_01993_));
 sky130_fd_sc_hd__nand2_1 _07909_ (.A(_01993_),
    .B(_01988_),
    .Y(_01995_));
 sky130_fd_sc_hd__nor2_1 _07910_ (.A(_01880_),
    .B(_01985_),
    .Y(_01996_));
 sky130_fd_sc_hd__nand3_2 _07911_ (.A(_01996_),
    .B(_01992_),
    .C(_01673_),
    .Y(_01997_));
 sky130_fd_sc_hd__nand3_1 _07912_ (.A(_01990_),
    .B(_01995_),
    .C(_01997_),
    .Y(_01998_));
 sky130_fd_sc_hd__nand2_1 _07913_ (.A(_01579_),
    .B(_01677_),
    .Y(_01999_));
 sky130_fd_sc_hd__nand2_1 _07914_ (.A(_01999_),
    .B(_01673_),
    .Y(_02000_));
 sky130_fd_sc_hd__nand2_1 _07915_ (.A(_02000_),
    .B(_01678_),
    .Y(_02001_));
 sky130_fd_sc_hd__nand2_1 _07916_ (.A(_02001_),
    .B(_01997_),
    .Y(_02002_));
 sky130_fd_sc_hd__inv_2 _07917_ (.A(_01997_),
    .Y(_02003_));
 sky130_fd_sc_hd__nand3_1 _07918_ (.A(_02000_),
    .B(_02003_),
    .C(_01678_),
    .Y(_02004_));
 sky130_fd_sc_hd__nand2_1 _07919_ (.A(_02002_),
    .B(_02004_),
    .Y(_02006_));
 sky130_fd_sc_hd__o21ai_1 _07920_ (.A1(_01998_),
    .A2(_02006_),
    .B1(_02004_),
    .Y(_02007_));
 sky130_fd_sc_hd__nand3_1 _07921_ (.A(_01964_),
    .B(_01891_),
    .C(_01896_),
    .Y(_02008_));
 sky130_fd_sc_hd__nand3_1 _07922_ (.A(_01947_),
    .B(_01927_),
    .C(_01944_),
    .Y(_02009_));
 sky130_fd_sc_hd__nand2_1 _07923_ (.A(_02009_),
    .B(_01947_),
    .Y(_02010_));
 sky130_fd_sc_hd__nand2_1 _07924_ (.A(_01951_),
    .B(_01856_),
    .Y(_02011_));
 sky130_fd_sc_hd__nand3_1 _07925_ (.A(_01835_),
    .B(_01888_),
    .C(_01882_),
    .Y(_02012_));
 sky130_fd_sc_hd__nand2_1 _07926_ (.A(_02011_),
    .B(_02012_),
    .Y(_02013_));
 sky130_fd_sc_hd__nand2_1 _07927_ (.A(_02010_),
    .B(_02013_),
    .Y(_02014_));
 sky130_fd_sc_hd__nand3_1 _07928_ (.A(_02014_),
    .B(_01955_),
    .C(_01962_),
    .Y(_02015_));
 sky130_fd_sc_hd__nand2_1 _07929_ (.A(_02015_),
    .B(_02014_),
    .Y(_02017_));
 sky130_fd_sc_hd__nand2_1 _07930_ (.A(_02017_),
    .B(_01897_),
    .Y(_02018_));
 sky130_fd_sc_hd__nand2_1 _07931_ (.A(_02008_),
    .B(_02018_),
    .Y(_02019_));
 sky130_fd_sc_hd__nand2_1 _07932_ (.A(_02019_),
    .B(_01959_),
    .Y(_02020_));
 sky130_fd_sc_hd__nand3b_1 _07933_ (.A_N(_01959_),
    .B(_02008_),
    .C(_02018_),
    .Y(_02021_));
 sky130_fd_sc_hd__nand2_1 _07934_ (.A(_02020_),
    .B(_02021_),
    .Y(_02022_));
 sky130_fd_sc_hd__nand2_1 _07935_ (.A(_01947_),
    .B(_01927_),
    .Y(_02023_));
 sky130_fd_sc_hd__nand3_1 _07936_ (.A(_02023_),
    .B(_01943_),
    .C(_01941_),
    .Y(_02024_));
 sky130_fd_sc_hd__nand2_1 _07937_ (.A(_02024_),
    .B(_02009_),
    .Y(_02025_));
 sky130_fd_sc_hd__nand2_1 _07938_ (.A(_01914_),
    .B(_01925_),
    .Y(_02026_));
 sky130_fd_sc_hd__inv_2 _07939_ (.A(_01924_),
    .Y(_02028_));
 sky130_fd_sc_hd__nand2_1 _07940_ (.A(_02026_),
    .B(_02028_),
    .Y(_02029_));
 sky130_fd_sc_hd__nand2_1 _07941_ (.A(_02029_),
    .B(_01926_),
    .Y(_02030_));
 sky130_fd_sc_hd__nand2b_1 _07942_ (.A_N(_01911_),
    .B(_01908_),
    .Y(_02031_));
 sky130_fd_sc_hd__or2_1 _07943_ (.A(_01909_),
    .B(_02031_),
    .X(_02032_));
 sky130_fd_sc_hd__nand2_1 _07944_ (.A(_02031_),
    .B(_01909_),
    .Y(_02033_));
 sky130_fd_sc_hd__nand2_1 _07945_ (.A(_02032_),
    .B(_02033_),
    .Y(_02034_));
 sky130_fd_sc_hd__nand2_1 _07946_ (.A(_00522_),
    .B(_01535_),
    .Y(_02035_));
 sky130_fd_sc_hd__nand2_1 _07947_ (.A(_00254_),
    .B(_00751_),
    .Y(_02036_));
 sky130_fd_sc_hd__nand2_1 _07948_ (.A(_00656_),
    .B(_02379_),
    .Y(_02037_));
 sky130_fd_sc_hd__or2_1 _07949_ (.A(_02036_),
    .B(_02037_),
    .X(_02039_));
 sky130_fd_sc_hd__nand2_1 _07950_ (.A(_02036_),
    .B(_02037_),
    .Y(_02040_));
 sky130_fd_sc_hd__nand2_1 _07951_ (.A(_02039_),
    .B(_02040_),
    .Y(_02041_));
 sky130_fd_sc_hd__o21ai_1 _07952_ (.A1(_02035_),
    .A2(_02041_),
    .B1(_02039_),
    .Y(_02042_));
 sky130_fd_sc_hd__inv_2 _07953_ (.A(_02042_),
    .Y(_02043_));
 sky130_fd_sc_hd__nand2_1 _07954_ (.A(_02034_),
    .B(_02043_),
    .Y(_02044_));
 sky130_fd_sc_hd__nand2_1 _07955_ (.A(_04827_),
    .B(_01048_),
    .Y(_02045_));
 sky130_fd_sc_hd__nand2_1 _07956_ (.A(_04819_),
    .B(_01092_),
    .Y(_02046_));
 sky130_fd_sc_hd__nor2_1 _07957_ (.A(_02045_),
    .B(_02046_),
    .Y(_02047_));
 sky130_fd_sc_hd__inv_2 _07958_ (.A(_02047_),
    .Y(_02048_));
 sky130_fd_sc_hd__nand2_1 _07959_ (.A(_02045_),
    .B(_02046_),
    .Y(_02050_));
 sky130_fd_sc_hd__nand2_1 _07960_ (.A(_04911_),
    .B(_01158_),
    .Y(_02051_));
 sky130_fd_sc_hd__inv_2 _07961_ (.A(_02051_),
    .Y(_02052_));
 sky130_fd_sc_hd__a21o_1 _07962_ (.A1(_02048_),
    .A2(_02050_),
    .B1(_02052_),
    .X(_02053_));
 sky130_fd_sc_hd__nand3_1 _07963_ (.A(_02048_),
    .B(_02052_),
    .C(_02050_),
    .Y(_02054_));
 sky130_fd_sc_hd__nand2_1 _07964_ (.A(_02053_),
    .B(_02054_),
    .Y(_02055_));
 sky130_fd_sc_hd__inv_2 _07965_ (.A(_02055_),
    .Y(_02056_));
 sky130_fd_sc_hd__nand3_1 _07966_ (.A(_02032_),
    .B(_02042_),
    .C(_02033_),
    .Y(_02057_));
 sky130_fd_sc_hd__a21boi_2 _07967_ (.A1(_02044_),
    .A2(_02056_),
    .B1_N(_02057_),
    .Y(_02058_));
 sky130_fd_sc_hd__nand2_1 _07968_ (.A(_02030_),
    .B(_02058_),
    .Y(_02059_));
 sky130_fd_sc_hd__o21ai_1 _07969_ (.A1(_00264_),
    .A2(_01937_),
    .B1(_01938_),
    .Y(_02061_));
 sky130_fd_sc_hd__nand2_1 _07970_ (.A(_01942_),
    .B(_02061_),
    .Y(_02062_));
 sky130_fd_sc_hd__and2_1 _07971_ (.A(_02054_),
    .B(_02048_),
    .X(_02063_));
 sky130_fd_sc_hd__nor2_1 _07972_ (.A(_02062_),
    .B(_02063_),
    .Y(_02064_));
 sky130_fd_sc_hd__inv_2 _07973_ (.A(_02064_),
    .Y(_02065_));
 sky130_fd_sc_hd__nand2_1 _07974_ (.A(_02063_),
    .B(_02062_),
    .Y(_02066_));
 sky130_fd_sc_hd__nand2_1 _07975_ (.A(_02065_),
    .B(_02066_),
    .Y(_02067_));
 sky130_fd_sc_hd__inv_2 _07976_ (.A(_02067_),
    .Y(_02068_));
 sky130_fd_sc_hd__nor2_1 _07977_ (.A(_02058_),
    .B(_02030_),
    .Y(_02069_));
 sky130_fd_sc_hd__a21oi_2 _07978_ (.A1(_02059_),
    .A2(_02068_),
    .B1(_02069_),
    .Y(_02070_));
 sky130_fd_sc_hd__nand2_1 _07979_ (.A(_02025_),
    .B(_02070_),
    .Y(_02072_));
 sky130_fd_sc_hd__nor2_1 _07980_ (.A(_02070_),
    .B(_02025_),
    .Y(_02073_));
 sky130_fd_sc_hd__a21o_1 _07981_ (.A1(_02072_),
    .A2(_02064_),
    .B1(_02073_),
    .X(_02074_));
 sky130_fd_sc_hd__a21o_1 _07982_ (.A1(_02014_),
    .A2(_01955_),
    .B1(_01962_),
    .X(_02075_));
 sky130_fd_sc_hd__nand3_2 _07983_ (.A(_02074_),
    .B(_02015_),
    .C(_02075_),
    .Y(_02076_));
 sky130_fd_sc_hd__nand2_1 _07984_ (.A(_02022_),
    .B(_02076_),
    .Y(_02077_));
 sky130_fd_sc_hd__inv_2 _07985_ (.A(_02076_),
    .Y(_02078_));
 sky130_fd_sc_hd__nand3_2 _07986_ (.A(_02020_),
    .B(_02078_),
    .C(_02021_),
    .Y(_02079_));
 sky130_fd_sc_hd__nand2_1 _07987_ (.A(_02044_),
    .B(_02057_),
    .Y(_02080_));
 sky130_fd_sc_hd__nand2_1 _07988_ (.A(_02080_),
    .B(_02055_),
    .Y(_02081_));
 sky130_fd_sc_hd__nand3_1 _07989_ (.A(_02044_),
    .B(_02057_),
    .C(_02056_),
    .Y(_02083_));
 sky130_fd_sc_hd__nand2_1 _07990_ (.A(_02081_),
    .B(_02083_),
    .Y(_02084_));
 sky130_fd_sc_hd__inv_2 _07991_ (.A(_04827_),
    .Y(_02085_));
 sky130_fd_sc_hd__inv_2 _07992_ (.A(_01092_),
    .Y(_02086_));
 sky130_fd_sc_hd__nand2_1 _07993_ (.A(_04911_),
    .B(_04260_),
    .Y(_02087_));
 sky130_fd_sc_hd__nor3_1 _07994_ (.A(_02085_),
    .B(_02086_),
    .C(_02087_),
    .Y(_02088_));
 sky130_fd_sc_hd__inv_2 _07995_ (.A(_02088_),
    .Y(_02089_));
 sky130_fd_sc_hd__o21ai_1 _07996_ (.A1(_02085_),
    .A2(_02086_),
    .B1(_02087_),
    .Y(_02090_));
 sky130_fd_sc_hd__nand2_1 _07997_ (.A(_04895_),
    .B(_01565_),
    .Y(_02091_));
 sky130_fd_sc_hd__inv_2 _07998_ (.A(_02091_),
    .Y(_02092_));
 sky130_fd_sc_hd__a21o_1 _07999_ (.A1(_02089_),
    .A2(_02090_),
    .B1(_02092_),
    .X(_02094_));
 sky130_fd_sc_hd__nand3_1 _08000_ (.A(_02089_),
    .B(_02092_),
    .C(_02090_),
    .Y(_02095_));
 sky130_fd_sc_hd__nand2_1 _08001_ (.A(_02094_),
    .B(_02095_),
    .Y(_02096_));
 sky130_fd_sc_hd__inv_2 _08002_ (.A(_02096_),
    .Y(_02097_));
 sky130_fd_sc_hd__xnor2_1 _08003_ (.A(_02035_),
    .B(_02041_),
    .Y(_02098_));
 sky130_fd_sc_hd__a22o_1 _08004_ (.A1(_00254_),
    .A2(_02379_),
    .B1(_00522_),
    .B2(_02357_),
    .X(_02099_));
 sky130_fd_sc_hd__nand2_1 _08005_ (.A(_04828_),
    .B(_01535_),
    .Y(_02100_));
 sky130_fd_sc_hd__inv_2 _08006_ (.A(_02100_),
    .Y(_02101_));
 sky130_fd_sc_hd__and4_1 _08007_ (.A(_00254_),
    .B(_00522_),
    .C(_02379_),
    .D(_02357_),
    .X(_02102_));
 sky130_fd_sc_hd__a21oi_1 _08008_ (.A1(_02099_),
    .A2(_02101_),
    .B1(_02102_),
    .Y(_02103_));
 sky130_fd_sc_hd__nand2_1 _08009_ (.A(_02098_),
    .B(_02103_),
    .Y(_02105_));
 sky130_fd_sc_hd__nor2_1 _08010_ (.A(_02103_),
    .B(_02098_),
    .Y(_02106_));
 sky130_fd_sc_hd__a21oi_1 _08011_ (.A1(_02097_),
    .A2(_02105_),
    .B1(_02106_),
    .Y(_02107_));
 sky130_fd_sc_hd__nand2_1 _08012_ (.A(_02084_),
    .B(_02107_),
    .Y(_02108_));
 sky130_fd_sc_hd__nand2_1 _08013_ (.A(_04895_),
    .B(_00204_),
    .Y(_02109_));
 sky130_fd_sc_hd__and2_1 _08014_ (.A(_02095_),
    .B(_02089_),
    .X(_02110_));
 sky130_fd_sc_hd__nor2_2 _08015_ (.A(_02109_),
    .B(_02110_),
    .Y(_02111_));
 sky130_fd_sc_hd__inv_2 _08016_ (.A(_02111_),
    .Y(_02112_));
 sky130_fd_sc_hd__nand2_1 _08017_ (.A(_02110_),
    .B(_02109_),
    .Y(_02113_));
 sky130_fd_sc_hd__nand2_1 _08018_ (.A(_02112_),
    .B(_02113_),
    .Y(_02114_));
 sky130_fd_sc_hd__inv_2 _08019_ (.A(_02114_),
    .Y(_02116_));
 sky130_fd_sc_hd__nor2_1 _08020_ (.A(_02107_),
    .B(_02084_),
    .Y(_02117_));
 sky130_fd_sc_hd__a21oi_1 _08021_ (.A1(_02108_),
    .A2(_02116_),
    .B1(_02117_),
    .Y(_02118_));
 sky130_fd_sc_hd__inv_2 _08022_ (.A(_02118_),
    .Y(_02119_));
 sky130_fd_sc_hd__inv_2 _08023_ (.A(_02030_),
    .Y(_02120_));
 sky130_fd_sc_hd__inv_2 _08024_ (.A(_02058_),
    .Y(_02121_));
 sky130_fd_sc_hd__nand2_1 _08025_ (.A(_02120_),
    .B(_02121_),
    .Y(_02122_));
 sky130_fd_sc_hd__nand3_1 _08026_ (.A(_02122_),
    .B(_02059_),
    .C(_02068_),
    .Y(_02123_));
 sky130_fd_sc_hd__nand2_1 _08027_ (.A(_02122_),
    .B(_02059_),
    .Y(_02124_));
 sky130_fd_sc_hd__nand2_1 _08028_ (.A(_02124_),
    .B(_02067_),
    .Y(_02125_));
 sky130_fd_sc_hd__nand3_2 _08029_ (.A(_02119_),
    .B(_02123_),
    .C(_02125_),
    .Y(_02127_));
 sky130_fd_sc_hd__nand2_1 _08030_ (.A(_02125_),
    .B(_02123_),
    .Y(_02128_));
 sky130_fd_sc_hd__nand2_1 _08031_ (.A(_02128_),
    .B(_02118_),
    .Y(_02129_));
 sky130_fd_sc_hd__nand3_2 _08032_ (.A(_02127_),
    .B(_02129_),
    .C(_02111_),
    .Y(_02130_));
 sky130_fd_sc_hd__nand2_1 _08033_ (.A(_02130_),
    .B(_02127_),
    .Y(_02131_));
 sky130_fd_sc_hd__inv_2 _08034_ (.A(_02070_),
    .Y(_02132_));
 sky130_fd_sc_hd__nand3_1 _08035_ (.A(_02132_),
    .B(_02009_),
    .C(_02024_),
    .Y(_02133_));
 sky130_fd_sc_hd__nand3_1 _08036_ (.A(_02133_),
    .B(_02064_),
    .C(_02072_),
    .Y(_02134_));
 sky130_fd_sc_hd__nand2_1 _08037_ (.A(_02133_),
    .B(_02072_),
    .Y(_02135_));
 sky130_fd_sc_hd__nand2_1 _08038_ (.A(_02135_),
    .B(_02065_),
    .Y(_02136_));
 sky130_fd_sc_hd__nand3_2 _08039_ (.A(_02131_),
    .B(_02134_),
    .C(_02136_),
    .Y(_02138_));
 sky130_fd_sc_hd__nand2_1 _08040_ (.A(_02075_),
    .B(_02015_),
    .Y(_02139_));
 sky130_fd_sc_hd__a21oi_1 _08041_ (.A1(_02072_),
    .A2(_02064_),
    .B1(_02073_),
    .Y(_02140_));
 sky130_fd_sc_hd__nand2_1 _08042_ (.A(_02139_),
    .B(_02140_),
    .Y(_02141_));
 sky130_fd_sc_hd__nand2_1 _08043_ (.A(_02076_),
    .B(_02141_),
    .Y(_02142_));
 sky130_fd_sc_hd__nor2_1 _08044_ (.A(_02138_),
    .B(_02142_),
    .Y(_02143_));
 sky130_fd_sc_hd__nand3_2 _08045_ (.A(_02077_),
    .B(_02079_),
    .C(_02143_),
    .Y(_02144_));
 sky130_fd_sc_hd__inv_2 _08046_ (.A(_02144_),
    .Y(_02145_));
 sky130_fd_sc_hd__a21o_1 _08047_ (.A1(_01965_),
    .A2(_01959_),
    .B1(_01966_),
    .X(_02146_));
 sky130_fd_sc_hd__nand3_1 _08048_ (.A(_02146_),
    .B(_01973_),
    .C(_01974_),
    .Y(_02147_));
 sky130_fd_sc_hd__nand2_1 _08049_ (.A(_01975_),
    .B(_01967_),
    .Y(_02149_));
 sky130_fd_sc_hd__nand2_1 _08050_ (.A(_02147_),
    .B(_02149_),
    .Y(_02150_));
 sky130_fd_sc_hd__nand2_1 _08051_ (.A(_02150_),
    .B(_02079_),
    .Y(_02151_));
 sky130_fd_sc_hd__inv_2 _08052_ (.A(_02079_),
    .Y(_02152_));
 sky130_fd_sc_hd__nand3_2 _08053_ (.A(_02152_),
    .B(_02147_),
    .C(_02149_),
    .Y(_02153_));
 sky130_fd_sc_hd__nand3_2 _08054_ (.A(_02145_),
    .B(_02151_),
    .C(_02153_),
    .Y(_02154_));
 sky130_fd_sc_hd__nand2_1 _08055_ (.A(_01880_),
    .B(_01979_),
    .Y(_02155_));
 sky130_fd_sc_hd__nand2_1 _08056_ (.A(_02155_),
    .B(_02147_),
    .Y(_02156_));
 sky130_fd_sc_hd__nand2_1 _08057_ (.A(_02156_),
    .B(_01980_),
    .Y(_02157_));
 sky130_fd_sc_hd__nand2_1 _08058_ (.A(_02157_),
    .B(_02153_),
    .Y(_02158_));
 sky130_fd_sc_hd__nor2_1 _08059_ (.A(_02079_),
    .B(_02150_),
    .Y(_02160_));
 sky130_fd_sc_hd__nand3_1 _08060_ (.A(_02160_),
    .B(_02156_),
    .C(_01980_),
    .Y(_02161_));
 sky130_fd_sc_hd__nand2_1 _08061_ (.A(_02158_),
    .B(_02161_),
    .Y(_02162_));
 sky130_fd_sc_hd__nor2_1 _08062_ (.A(_02154_),
    .B(_02162_),
    .Y(_02163_));
 sky130_fd_sc_hd__inv_2 _08063_ (.A(_01980_),
    .Y(_02164_));
 sky130_fd_sc_hd__nand3_1 _08064_ (.A(_02164_),
    .B(_01988_),
    .C(_01986_),
    .Y(_02165_));
 sky130_fd_sc_hd__nand2_1 _08065_ (.A(_01989_),
    .B(_01980_),
    .Y(_02166_));
 sky130_fd_sc_hd__nand2_1 _08066_ (.A(_02165_),
    .B(_02166_),
    .Y(_02167_));
 sky130_fd_sc_hd__nand2_1 _08067_ (.A(_02167_),
    .B(_02161_),
    .Y(_02168_));
 sky130_fd_sc_hd__nor2_1 _08068_ (.A(_02153_),
    .B(_02157_),
    .Y(_02169_));
 sky130_fd_sc_hd__nand3_1 _08069_ (.A(_02169_),
    .B(_02165_),
    .C(_02166_),
    .Y(_02171_));
 sky130_fd_sc_hd__a21boi_1 _08070_ (.A1(_02163_),
    .A2(_02168_),
    .B1_N(_02171_),
    .Y(_02172_));
 sky130_fd_sc_hd__nand2_1 _08071_ (.A(_01995_),
    .B(_01997_),
    .Y(_02173_));
 sky130_fd_sc_hd__nand2_1 _08072_ (.A(_02173_),
    .B(_02165_),
    .Y(_02174_));
 sky130_fd_sc_hd__nand2_1 _08073_ (.A(_02174_),
    .B(_01998_),
    .Y(_02175_));
 sky130_fd_sc_hd__inv_2 _08074_ (.A(_02175_),
    .Y(_02176_));
 sky130_fd_sc_hd__nand3_1 _08075_ (.A(_02176_),
    .B(_02004_),
    .C(_02002_),
    .Y(_02177_));
 sky130_fd_sc_hd__nor2_1 _08076_ (.A(_02172_),
    .B(_02177_),
    .Y(_02178_));
 sky130_fd_sc_hd__nor2_1 _08077_ (.A(_02007_),
    .B(_02178_),
    .Y(_02179_));
 sky130_fd_sc_hd__inv_2 _08078_ (.A(_02154_),
    .Y(_02180_));
 sky130_fd_sc_hd__nand3_1 _08079_ (.A(_02180_),
    .B(_02161_),
    .C(_02158_),
    .Y(_02182_));
 sky130_fd_sc_hd__nand2_1 _08080_ (.A(_02162_),
    .B(_02154_),
    .Y(_02183_));
 sky130_fd_sc_hd__nand2_1 _08081_ (.A(_02182_),
    .B(_02183_),
    .Y(_02184_));
 sky130_fd_sc_hd__inv_2 _08082_ (.A(_02184_),
    .Y(_02185_));
 sky130_fd_sc_hd__nand2_1 _08083_ (.A(_02168_),
    .B(_02171_),
    .Y(_02186_));
 sky130_fd_sc_hd__inv_2 _08084_ (.A(_02186_),
    .Y(_02187_));
 sky130_fd_sc_hd__nand2_1 _08085_ (.A(_02185_),
    .B(_02187_),
    .Y(_02188_));
 sky130_fd_sc_hd__nor2_1 _08086_ (.A(_02188_),
    .B(_02177_),
    .Y(_02189_));
 sky130_fd_sc_hd__nand2_1 _08087_ (.A(_02077_),
    .B(_02079_),
    .Y(_02190_));
 sky130_fd_sc_hd__nand2_1 _08088_ (.A(_02136_),
    .B(_02134_),
    .Y(_02191_));
 sky130_fd_sc_hd__a21boi_1 _08089_ (.A1(_02111_),
    .A2(_02129_),
    .B1_N(_02127_),
    .Y(_02193_));
 sky130_fd_sc_hd__nor2_1 _08090_ (.A(_02191_),
    .B(_02193_),
    .Y(_02194_));
 sky130_fd_sc_hd__nand3_1 _08091_ (.A(_02194_),
    .B(_02076_),
    .C(_02141_),
    .Y(_02195_));
 sky130_fd_sc_hd__nand2_1 _08092_ (.A(_02190_),
    .B(_02195_),
    .Y(_02196_));
 sky130_fd_sc_hd__nand2_1 _08093_ (.A(_02196_),
    .B(_02144_),
    .Y(_02197_));
 sky130_fd_sc_hd__a21o_1 _08094_ (.A1(_02127_),
    .A2(_02129_),
    .B1(_02111_),
    .X(_02198_));
 sky130_fd_sc_hd__nand2b_1 _08095_ (.A_N(_02106_),
    .B(_02105_),
    .Y(_02199_));
 sky130_fd_sc_hd__xor2_1 _08096_ (.A(_02097_),
    .B(_02199_),
    .X(_02200_));
 sky130_fd_sc_hd__nand2_1 _08097_ (.A(_04991_),
    .B(_01535_),
    .Y(_02201_));
 sky130_fd_sc_hd__and4_1 _08098_ (.A(_00522_),
    .B(_04828_),
    .C(_02379_),
    .D(_02357_),
    .X(_02202_));
 sky130_fd_sc_hd__a22o_1 _08099_ (.A1(_00522_),
    .A2(_02379_),
    .B1(_04828_),
    .B2(_02357_),
    .X(_02204_));
 sky130_fd_sc_hd__nand2b_1 _08100_ (.A_N(_02202_),
    .B(_02204_),
    .Y(_02205_));
 sky130_fd_sc_hd__o21ba_1 _08101_ (.A1(_02201_),
    .A2(_02205_),
    .B1_N(_02202_),
    .X(_02206_));
 sky130_fd_sc_hd__nor2b_1 _08102_ (.A(_02102_),
    .B_N(_02099_),
    .Y(_02207_));
 sky130_fd_sc_hd__xor2_1 _08103_ (.A(_02100_),
    .B(_02207_),
    .X(_02208_));
 sky130_fd_sc_hd__nand2_1 _08104_ (.A(_02206_),
    .B(_02208_),
    .Y(_02209_));
 sky130_fd_sc_hd__and4_1 _08105_ (.A(_04991_),
    .B(_04992_),
    .C(_04293_),
    .D(_04260_),
    .X(_02210_));
 sky130_fd_sc_hd__inv_2 _08106_ (.A(_02210_),
    .Y(_02211_));
 sky130_fd_sc_hd__a22o_1 _08107_ (.A1(_04991_),
    .A2(_04293_),
    .B1(_04992_),
    .B2(_04260_),
    .X(_02212_));
 sky130_fd_sc_hd__and2_1 _08108_ (.A(_02211_),
    .B(_02212_),
    .X(_02213_));
 sky130_fd_sc_hd__nor2_1 _08109_ (.A(_02208_),
    .B(_02206_),
    .Y(_02215_));
 sky130_fd_sc_hd__a21oi_1 _08110_ (.A1(_02209_),
    .A2(_02213_),
    .B1(_02215_),
    .Y(_02216_));
 sky130_fd_sc_hd__nand2_1 _08111_ (.A(_02200_),
    .B(_02216_),
    .Y(_02217_));
 sky130_fd_sc_hd__nor2_1 _08112_ (.A(_02216_),
    .B(_02200_),
    .Y(_02218_));
 sky130_fd_sc_hd__a21oi_1 _08113_ (.A1(_02217_),
    .A2(_02210_),
    .B1(_02218_),
    .Y(_02219_));
 sky130_fd_sc_hd__nand2b_1 _08114_ (.A_N(_02117_),
    .B(_02108_),
    .Y(_02220_));
 sky130_fd_sc_hd__or2_1 _08115_ (.A(_02114_),
    .B(_02220_),
    .X(_02221_));
 sky130_fd_sc_hd__nand2_1 _08116_ (.A(_02220_),
    .B(_02114_),
    .Y(_02222_));
 sky130_fd_sc_hd__nand2_1 _08117_ (.A(_02221_),
    .B(_02222_),
    .Y(_02223_));
 sky130_fd_sc_hd__nor2_1 _08118_ (.A(_02219_),
    .B(_02223_),
    .Y(_02224_));
 sky130_fd_sc_hd__nand3_2 _08119_ (.A(_02198_),
    .B(_02130_),
    .C(_02224_),
    .Y(_02226_));
 sky130_fd_sc_hd__nand2_1 _08120_ (.A(_02193_),
    .B(_02191_),
    .Y(_02227_));
 sky130_fd_sc_hd__nand2_1 _08121_ (.A(_02138_),
    .B(_02227_),
    .Y(_02228_));
 sky130_fd_sc_hd__nor2_1 _08122_ (.A(_02226_),
    .B(_02228_),
    .Y(_02229_));
 sky130_fd_sc_hd__nand2_1 _08123_ (.A(_02142_),
    .B(_02138_),
    .Y(_02230_));
 sky130_fd_sc_hd__nand3_1 _08124_ (.A(_02229_),
    .B(_02195_),
    .C(_02230_),
    .Y(_02231_));
 sky130_fd_sc_hd__nand2_1 _08125_ (.A(_02197_),
    .B(_02231_),
    .Y(_02232_));
 sky130_fd_sc_hd__inv_2 _08126_ (.A(_02226_),
    .Y(_02233_));
 sky130_fd_sc_hd__nand3_2 _08127_ (.A(_02233_),
    .B(_02138_),
    .C(_02227_),
    .Y(_02234_));
 sky130_fd_sc_hd__nand2_1 _08128_ (.A(_02195_),
    .B(_02230_),
    .Y(_02235_));
 sky130_fd_sc_hd__nor2_1 _08129_ (.A(_02234_),
    .B(_02235_),
    .Y(_02237_));
 sky130_fd_sc_hd__nand3_2 _08130_ (.A(_02196_),
    .B(_02144_),
    .C(_02237_),
    .Y(_02238_));
 sky130_fd_sc_hd__nand2_1 _08131_ (.A(_02232_),
    .B(_02238_),
    .Y(_02239_));
 sky130_fd_sc_hd__nand2_1 _08132_ (.A(_02235_),
    .B(_02234_),
    .Y(_02240_));
 sky130_fd_sc_hd__nand2_1 _08133_ (.A(_02231_),
    .B(_02240_),
    .Y(_02241_));
 sky130_fd_sc_hd__nand2_1 _08134_ (.A(_02198_),
    .B(_02130_),
    .Y(_02242_));
 sky130_fd_sc_hd__nand3b_1 _08135_ (.A_N(_02219_),
    .B(_02221_),
    .C(_02222_),
    .Y(_02243_));
 sky130_fd_sc_hd__nand2_1 _08136_ (.A(_02242_),
    .B(_02243_),
    .Y(_02244_));
 sky130_fd_sc_hd__nand2b_1 _08137_ (.A_N(_02215_),
    .B(_02209_),
    .Y(_02245_));
 sky130_fd_sc_hd__xor2_1 _08138_ (.A(_02213_),
    .B(_02245_),
    .X(_02246_));
 sky130_fd_sc_hd__nand2_1 _08139_ (.A(_04992_),
    .B(_04293_),
    .Y(_02248_));
 sky130_fd_sc_hd__nand2_1 _08140_ (.A(_04992_),
    .B(_01535_),
    .Y(_02249_));
 sky130_fd_sc_hd__nand2_1 _08141_ (.A(_04991_),
    .B(_02357_),
    .Y(_02250_));
 sky130_fd_sc_hd__or3_1 _08142_ (.A(_02085_),
    .B(_01597_),
    .C(_02250_),
    .X(_02251_));
 sky130_fd_sc_hd__o21ai_1 _08143_ (.A1(_02085_),
    .A2(_01597_),
    .B1(_02250_),
    .Y(_02252_));
 sky130_fd_sc_hd__nand2_1 _08144_ (.A(_02251_),
    .B(_02252_),
    .Y(_02253_));
 sky130_fd_sc_hd__o21a_1 _08145_ (.A1(_02249_),
    .A2(_02253_),
    .B1(_02251_),
    .X(_02254_));
 sky130_fd_sc_hd__or2_1 _08146_ (.A(_02201_),
    .B(_02205_),
    .X(_02255_));
 sky130_fd_sc_hd__nand2_1 _08147_ (.A(_02205_),
    .B(_02201_),
    .Y(_02256_));
 sky130_fd_sc_hd__nand2_1 _08148_ (.A(_02255_),
    .B(_02256_),
    .Y(_02257_));
 sky130_fd_sc_hd__nor2_1 _08149_ (.A(_02254_),
    .B(_02257_),
    .Y(_02259_));
 sky130_fd_sc_hd__inv_2 _08150_ (.A(_02259_),
    .Y(_02260_));
 sky130_fd_sc_hd__nand2_1 _08151_ (.A(_02257_),
    .B(_02254_),
    .Y(_02261_));
 sky130_fd_sc_hd__nand2_1 _08152_ (.A(_02260_),
    .B(_02261_),
    .Y(_02262_));
 sky130_fd_sc_hd__or2_1 _08153_ (.A(_02248_),
    .B(_02262_),
    .X(_02263_));
 sky130_fd_sc_hd__and2_1 _08154_ (.A(_02263_),
    .B(_02260_),
    .X(_02264_));
 sky130_fd_sc_hd__nor2_1 _08155_ (.A(_02246_),
    .B(_02264_),
    .Y(_02265_));
 sky130_fd_sc_hd__nand2b_1 _08156_ (.A_N(_02218_),
    .B(_02217_),
    .Y(_02266_));
 sky130_fd_sc_hd__nand2_1 _08157_ (.A(_02266_),
    .B(_02211_),
    .Y(_02267_));
 sky130_fd_sc_hd__nand3b_1 _08158_ (.A_N(_02218_),
    .B(_02210_),
    .C(_02217_),
    .Y(_02268_));
 sky130_fd_sc_hd__nand3_1 _08159_ (.A(_02265_),
    .B(_02267_),
    .C(_02268_),
    .Y(_02270_));
 sky130_fd_sc_hd__nand2_1 _08160_ (.A(_02223_),
    .B(_02219_),
    .Y(_02271_));
 sky130_fd_sc_hd__nand2_1 _08161_ (.A(_02243_),
    .B(_02271_),
    .Y(_02272_));
 sky130_fd_sc_hd__nor2_1 _08162_ (.A(_02270_),
    .B(_02272_),
    .Y(_02273_));
 sky130_fd_sc_hd__nand3_1 _08163_ (.A(_02244_),
    .B(_02273_),
    .C(_02226_),
    .Y(_02274_));
 sky130_fd_sc_hd__nand2_1 _08164_ (.A(_02228_),
    .B(_02226_),
    .Y(_02275_));
 sky130_fd_sc_hd__nand3b_1 _08165_ (.A_N(_02274_),
    .B(_02234_),
    .C(_02275_),
    .Y(_02276_));
 sky130_fd_sc_hd__nor2_1 _08166_ (.A(_02241_),
    .B(_02276_),
    .Y(_02277_));
 sky130_fd_sc_hd__inv_2 _08167_ (.A(_02277_),
    .Y(_02278_));
 sky130_fd_sc_hd__nand2_1 _08168_ (.A(_02239_),
    .B(_02278_),
    .Y(_02279_));
 sky130_fd_sc_hd__nand3_2 _08169_ (.A(_02277_),
    .B(_02232_),
    .C(_02238_),
    .Y(_02281_));
 sky130_fd_sc_hd__nand2_1 _08170_ (.A(_02279_),
    .B(_02281_),
    .Y(_02282_));
 sky130_fd_sc_hd__nand2_1 _08171_ (.A(_02151_),
    .B(_02153_),
    .Y(_02283_));
 sky130_fd_sc_hd__nand2_1 _08172_ (.A(_02283_),
    .B(_02144_),
    .Y(_02284_));
 sky130_fd_sc_hd__nand2_1 _08173_ (.A(_02284_),
    .B(_02154_),
    .Y(_02285_));
 sky130_fd_sc_hd__nand2_1 _08174_ (.A(_02285_),
    .B(_02238_),
    .Y(_02286_));
 sky130_fd_sc_hd__inv_2 _08175_ (.A(_02238_),
    .Y(_02287_));
 sky130_fd_sc_hd__nand3_1 _08176_ (.A(_02287_),
    .B(_02284_),
    .C(_02154_),
    .Y(_02288_));
 sky130_fd_sc_hd__nand2_1 _08177_ (.A(_02286_),
    .B(_02288_),
    .Y(_02289_));
 sky130_fd_sc_hd__nor2_1 _08178_ (.A(_02282_),
    .B(_02289_),
    .Y(_02290_));
 sky130_fd_sc_hd__and2_1 _08179_ (.A(_02272_),
    .B(_02270_),
    .X(_02292_));
 sky130_fd_sc_hd__nand2_1 _08180_ (.A(_02264_),
    .B(_02246_),
    .Y(_02293_));
 sky130_fd_sc_hd__inv_2 _08181_ (.A(_02293_),
    .Y(_02294_));
 sky130_fd_sc_hd__a2111o_1 _08182_ (.A1(_02085_),
    .A2(_01535_),
    .B1(_01956_),
    .C1(_01597_),
    .D1(_02250_),
    .X(_02295_));
 sky130_fd_sc_hd__a21oi_1 _08183_ (.A1(_02249_),
    .A2(_02253_),
    .B1(_02295_),
    .Y(_02296_));
 sky130_fd_sc_hd__nand2_1 _08184_ (.A(_02263_),
    .B(_02296_),
    .Y(_02297_));
 sky130_fd_sc_hd__a21o_1 _08185_ (.A1(_02248_),
    .A2(_02262_),
    .B1(_02297_),
    .X(_02298_));
 sky130_fd_sc_hd__nor3_1 _08186_ (.A(_02265_),
    .B(_02294_),
    .C(_02298_),
    .Y(_02299_));
 sky130_fd_sc_hd__a21o_1 _08187_ (.A1(_02267_),
    .A2(_02268_),
    .B1(_02265_),
    .X(_02300_));
 sky130_fd_sc_hd__nand3_1 _08188_ (.A(_02299_),
    .B(_02270_),
    .C(_02300_),
    .Y(_02301_));
 sky130_fd_sc_hd__nor3_1 _08189_ (.A(_02273_),
    .B(_02292_),
    .C(_02301_),
    .Y(_02303_));
 sky130_fd_sc_hd__a21o_1 _08190_ (.A1(_02244_),
    .A2(_02226_),
    .B1(_02273_),
    .X(_02304_));
 sky130_fd_sc_hd__nand3_1 _08191_ (.A(_02303_),
    .B(_02304_),
    .C(_02274_),
    .Y(_02305_));
 sky130_fd_sc_hd__inv_2 _08192_ (.A(_02305_),
    .Y(_02306_));
 sky130_fd_sc_hd__inv_2 _08193_ (.A(_02241_),
    .Y(_02307_));
 sky130_fd_sc_hd__nand2_1 _08194_ (.A(_02234_),
    .B(_02275_),
    .Y(_02308_));
 sky130_fd_sc_hd__nand2_1 _08195_ (.A(_02308_),
    .B(_02274_),
    .Y(_02309_));
 sky130_fd_sc_hd__and4_1 _08196_ (.A(_02306_),
    .B(_02307_),
    .C(_02276_),
    .D(_02309_),
    .X(_02310_));
 sky130_fd_sc_hd__nand2_1 _08197_ (.A(_02290_),
    .B(_02310_),
    .Y(_02311_));
 sky130_fd_sc_hd__inv_2 _08198_ (.A(_02281_),
    .Y(_02312_));
 sky130_fd_sc_hd__a21boi_1 _08199_ (.A1(_02312_),
    .A2(_02286_),
    .B1_N(_02288_),
    .Y(_02314_));
 sky130_fd_sc_hd__nand2_1 _08200_ (.A(_02311_),
    .B(_02314_),
    .Y(_02315_));
 sky130_fd_sc_hd__nand2_1 _08201_ (.A(_02189_),
    .B(_02315_),
    .Y(_02316_));
 sky130_fd_sc_hd__nand2_2 _08202_ (.A(_02179_),
    .B(_02316_),
    .Y(_02317_));
 sky130_fd_sc_hd__xor2_1 _08203_ (.A(_01711_),
    .B(_01737_),
    .X(_02318_));
 sky130_fd_sc_hd__inv_2 _08204_ (.A(_02318_),
    .Y(_02319_));
 sky130_fd_sc_hd__nand2_1 _08205_ (.A(_01709_),
    .B(_01711_),
    .Y(_02320_));
 sky130_fd_sc_hd__nand2_1 _08206_ (.A(_02320_),
    .B(_01678_),
    .Y(_02321_));
 sky130_fd_sc_hd__nand2_1 _08207_ (.A(_02321_),
    .B(_01712_),
    .Y(_02322_));
 sky130_fd_sc_hd__inv_2 _08208_ (.A(_02322_),
    .Y(_02323_));
 sky130_fd_sc_hd__and3_1 _08209_ (.A(_02319_),
    .B(_01767_),
    .C(_02323_),
    .X(_02325_));
 sky130_fd_sc_hd__nand3_1 _08210_ (.A(_01782_),
    .B(_02317_),
    .C(_02325_),
    .Y(_02326_));
 sky130_fd_sc_hd__nand2_2 _08211_ (.A(_01781_),
    .B(_02326_),
    .Y(_02327_));
 sky130_fd_sc_hd__inv_2 _08212_ (.A(_00390_),
    .Y(_02328_));
 sky130_fd_sc_hd__a21boi_1 _08213_ (.A1(_02328_),
    .A2(_00406_),
    .B1_N(_00407_),
    .Y(_02329_));
 sky130_fd_sc_hd__nand2_1 _08214_ (.A(_00861_),
    .B(_05160_),
    .Y(_02330_));
 sky130_fd_sc_hd__inv_2 _08215_ (.A(_02330_),
    .Y(_02331_));
 sky130_fd_sc_hd__nand2_1 _08216_ (.A(_00751_),
    .B(_00393_),
    .Y(_02332_));
 sky130_fd_sc_hd__nand2_1 _08217_ (.A(_00795_),
    .B(net17),
    .Y(_02333_));
 sky130_fd_sc_hd__nor2_1 _08218_ (.A(_02332_),
    .B(_02333_),
    .Y(_02334_));
 sky130_fd_sc_hd__nand2_1 _08219_ (.A(_02332_),
    .B(_02333_),
    .Y(_02336_));
 sky130_fd_sc_hd__inv_2 _08220_ (.A(_02336_),
    .Y(_02337_));
 sky130_fd_sc_hd__nor2_1 _08221_ (.A(_02334_),
    .B(_02337_),
    .Y(_02338_));
 sky130_fd_sc_hd__or2_1 _08222_ (.A(_02331_),
    .B(_02338_),
    .X(_02339_));
 sky130_fd_sc_hd__nand2_1 _08223_ (.A(_02338_),
    .B(_02331_),
    .Y(_02340_));
 sky130_fd_sc_hd__nand2_1 _08224_ (.A(_02339_),
    .B(_02340_),
    .Y(_02341_));
 sky130_fd_sc_hd__nand2_1 _08225_ (.A(_00401_),
    .B(_00396_),
    .Y(_02342_));
 sky130_fd_sc_hd__inv_2 _08226_ (.A(_02342_),
    .Y(_02343_));
 sky130_fd_sc_hd__nand2_1 _08227_ (.A(_02341_),
    .B(_02343_),
    .Y(_02344_));
 sky130_fd_sc_hd__nand3_2 _08228_ (.A(_02339_),
    .B(_02342_),
    .C(_02340_),
    .Y(_02345_));
 sky130_fd_sc_hd__nand2_1 _08229_ (.A(_02344_),
    .B(_02345_),
    .Y(_02347_));
 sky130_fd_sc_hd__nand2_1 _08230_ (.A(_00784_),
    .B(_01565_),
    .Y(_02348_));
 sky130_fd_sc_hd__inv_2 _08231_ (.A(_02348_),
    .Y(_02349_));
 sky130_fd_sc_hd__nand2_1 _08232_ (.A(_01323_),
    .B(_01048_),
    .Y(_02350_));
 sky130_fd_sc_hd__nand2_1 _08233_ (.A(_04293_),
    .B(_04084_),
    .Y(_02351_));
 sky130_fd_sc_hd__or2_1 _08234_ (.A(_02350_),
    .B(_02351_),
    .X(_02352_));
 sky130_fd_sc_hd__nand2_1 _08235_ (.A(_02350_),
    .B(_02351_),
    .Y(_02353_));
 sky130_fd_sc_hd__nand2_1 _08236_ (.A(_02352_),
    .B(_02353_),
    .Y(_02354_));
 sky130_fd_sc_hd__xor2_1 _08237_ (.A(_02349_),
    .B(_02354_),
    .X(_02355_));
 sky130_fd_sc_hd__nand2_1 _08238_ (.A(_02347_),
    .B(_02355_),
    .Y(_02356_));
 sky130_fd_sc_hd__inv_2 _08239_ (.A(_02355_),
    .Y(_02358_));
 sky130_fd_sc_hd__nand3_2 _08240_ (.A(_02344_),
    .B(_02358_),
    .C(_02345_),
    .Y(_02359_));
 sky130_fd_sc_hd__nand2_1 _08241_ (.A(_02356_),
    .B(_02359_),
    .Y(_02360_));
 sky130_fd_sc_hd__nor2_1 _08242_ (.A(_02329_),
    .B(_02360_),
    .Y(_02361_));
 sky130_fd_sc_hd__inv_2 _08243_ (.A(_02361_),
    .Y(_02362_));
 sky130_fd_sc_hd__nand2_1 _08244_ (.A(_02360_),
    .B(_02329_),
    .Y(_02363_));
 sky130_fd_sc_hd__nand2_1 _08245_ (.A(_02362_),
    .B(_02363_),
    .Y(_02364_));
 sky130_fd_sc_hd__nand2_1 _08246_ (.A(_01081_),
    .B(_00003_),
    .Y(_02365_));
 sky130_fd_sc_hd__nand2_1 _08247_ (.A(_00850_),
    .B(_01774_),
    .Y(_02366_));
 sky130_fd_sc_hd__nand2_1 _08248_ (.A(_00740_),
    .B(_01807_),
    .Y(_02367_));
 sky130_fd_sc_hd__or2_1 _08249_ (.A(_02366_),
    .B(_02367_),
    .X(_02369_));
 sky130_fd_sc_hd__nand2_1 _08250_ (.A(_02366_),
    .B(_02367_),
    .Y(_02370_));
 sky130_fd_sc_hd__nand2_1 _08251_ (.A(_02369_),
    .B(_02370_),
    .Y(_02371_));
 sky130_fd_sc_hd__or2_1 _08252_ (.A(_02365_),
    .B(_02371_),
    .X(_02372_));
 sky130_fd_sc_hd__nand2_1 _08253_ (.A(_02371_),
    .B(_02365_),
    .Y(_02373_));
 sky130_fd_sc_hd__nand2_1 _08254_ (.A(_02372_),
    .B(_02373_),
    .Y(_02374_));
 sky130_fd_sc_hd__nand2_1 _08255_ (.A(_00389_),
    .B(_00382_),
    .Y(_02375_));
 sky130_fd_sc_hd__nand2_1 _08256_ (.A(_02374_),
    .B(_02375_),
    .Y(_02376_));
 sky130_fd_sc_hd__inv_2 _08257_ (.A(_02375_),
    .Y(_02377_));
 sky130_fd_sc_hd__nand3_1 _08258_ (.A(_02372_),
    .B(_02377_),
    .C(_02373_),
    .Y(_02378_));
 sky130_fd_sc_hd__nand2_1 _08259_ (.A(_02376_),
    .B(_02378_),
    .Y(_02380_));
 sky130_fd_sc_hd__nand2_1 _08260_ (.A(_00420_),
    .B(_00415_),
    .Y(_02381_));
 sky130_fd_sc_hd__nand2_1 _08261_ (.A(_02380_),
    .B(_02381_),
    .Y(_02382_));
 sky130_fd_sc_hd__nand3b_1 _08262_ (.A_N(_02381_),
    .B(_02376_),
    .C(_02378_),
    .Y(_02383_));
 sky130_fd_sc_hd__nand2_1 _08263_ (.A(_02382_),
    .B(_02383_),
    .Y(_02384_));
 sky130_fd_sc_hd__nand2_1 _08264_ (.A(_02364_),
    .B(_02384_),
    .Y(_02385_));
 sky130_fd_sc_hd__inv_2 _08265_ (.A(_02384_),
    .Y(_02386_));
 sky130_fd_sc_hd__nand3_2 _08266_ (.A(_02362_),
    .B(_02386_),
    .C(_02363_),
    .Y(_02387_));
 sky130_fd_sc_hd__nand2_1 _08267_ (.A(_02385_),
    .B(_02387_),
    .Y(_02388_));
 sky130_fd_sc_hd__nand2_2 _08268_ (.A(_00437_),
    .B(_00411_),
    .Y(_02389_));
 sky130_fd_sc_hd__inv_2 _08269_ (.A(_02389_),
    .Y(_02391_));
 sky130_fd_sc_hd__nand2_1 _08270_ (.A(_02388_),
    .B(_02391_),
    .Y(_02392_));
 sky130_fd_sc_hd__nand2_1 _08271_ (.A(net6),
    .B(_02995_),
    .Y(_02393_));
 sky130_fd_sc_hd__nand2_1 _08272_ (.A(_01037_),
    .B(_03028_),
    .Y(_02394_));
 sky130_fd_sc_hd__or2_1 _08273_ (.A(_02393_),
    .B(_02394_),
    .X(_02395_));
 sky130_fd_sc_hd__nand2_1 _08274_ (.A(_02393_),
    .B(_02394_),
    .Y(_02396_));
 sky130_fd_sc_hd__nand2_1 _08275_ (.A(_02395_),
    .B(_02396_),
    .Y(_02397_));
 sky130_fd_sc_hd__nand2_1 _08276_ (.A(_03215_),
    .B(_02544_),
    .Y(_02398_));
 sky130_fd_sc_hd__inv_2 _08277_ (.A(_02398_),
    .Y(_02399_));
 sky130_fd_sc_hd__nand2b_1 _08278_ (.A_N(_02397_),
    .B(_02399_),
    .Y(_02400_));
 sky130_fd_sc_hd__nand2_1 _08279_ (.A(_02397_),
    .B(_02398_),
    .Y(_02402_));
 sky130_fd_sc_hd__nand2_1 _08280_ (.A(_02400_),
    .B(_02402_),
    .Y(_02403_));
 sky130_fd_sc_hd__nand2_1 _08281_ (.A(_00453_),
    .B(_00447_),
    .Y(_02404_));
 sky130_fd_sc_hd__nand2_1 _08282_ (.A(_02403_),
    .B(_02404_),
    .Y(_02405_));
 sky130_fd_sc_hd__inv_2 _08283_ (.A(_02404_),
    .Y(_02406_));
 sky130_fd_sc_hd__nand3_1 _08284_ (.A(_02406_),
    .B(_02400_),
    .C(_02402_),
    .Y(_02407_));
 sky130_fd_sc_hd__nand2_1 _08285_ (.A(_02405_),
    .B(_02407_),
    .Y(_02408_));
 sky130_fd_sc_hd__nand2_1 _08286_ (.A(_03809_),
    .B(_02753_),
    .Y(_02409_));
 sky130_fd_sc_hd__inv_2 _08287_ (.A(_01873_),
    .Y(_02410_));
 sky130_fd_sc_hd__nand2_1 _08288_ (.A(_04962_),
    .B(_02049_),
    .Y(_02411_));
 sky130_fd_sc_hd__nor3_1 _08289_ (.A(_01330_),
    .B(_02410_),
    .C(_02411_),
    .Y(_02413_));
 sky130_fd_sc_hd__inv_2 _08290_ (.A(_02413_),
    .Y(_02414_));
 sky130_fd_sc_hd__o21ai_1 _08291_ (.A1(_01330_),
    .A2(_02410_),
    .B1(_02411_),
    .Y(_02415_));
 sky130_fd_sc_hd__nand2_1 _08292_ (.A(_02414_),
    .B(_02415_),
    .Y(_02416_));
 sky130_fd_sc_hd__or2_1 _08293_ (.A(_02409_),
    .B(_02416_),
    .X(_02417_));
 sky130_fd_sc_hd__nand2_1 _08294_ (.A(_02416_),
    .B(_02409_),
    .Y(_02418_));
 sky130_fd_sc_hd__nand3_1 _08295_ (.A(_02408_),
    .B(_02417_),
    .C(_02418_),
    .Y(_02419_));
 sky130_fd_sc_hd__nand2_1 _08296_ (.A(_02417_),
    .B(_02418_),
    .Y(_02420_));
 sky130_fd_sc_hd__nand3_1 _08297_ (.A(_02420_),
    .B(_02405_),
    .C(_02407_),
    .Y(_02421_));
 sky130_fd_sc_hd__nand2_1 _08298_ (.A(_02419_),
    .B(_02421_),
    .Y(_02422_));
 sky130_fd_sc_hd__nand2_1 _08299_ (.A(_00421_),
    .B(_00423_),
    .Y(_02424_));
 sky130_fd_sc_hd__nor2_1 _08300_ (.A(_00423_),
    .B(_00421_),
    .Y(_02425_));
 sky130_fd_sc_hd__a21oi_4 _08301_ (.A1(_02424_),
    .A2(_00428_),
    .B1(_02425_),
    .Y(_02426_));
 sky130_fd_sc_hd__inv_2 _08302_ (.A(_02426_),
    .Y(_02427_));
 sky130_fd_sc_hd__nand2_1 _08303_ (.A(_02422_),
    .B(_02427_),
    .Y(_02428_));
 sky130_fd_sc_hd__nand3_1 _08304_ (.A(_02419_),
    .B(_02421_),
    .C(_02426_),
    .Y(_02429_));
 sky130_fd_sc_hd__nand2_1 _08305_ (.A(_02428_),
    .B(_02429_),
    .Y(_02430_));
 sky130_fd_sc_hd__nand2_1 _08306_ (.A(_00470_),
    .B(_00469_),
    .Y(_02431_));
 sky130_fd_sc_hd__nand2_1 _08307_ (.A(_02430_),
    .B(_02431_),
    .Y(_02432_));
 sky130_fd_sc_hd__nand3b_1 _08308_ (.A_N(_02431_),
    .B(_02428_),
    .C(_02429_),
    .Y(_02433_));
 sky130_fd_sc_hd__nand2_1 _08309_ (.A(_02432_),
    .B(_02433_),
    .Y(_02435_));
 sky130_fd_sc_hd__inv_2 _08310_ (.A(_02435_),
    .Y(_02436_));
 sky130_fd_sc_hd__nand3_2 _08311_ (.A(_02385_),
    .B(_02389_),
    .C(_02387_),
    .Y(_02437_));
 sky130_fd_sc_hd__nand3_2 _08312_ (.A(_02392_),
    .B(_02436_),
    .C(_02437_),
    .Y(_02438_));
 sky130_fd_sc_hd__nand2_1 _08313_ (.A(_02388_),
    .B(_02389_),
    .Y(_02439_));
 sky130_fd_sc_hd__nand3_1 _08314_ (.A(_02385_),
    .B(_02391_),
    .C(_02387_),
    .Y(_02440_));
 sky130_fd_sc_hd__nand3_1 _08315_ (.A(_02439_),
    .B(_02435_),
    .C(_02440_),
    .Y(_02441_));
 sky130_fd_sc_hd__nand2_1 _08316_ (.A(_02438_),
    .B(_02441_),
    .Y(_02442_));
 sky130_fd_sc_hd__nand2_2 _08317_ (.A(_00487_),
    .B(_00441_),
    .Y(_02443_));
 sky130_fd_sc_hd__nand2_1 _08318_ (.A(_02442_),
    .B(_02443_),
    .Y(_02444_));
 sky130_fd_sc_hd__inv_2 _08319_ (.A(_02443_),
    .Y(_02446_));
 sky130_fd_sc_hd__nand3_1 _08320_ (.A(_02438_),
    .B(_02441_),
    .C(_02446_),
    .Y(_02447_));
 sky130_fd_sc_hd__nand2_1 _08321_ (.A(_02444_),
    .B(_02447_),
    .Y(_02448_));
 sky130_fd_sc_hd__and2_1 _08322_ (.A(_00525_),
    .B(_00519_),
    .X(_02449_));
 sky130_fd_sc_hd__nand2_1 _08323_ (.A(_04876_),
    .B(_04809_),
    .Y(_02450_));
 sky130_fd_sc_hd__inv_2 _08324_ (.A(_03402_),
    .Y(_02451_));
 sky130_fd_sc_hd__nand2_1 _08325_ (.A(_04871_),
    .B(_03820_),
    .Y(_02452_));
 sky130_fd_sc_hd__nor3_1 _08326_ (.A(_00110_),
    .B(_02451_),
    .C(_02452_),
    .Y(_02453_));
 sky130_fd_sc_hd__o21ai_1 _08327_ (.A1(_00110_),
    .A2(_02451_),
    .B1(_02452_),
    .Y(_02454_));
 sky130_fd_sc_hd__inv_2 _08328_ (.A(_02454_),
    .Y(_02455_));
 sky130_fd_sc_hd__nor2_1 _08329_ (.A(_02453_),
    .B(_02455_),
    .Y(_02457_));
 sky130_fd_sc_hd__xor2_1 _08330_ (.A(_02450_),
    .B(_02457_),
    .X(_02458_));
 sky130_fd_sc_hd__nor2_1 _08331_ (.A(_02449_),
    .B(_02458_),
    .Y(_02459_));
 sky130_fd_sc_hd__nand2_1 _08332_ (.A(_02458_),
    .B(_02449_),
    .Y(_02460_));
 sky130_fd_sc_hd__inv_2 _08333_ (.A(_02460_),
    .Y(_02461_));
 sky130_fd_sc_hd__nand2_1 _08334_ (.A(_00529_),
    .B(_04991_),
    .Y(_02462_));
 sky130_fd_sc_hd__inv_2 _08335_ (.A(net46),
    .Y(_02463_));
 sky130_fd_sc_hd__inv_2 _08336_ (.A(_04819_),
    .Y(_02464_));
 sky130_fd_sc_hd__nand2_1 _08337_ (.A(_00124_),
    .B(_04827_),
    .Y(_02465_));
 sky130_fd_sc_hd__nor3_1 _08338_ (.A(_02463_),
    .B(_02464_),
    .C(_02465_),
    .Y(_02466_));
 sky130_fd_sc_hd__o21ai_1 _08339_ (.A1(_02463_),
    .A2(_02464_),
    .B1(_02465_),
    .Y(_02468_));
 sky130_fd_sc_hd__inv_2 _08340_ (.A(_02468_),
    .Y(_02469_));
 sky130_fd_sc_hd__nor2_1 _08341_ (.A(_02466_),
    .B(_02469_),
    .Y(_02470_));
 sky130_fd_sc_hd__xor2_1 _08342_ (.A(_02462_),
    .B(_02470_),
    .X(_02471_));
 sky130_fd_sc_hd__o21ai_1 _08343_ (.A1(_02459_),
    .A2(_02461_),
    .B1(_02471_),
    .Y(_02472_));
 sky130_fd_sc_hd__inv_2 _08344_ (.A(_02471_),
    .Y(_02473_));
 sky130_fd_sc_hd__nand3b_1 _08345_ (.A_N(_02459_),
    .B(_02473_),
    .C(_02460_),
    .Y(_02474_));
 sky130_fd_sc_hd__nand2_1 _08346_ (.A(_02472_),
    .B(_02474_),
    .Y(_02475_));
 sky130_fd_sc_hd__nand2_1 _08347_ (.A(_04818_),
    .B(_05028_),
    .Y(_02476_));
 sky130_fd_sc_hd__nand2_1 _08348_ (.A(net40),
    .B(_03226_),
    .Y(_02477_));
 sky130_fd_sc_hd__nand2_1 _08349_ (.A(_04812_),
    .B(_03094_),
    .Y(_02479_));
 sky130_fd_sc_hd__or2_1 _08350_ (.A(_02477_),
    .B(_02479_),
    .X(_02480_));
 sky130_fd_sc_hd__nand2_1 _08351_ (.A(_02477_),
    .B(_02479_),
    .Y(_02481_));
 sky130_fd_sc_hd__nand2_1 _08352_ (.A(_02480_),
    .B(_02481_),
    .Y(_02482_));
 sky130_fd_sc_hd__or2_1 _08353_ (.A(_02476_),
    .B(_02482_),
    .X(_02483_));
 sky130_fd_sc_hd__nand2_1 _08354_ (.A(_02482_),
    .B(_02476_),
    .Y(_02484_));
 sky130_fd_sc_hd__nand2_1 _08355_ (.A(_02483_),
    .B(_02484_),
    .Y(_02485_));
 sky130_fd_sc_hd__nand2_1 _08356_ (.A(_00465_),
    .B(_00460_),
    .Y(_02486_));
 sky130_fd_sc_hd__nand2_1 _08357_ (.A(_02485_),
    .B(_02486_),
    .Y(_02487_));
 sky130_fd_sc_hd__inv_2 _08358_ (.A(_02486_),
    .Y(_02488_));
 sky130_fd_sc_hd__nand3_1 _08359_ (.A(_02488_),
    .B(_02483_),
    .C(_02484_),
    .Y(_02490_));
 sky130_fd_sc_hd__nand2_1 _08360_ (.A(_02487_),
    .B(_02490_),
    .Y(_02491_));
 sky130_fd_sc_hd__nand2_1 _08361_ (.A(_00499_),
    .B(_00494_),
    .Y(_02492_));
 sky130_fd_sc_hd__nand2_1 _08362_ (.A(_02491_),
    .B(_02492_),
    .Y(_02493_));
 sky130_fd_sc_hd__nand3b_1 _08363_ (.A_N(_02492_),
    .B(_02487_),
    .C(_02490_),
    .Y(_02494_));
 sky130_fd_sc_hd__nand2_1 _08364_ (.A(_02493_),
    .B(_02494_),
    .Y(_02495_));
 sky130_fd_sc_hd__nand2_1 _08365_ (.A(_00506_),
    .B(_00504_),
    .Y(_02496_));
 sky130_fd_sc_hd__nand2_1 _08366_ (.A(_02495_),
    .B(_02496_),
    .Y(_02497_));
 sky130_fd_sc_hd__inv_2 _08367_ (.A(_02496_),
    .Y(_02498_));
 sky130_fd_sc_hd__nand3_1 _08368_ (.A(_02498_),
    .B(_02493_),
    .C(_02494_),
    .Y(_02499_));
 sky130_fd_sc_hd__nand3_1 _08369_ (.A(_02475_),
    .B(_02497_),
    .C(_02499_),
    .Y(_02501_));
 sky130_fd_sc_hd__inv_2 _08370_ (.A(_02475_),
    .Y(_02502_));
 sky130_fd_sc_hd__nand2_1 _08371_ (.A(_02497_),
    .B(_02499_),
    .Y(_02503_));
 sky130_fd_sc_hd__nand2_1 _08372_ (.A(_02502_),
    .B(_02503_),
    .Y(_02504_));
 sky130_fd_sc_hd__nand2_1 _08373_ (.A(_02501_),
    .B(_02504_),
    .Y(_02505_));
 sky130_fd_sc_hd__or2_1 _08374_ (.A(_00477_),
    .B(_00474_),
    .X(_02506_));
 sky130_fd_sc_hd__nand2_2 _08375_ (.A(_00483_),
    .B(_02506_),
    .Y(_02507_));
 sky130_fd_sc_hd__nand2_1 _08376_ (.A(_02505_),
    .B(_02507_),
    .Y(_02508_));
 sky130_fd_sc_hd__inv_2 _08377_ (.A(_02507_),
    .Y(_02509_));
 sky130_fd_sc_hd__nand3_1 _08378_ (.A(_02501_),
    .B(_02504_),
    .C(_02509_),
    .Y(_02510_));
 sky130_fd_sc_hd__nand2_1 _08379_ (.A(_02508_),
    .B(_02510_),
    .Y(_02512_));
 sky130_fd_sc_hd__o21ai_2 _08380_ (.A1(_00512_),
    .A2(_00511_),
    .B1(_00546_),
    .Y(_02513_));
 sky130_fd_sc_hd__nand2_1 _08381_ (.A(_02512_),
    .B(_02513_),
    .Y(_02514_));
 sky130_fd_sc_hd__nand3b_1 _08382_ (.A_N(_02513_),
    .B(_02508_),
    .C(_02510_),
    .Y(_02515_));
 sky130_fd_sc_hd__nand2_1 _08383_ (.A(_02514_),
    .B(_02515_),
    .Y(_02516_));
 sky130_fd_sc_hd__inv_2 _08384_ (.A(_02516_),
    .Y(_02517_));
 sky130_fd_sc_hd__nand2_1 _08385_ (.A(_02448_),
    .B(_02517_),
    .Y(_02518_));
 sky130_fd_sc_hd__nand3_1 _08386_ (.A(_02444_),
    .B(_02447_),
    .C(_02516_),
    .Y(_02519_));
 sky130_fd_sc_hd__nand2_1 _08387_ (.A(_02518_),
    .B(_02519_),
    .Y(_02520_));
 sky130_fd_sc_hd__nand2_2 _08388_ (.A(_00568_),
    .B(_00491_),
    .Y(_02521_));
 sky130_fd_sc_hd__nand2_1 _08389_ (.A(_02520_),
    .B(_02521_),
    .Y(_02523_));
 sky130_fd_sc_hd__inv_2 _08390_ (.A(_02521_),
    .Y(_02524_));
 sky130_fd_sc_hd__nand3_1 _08391_ (.A(_02518_),
    .B(_02524_),
    .C(_02519_),
    .Y(_02525_));
 sky130_fd_sc_hd__nand2_1 _08392_ (.A(_02523_),
    .B(_02525_),
    .Y(_02526_));
 sky130_fd_sc_hd__nand2_1 _08393_ (.A(net49),
    .B(_04992_),
    .Y(_02527_));
 sky130_fd_sc_hd__o21a_1 _08394_ (.A1(_00530_),
    .A2(_00536_),
    .B1(_00534_),
    .X(_02528_));
 sky130_fd_sc_hd__nor2_1 _08395_ (.A(_02527_),
    .B(_02528_),
    .Y(_02529_));
 sky130_fd_sc_hd__inv_2 _08396_ (.A(_02529_),
    .Y(_02530_));
 sky130_fd_sc_hd__nand2_1 _08397_ (.A(_02528_),
    .B(_02527_),
    .Y(_02531_));
 sky130_fd_sc_hd__nand2_1 _08398_ (.A(_02530_),
    .B(_02531_),
    .Y(_02532_));
 sky130_fd_sc_hd__and2_1 _08399_ (.A(_00540_),
    .B(_00528_),
    .X(_02534_));
 sky130_fd_sc_hd__or2_1 _08400_ (.A(_02532_),
    .B(_02534_),
    .X(_02535_));
 sky130_fd_sc_hd__nand2_1 _08401_ (.A(_02534_),
    .B(_02532_),
    .Y(_02536_));
 sky130_fd_sc_hd__nand2_1 _08402_ (.A(_02535_),
    .B(_02536_),
    .Y(_02537_));
 sky130_fd_sc_hd__or2_1 _08403_ (.A(_00574_),
    .B(_02537_),
    .X(_02538_));
 sky130_fd_sc_hd__nand2_1 _08404_ (.A(_02537_),
    .B(_00574_),
    .Y(_02539_));
 sky130_fd_sc_hd__nand2_1 _08405_ (.A(_02538_),
    .B(_02539_),
    .Y(_02540_));
 sky130_fd_sc_hd__o21a_1 _08406_ (.A1(_00548_),
    .A2(_00551_),
    .B1(_00560_),
    .X(_02541_));
 sky130_fd_sc_hd__nor2_2 _08407_ (.A(_02540_),
    .B(_02541_),
    .Y(_02542_));
 sky130_fd_sc_hd__nand2_1 _08408_ (.A(_02541_),
    .B(_02540_),
    .Y(_02543_));
 sky130_fd_sc_hd__nor2b_1 _08409_ (.A(_02542_),
    .B_N(_02543_),
    .Y(_02545_));
 sky130_fd_sc_hd__nand2_1 _08410_ (.A(_02526_),
    .B(_02545_),
    .Y(_02546_));
 sky130_fd_sc_hd__nand3b_1 _08411_ (.A_N(_02545_),
    .B(_02523_),
    .C(_02525_),
    .Y(_02547_));
 sky130_fd_sc_hd__nand2_1 _08412_ (.A(_02546_),
    .B(_02547_),
    .Y(_02548_));
 sky130_fd_sc_hd__nand2_2 _08413_ (.A(_00586_),
    .B(_00572_),
    .Y(_02549_));
 sky130_fd_sc_hd__inv_2 _08414_ (.A(_02549_),
    .Y(_02550_));
 sky130_fd_sc_hd__nand2_1 _08415_ (.A(_02548_),
    .B(_02550_),
    .Y(_02551_));
 sky130_fd_sc_hd__nor2_1 _08416_ (.A(_02550_),
    .B(_02548_),
    .Y(_02552_));
 sky130_fd_sc_hd__a21o_1 _08417_ (.A1(_02551_),
    .A2(_00578_),
    .B1(_02552_),
    .X(_02553_));
 sky130_fd_sc_hd__a21boi_1 _08418_ (.A1(_02392_),
    .A2(_02436_),
    .B1_N(_02437_),
    .Y(_02554_));
 sky130_fd_sc_hd__nand2_1 _08419_ (.A(_01535_),
    .B(_00393_),
    .Y(_02556_));
 sky130_fd_sc_hd__nand2_1 _08420_ (.A(_00751_),
    .B(net17),
    .Y(_02557_));
 sky130_fd_sc_hd__inv_2 _08421_ (.A(_02557_),
    .Y(_02558_));
 sky130_fd_sc_hd__nand2_1 _08422_ (.A(_00795_),
    .B(net18),
    .Y(_02559_));
 sky130_fd_sc_hd__inv_2 _08423_ (.A(_02559_),
    .Y(_02560_));
 sky130_fd_sc_hd__nand2_1 _08424_ (.A(_02558_),
    .B(_02560_),
    .Y(_02561_));
 sky130_fd_sc_hd__nand2_1 _08425_ (.A(_02557_),
    .B(_02559_),
    .Y(_02562_));
 sky130_fd_sc_hd__nand2_1 _08426_ (.A(_02561_),
    .B(_02562_),
    .Y(_02563_));
 sky130_fd_sc_hd__or2_1 _08427_ (.A(_02556_),
    .B(_02563_),
    .X(_02564_));
 sky130_fd_sc_hd__nand2_1 _08428_ (.A(_02563_),
    .B(_02556_),
    .Y(_02565_));
 sky130_fd_sc_hd__nand2_1 _08429_ (.A(_02564_),
    .B(_02565_),
    .Y(_02567_));
 sky130_fd_sc_hd__a21oi_1 _08430_ (.A1(_02336_),
    .A2(_02331_),
    .B1(_02334_),
    .Y(_02568_));
 sky130_fd_sc_hd__nand2_1 _08431_ (.A(_02567_),
    .B(_02568_),
    .Y(_02569_));
 sky130_fd_sc_hd__nand3b_1 _08432_ (.A_N(_02568_),
    .B(_02564_),
    .C(_02565_),
    .Y(_02570_));
 sky130_fd_sc_hd__nand2_1 _08433_ (.A(_02569_),
    .B(_02570_),
    .Y(_02571_));
 sky130_fd_sc_hd__nand2_1 _08434_ (.A(_04260_),
    .B(_04084_),
    .Y(_02572_));
 sky130_fd_sc_hd__nand2_1 _08435_ (.A(_04293_),
    .B(_05160_),
    .Y(_02573_));
 sky130_fd_sc_hd__or2_1 _08436_ (.A(_02572_),
    .B(_02573_),
    .X(_02574_));
 sky130_fd_sc_hd__nand2_1 _08437_ (.A(_02572_),
    .B(_02573_),
    .Y(_02575_));
 sky130_fd_sc_hd__nand2_1 _08438_ (.A(_01323_),
    .B(_01565_),
    .Y(_02576_));
 sky130_fd_sc_hd__inv_2 _08439_ (.A(_02576_),
    .Y(_02578_));
 sky130_fd_sc_hd__a21o_1 _08440_ (.A1(_02574_),
    .A2(_02575_),
    .B1(_02578_),
    .X(_02579_));
 sky130_fd_sc_hd__nand3_1 _08441_ (.A(_02574_),
    .B(_02578_),
    .C(_02575_),
    .Y(_02580_));
 sky130_fd_sc_hd__nand2_1 _08442_ (.A(_02579_),
    .B(_02580_),
    .Y(_02581_));
 sky130_fd_sc_hd__nand2_1 _08443_ (.A(_02571_),
    .B(_02581_),
    .Y(_02582_));
 sky130_fd_sc_hd__inv_2 _08444_ (.A(_02581_),
    .Y(_02583_));
 sky130_fd_sc_hd__nand3_1 _08445_ (.A(_02569_),
    .B(_02583_),
    .C(_02570_),
    .Y(_02584_));
 sky130_fd_sc_hd__nand2_1 _08446_ (.A(_02582_),
    .B(_02584_),
    .Y(_02585_));
 sky130_fd_sc_hd__nand2_1 _08447_ (.A(_02359_),
    .B(_02345_),
    .Y(_02586_));
 sky130_fd_sc_hd__nand2b_1 _08448_ (.A_N(_02585_),
    .B(_02586_),
    .Y(_02587_));
 sky130_fd_sc_hd__nand3_2 _08449_ (.A(_02585_),
    .B(_02345_),
    .C(_02359_),
    .Y(_02589_));
 sky130_fd_sc_hd__nand2_1 _08450_ (.A(_02587_),
    .B(_02589_),
    .Y(_02590_));
 sky130_fd_sc_hd__nand2_1 _08451_ (.A(_00740_),
    .B(_00412_),
    .Y(_02591_));
 sky130_fd_sc_hd__nand2_1 _08452_ (.A(_00784_),
    .B(_00204_),
    .Y(_02592_));
 sky130_fd_sc_hd__or2_1 _08453_ (.A(_02591_),
    .B(_02592_),
    .X(_02593_));
 sky130_fd_sc_hd__nand2_1 _08454_ (.A(_02591_),
    .B(_02592_),
    .Y(_02594_));
 sky130_fd_sc_hd__nand2_1 _08455_ (.A(_00850_),
    .B(_00003_),
    .Y(_02595_));
 sky130_fd_sc_hd__inv_2 _08456_ (.A(_02595_),
    .Y(_02596_));
 sky130_fd_sc_hd__a21o_1 _08457_ (.A1(_02593_),
    .A2(_02594_),
    .B1(_02596_),
    .X(_02597_));
 sky130_fd_sc_hd__nand3_1 _08458_ (.A(_02593_),
    .B(_02596_),
    .C(_02594_),
    .Y(_02598_));
 sky130_fd_sc_hd__nand2_1 _08459_ (.A(_02597_),
    .B(_02598_),
    .Y(_02600_));
 sky130_fd_sc_hd__a21boi_2 _08460_ (.A1(_02349_),
    .A2(_02353_),
    .B1_N(_02352_),
    .Y(_02601_));
 sky130_fd_sc_hd__inv_2 _08461_ (.A(_02601_),
    .Y(_02602_));
 sky130_fd_sc_hd__nand2_1 _08462_ (.A(_02600_),
    .B(_02602_),
    .Y(_02603_));
 sky130_fd_sc_hd__nand3_1 _08463_ (.A(_02597_),
    .B(_02601_),
    .C(_02598_),
    .Y(_02604_));
 sky130_fd_sc_hd__nand2_1 _08464_ (.A(_02372_),
    .B(_02369_),
    .Y(_02605_));
 sky130_fd_sc_hd__inv_2 _08465_ (.A(_02605_),
    .Y(_02606_));
 sky130_fd_sc_hd__a21o_1 _08466_ (.A1(_02603_),
    .A2(_02604_),
    .B1(_02606_),
    .X(_02607_));
 sky130_fd_sc_hd__nand3_1 _08467_ (.A(_02603_),
    .B(_02606_),
    .C(_02604_),
    .Y(_02608_));
 sky130_fd_sc_hd__nand2_1 _08468_ (.A(_02607_),
    .B(_02608_),
    .Y(_02609_));
 sky130_fd_sc_hd__nand2_1 _08469_ (.A(_02590_),
    .B(_02609_),
    .Y(_02611_));
 sky130_fd_sc_hd__inv_2 _08470_ (.A(_02609_),
    .Y(_02612_));
 sky130_fd_sc_hd__nand3_2 _08471_ (.A(_02587_),
    .B(_02612_),
    .C(_02589_),
    .Y(_02613_));
 sky130_fd_sc_hd__nand2_1 _08472_ (.A(_02611_),
    .B(_02613_),
    .Y(_02614_));
 sky130_fd_sc_hd__a21o_1 _08473_ (.A1(_02386_),
    .A2(_02363_),
    .B1(_02361_),
    .X(_02615_));
 sky130_fd_sc_hd__inv_2 _08474_ (.A(_02615_),
    .Y(_02616_));
 sky130_fd_sc_hd__nand2_1 _08475_ (.A(_02614_),
    .B(_02616_),
    .Y(_02617_));
 sky130_fd_sc_hd__nand3_2 _08476_ (.A(_02615_),
    .B(_02611_),
    .C(_02613_),
    .Y(_02618_));
 sky130_fd_sc_hd__inv_2 _08477_ (.A(net8),
    .Y(_02619_));
 sky130_fd_sc_hd__nand2_1 _08478_ (.A(net7),
    .B(_02995_),
    .Y(_02620_));
 sky130_fd_sc_hd__nor3_1 _08479_ (.A(_02619_),
    .B(_01957_),
    .C(_02620_),
    .Y(_02622_));
 sky130_fd_sc_hd__inv_2 _08480_ (.A(_02622_),
    .Y(_02623_));
 sky130_fd_sc_hd__o21ai_1 _08481_ (.A1(_02619_),
    .A2(_01957_),
    .B1(_02620_),
    .Y(_02624_));
 sky130_fd_sc_hd__nand2_1 _08482_ (.A(_03215_),
    .B(_01147_),
    .Y(_02625_));
 sky130_fd_sc_hd__inv_2 _08483_ (.A(_02625_),
    .Y(_02626_));
 sky130_fd_sc_hd__a21o_1 _08484_ (.A1(_02623_),
    .A2(_02624_),
    .B1(_02626_),
    .X(_02627_));
 sky130_fd_sc_hd__nand3_1 _08485_ (.A(_02623_),
    .B(_02626_),
    .C(_02624_),
    .Y(_02628_));
 sky130_fd_sc_hd__nand2_1 _08486_ (.A(_02627_),
    .B(_02628_),
    .Y(_02629_));
 sky130_fd_sc_hd__o21a_1 _08487_ (.A1(_02398_),
    .A2(_02397_),
    .B1(_02395_),
    .X(_02630_));
 sky130_fd_sc_hd__nand2_1 _08488_ (.A(_02629_),
    .B(_02630_),
    .Y(_02631_));
 sky130_fd_sc_hd__nand2_1 _08489_ (.A(_02400_),
    .B(_02395_),
    .Y(_02633_));
 sky130_fd_sc_hd__nand3_1 _08490_ (.A(_02633_),
    .B(_02627_),
    .C(_02628_),
    .Y(_02634_));
 sky130_fd_sc_hd__nand2_1 _08491_ (.A(_02631_),
    .B(_02634_),
    .Y(_02635_));
 sky130_fd_sc_hd__nand2_1 _08492_ (.A(net38),
    .B(net3),
    .Y(_02636_));
 sky130_fd_sc_hd__inv_2 _08493_ (.A(_02636_),
    .Y(_02637_));
 sky130_fd_sc_hd__nand2_1 _08494_ (.A(_04962_),
    .B(_01873_),
    .Y(_02638_));
 sky130_fd_sc_hd__nand2_1 _08495_ (.A(_04964_),
    .B(_02544_),
    .Y(_02639_));
 sky130_fd_sc_hd__xor2_1 _08496_ (.A(_02638_),
    .B(_02639_),
    .X(_02640_));
 sky130_fd_sc_hd__or2_1 _08497_ (.A(_02637_),
    .B(_02640_),
    .X(_02641_));
 sky130_fd_sc_hd__nand2_1 _08498_ (.A(_02640_),
    .B(_02637_),
    .Y(_02642_));
 sky130_fd_sc_hd__nand2_1 _08499_ (.A(_02641_),
    .B(_02642_),
    .Y(_02644_));
 sky130_fd_sc_hd__nand2_1 _08500_ (.A(_02635_),
    .B(_02644_),
    .Y(_02645_));
 sky130_fd_sc_hd__nand3b_1 _08501_ (.A_N(_02644_),
    .B(_02631_),
    .C(_02634_),
    .Y(_02646_));
 sky130_fd_sc_hd__nand2_1 _08502_ (.A(_02645_),
    .B(_02646_),
    .Y(_02647_));
 sky130_fd_sc_hd__nand2_1 _08503_ (.A(_02374_),
    .B(_02377_),
    .Y(_02648_));
 sky130_fd_sc_hd__nor2_1 _08504_ (.A(_02377_),
    .B(_02374_),
    .Y(_02649_));
 sky130_fd_sc_hd__a21oi_2 _08505_ (.A1(_02648_),
    .A2(_02381_),
    .B1(_02649_),
    .Y(_02650_));
 sky130_fd_sc_hd__inv_2 _08506_ (.A(_02650_),
    .Y(_02651_));
 sky130_fd_sc_hd__nand2_1 _08507_ (.A(_02647_),
    .B(_02651_),
    .Y(_02652_));
 sky130_fd_sc_hd__nand3_1 _08508_ (.A(_02645_),
    .B(_02646_),
    .C(_02650_),
    .Y(_02653_));
 sky130_fd_sc_hd__nand2_1 _08509_ (.A(_02652_),
    .B(_02653_),
    .Y(_02655_));
 sky130_fd_sc_hd__or2_1 _08510_ (.A(_02406_),
    .B(_02403_),
    .X(_02656_));
 sky130_fd_sc_hd__nand2_1 _08511_ (.A(_02419_),
    .B(_02656_),
    .Y(_02657_));
 sky130_fd_sc_hd__nand2_1 _08512_ (.A(_02655_),
    .B(_02657_),
    .Y(_02658_));
 sky130_fd_sc_hd__nand3b_1 _08513_ (.A_N(_02657_),
    .B(_02652_),
    .C(_02653_),
    .Y(_02659_));
 sky130_fd_sc_hd__nand2_1 _08514_ (.A(_02658_),
    .B(_02659_),
    .Y(_02660_));
 sky130_fd_sc_hd__inv_2 _08515_ (.A(_02660_),
    .Y(_02661_));
 sky130_fd_sc_hd__nand3_1 _08516_ (.A(_02617_),
    .B(_02618_),
    .C(_02661_),
    .Y(_02662_));
 sky130_fd_sc_hd__nand2_1 _08517_ (.A(_02617_),
    .B(_02618_),
    .Y(_02663_));
 sky130_fd_sc_hd__nand2_1 _08518_ (.A(_02663_),
    .B(_02660_),
    .Y(_02664_));
 sky130_fd_sc_hd__nand3_1 _08519_ (.A(_02554_),
    .B(_02662_),
    .C(_02664_),
    .Y(_02666_));
 sky130_fd_sc_hd__nand2_1 _08520_ (.A(_02664_),
    .B(_02662_),
    .Y(_02667_));
 sky130_fd_sc_hd__nand2_1 _08521_ (.A(_02438_),
    .B(_02437_),
    .Y(_02668_));
 sky130_fd_sc_hd__nand2_1 _08522_ (.A(_02667_),
    .B(_02668_),
    .Y(_02669_));
 sky130_fd_sc_hd__nand2_1 _08523_ (.A(_02666_),
    .B(_02669_),
    .Y(_02670_));
 sky130_fd_sc_hd__nand2_1 _08524_ (.A(net40),
    .B(_03094_),
    .Y(_02671_));
 sky130_fd_sc_hd__nand2_1 _08525_ (.A(_04812_),
    .B(_02753_),
    .Y(_02672_));
 sky130_fd_sc_hd__or2_1 _08526_ (.A(_02671_),
    .B(_02672_),
    .X(_02673_));
 sky130_fd_sc_hd__nand2_1 _08527_ (.A(_02671_),
    .B(_02672_),
    .Y(_02674_));
 sky130_fd_sc_hd__nand2_1 _08528_ (.A(_04818_),
    .B(_03226_),
    .Y(_02675_));
 sky130_fd_sc_hd__inv_2 _08529_ (.A(_02675_),
    .Y(_02677_));
 sky130_fd_sc_hd__a21o_1 _08530_ (.A1(_02673_),
    .A2(_02674_),
    .B1(_02677_),
    .X(_02678_));
 sky130_fd_sc_hd__nand3_2 _08531_ (.A(_02673_),
    .B(_02677_),
    .C(_02674_),
    .Y(_02679_));
 sky130_fd_sc_hd__inv_2 _08532_ (.A(_02409_),
    .Y(_02680_));
 sky130_fd_sc_hd__a21oi_2 _08533_ (.A1(_02415_),
    .A2(_02680_),
    .B1(_02413_),
    .Y(_02681_));
 sky130_fd_sc_hd__a21o_1 _08534_ (.A1(_02678_),
    .A2(_02679_),
    .B1(_02681_),
    .X(_02682_));
 sky130_fd_sc_hd__nand3_1 _08535_ (.A(_02678_),
    .B(_02681_),
    .C(_02679_),
    .Y(_02683_));
 sky130_fd_sc_hd__nand2_1 _08536_ (.A(_02682_),
    .B(_02683_),
    .Y(_02684_));
 sky130_fd_sc_hd__nand2_2 _08537_ (.A(_02483_),
    .B(_02480_),
    .Y(_02685_));
 sky130_fd_sc_hd__nand2_1 _08538_ (.A(_02684_),
    .B(_02685_),
    .Y(_02686_));
 sky130_fd_sc_hd__inv_2 _08539_ (.A(_02685_),
    .Y(_02688_));
 sky130_fd_sc_hd__nand3_1 _08540_ (.A(_02682_),
    .B(_02683_),
    .C(_02688_),
    .Y(_02689_));
 sky130_fd_sc_hd__nand2_1 _08541_ (.A(_02686_),
    .B(_02689_),
    .Y(_02690_));
 sky130_fd_sc_hd__nand2_1 _08542_ (.A(_02485_),
    .B(_02488_),
    .Y(_02691_));
 sky130_fd_sc_hd__nor2_1 _08543_ (.A(_02488_),
    .B(_02485_),
    .Y(_02692_));
 sky130_fd_sc_hd__a21oi_2 _08544_ (.A1(_02691_),
    .A2(_02492_),
    .B1(_02692_),
    .Y(_02693_));
 sky130_fd_sc_hd__inv_2 _08545_ (.A(_02693_),
    .Y(_02694_));
 sky130_fd_sc_hd__nand2_1 _08546_ (.A(_02690_),
    .B(_02694_),
    .Y(_02695_));
 sky130_fd_sc_hd__nand3_1 _08547_ (.A(_02686_),
    .B(_02693_),
    .C(_02689_),
    .Y(_02696_));
 sky130_fd_sc_hd__nand2_1 _08548_ (.A(_02695_),
    .B(_02696_),
    .Y(_02697_));
 sky130_fd_sc_hd__inv_2 _08549_ (.A(_03314_),
    .Y(_02699_));
 sky130_fd_sc_hd__nand2_1 _08550_ (.A(net43),
    .B(_03402_),
    .Y(_02700_));
 sky130_fd_sc_hd__nor3_1 _08551_ (.A(_00110_),
    .B(_02699_),
    .C(_02700_),
    .Y(_02701_));
 sky130_fd_sc_hd__o21ai_2 _08552_ (.A1(_00110_),
    .A2(_02699_),
    .B1(_02700_),
    .Y(_02702_));
 sky130_fd_sc_hd__inv_2 _08553_ (.A(_02702_),
    .Y(_02703_));
 sky130_fd_sc_hd__nand2_1 _08554_ (.A(_04876_),
    .B(_03820_),
    .Y(_02704_));
 sky130_fd_sc_hd__o21ai_1 _08555_ (.A1(_02701_),
    .A2(_02703_),
    .B1(_02704_),
    .Y(_02705_));
 sky130_fd_sc_hd__inv_2 _08556_ (.A(_02704_),
    .Y(_02706_));
 sky130_fd_sc_hd__nand3b_1 _08557_ (.A_N(_02701_),
    .B(_02706_),
    .C(_02702_),
    .Y(_02707_));
 sky130_fd_sc_hd__nand2_1 _08558_ (.A(_02705_),
    .B(_02707_),
    .Y(_02708_));
 sky130_fd_sc_hd__inv_2 _08559_ (.A(_02450_),
    .Y(_02710_));
 sky130_fd_sc_hd__a21oi_1 _08560_ (.A1(_02454_),
    .A2(_02710_),
    .B1(_02453_),
    .Y(_02711_));
 sky130_fd_sc_hd__inv_2 _08561_ (.A(_02711_),
    .Y(_02712_));
 sky130_fd_sc_hd__nand2b_1 _08562_ (.A_N(_02708_),
    .B(_02712_),
    .Y(_02713_));
 sky130_fd_sc_hd__nand2_1 _08563_ (.A(_02708_),
    .B(_02711_),
    .Y(_02714_));
 sky130_fd_sc_hd__nand2_1 _08564_ (.A(_02713_),
    .B(_02714_),
    .Y(_02715_));
 sky130_fd_sc_hd__nand2_1 _08565_ (.A(_00529_),
    .B(_04828_),
    .Y(_02716_));
 sky130_fd_sc_hd__nand2_1 _08566_ (.A(_00124_),
    .B(_04819_),
    .Y(_02717_));
 sky130_fd_sc_hd__nor3_1 _08567_ (.A(_02463_),
    .B(_00111_),
    .C(_02717_),
    .Y(_02718_));
 sky130_fd_sc_hd__o21ai_1 _08568_ (.A1(_02463_),
    .A2(_00111_),
    .B1(_02717_),
    .Y(_02719_));
 sky130_fd_sc_hd__nand2b_1 _08569_ (.A_N(_02718_),
    .B(_02719_),
    .Y(_02721_));
 sky130_fd_sc_hd__or2_1 _08570_ (.A(_02716_),
    .B(_02721_),
    .X(_02722_));
 sky130_fd_sc_hd__nand2_1 _08571_ (.A(_02721_),
    .B(_02716_),
    .Y(_02723_));
 sky130_fd_sc_hd__nand2_1 _08572_ (.A(_02722_),
    .B(_02723_),
    .Y(_02724_));
 sky130_fd_sc_hd__nand2_1 _08573_ (.A(_02715_),
    .B(_02724_),
    .Y(_02725_));
 sky130_fd_sc_hd__inv_2 _08574_ (.A(_02724_),
    .Y(_02726_));
 sky130_fd_sc_hd__nand3_1 _08575_ (.A(_02726_),
    .B(_02713_),
    .C(_02714_),
    .Y(_02727_));
 sky130_fd_sc_hd__nand2_1 _08576_ (.A(_02725_),
    .B(_02727_),
    .Y(_02728_));
 sky130_fd_sc_hd__inv_2 _08577_ (.A(_02728_),
    .Y(_02729_));
 sky130_fd_sc_hd__nand2_1 _08578_ (.A(_02697_),
    .B(_02729_),
    .Y(_02730_));
 sky130_fd_sc_hd__nand3_1 _08579_ (.A(_02695_),
    .B(_02696_),
    .C(_02728_),
    .Y(_02732_));
 sky130_fd_sc_hd__nand2_1 _08580_ (.A(_02730_),
    .B(_02732_),
    .Y(_02733_));
 sky130_fd_sc_hd__nand2_1 _08581_ (.A(_02422_),
    .B(_02426_),
    .Y(_02734_));
 sky130_fd_sc_hd__nor2_1 _08582_ (.A(_02426_),
    .B(_02422_),
    .Y(_02735_));
 sky130_fd_sc_hd__a21oi_2 _08583_ (.A1(_02734_),
    .A2(_02431_),
    .B1(_02735_),
    .Y(_02736_));
 sky130_fd_sc_hd__inv_2 _08584_ (.A(_02736_),
    .Y(_02737_));
 sky130_fd_sc_hd__nand2_1 _08585_ (.A(_02733_),
    .B(_02737_),
    .Y(_02738_));
 sky130_fd_sc_hd__nand3_1 _08586_ (.A(_02736_),
    .B(_02730_),
    .C(_02732_),
    .Y(_02739_));
 sky130_fd_sc_hd__nand2_1 _08587_ (.A(_02738_),
    .B(_02739_),
    .Y(_02740_));
 sky130_fd_sc_hd__o21ai_2 _08588_ (.A1(_02498_),
    .A2(_02495_),
    .B1(_02504_),
    .Y(_02741_));
 sky130_fd_sc_hd__nand2_1 _08589_ (.A(_02740_),
    .B(_02741_),
    .Y(_02743_));
 sky130_fd_sc_hd__nand3b_1 _08590_ (.A_N(_02741_),
    .B(_02738_),
    .C(_02739_),
    .Y(_02744_));
 sky130_fd_sc_hd__nand2_1 _08591_ (.A(_02743_),
    .B(_02744_),
    .Y(_02745_));
 sky130_fd_sc_hd__inv_2 _08592_ (.A(_02745_),
    .Y(_02746_));
 sky130_fd_sc_hd__nand2_1 _08593_ (.A(_02670_),
    .B(_02746_),
    .Y(_02747_));
 sky130_fd_sc_hd__nand3_2 _08594_ (.A(_02666_),
    .B(_02669_),
    .C(_02745_),
    .Y(_02748_));
 sky130_fd_sc_hd__nand2_1 _08595_ (.A(_02747_),
    .B(_02748_),
    .Y(_02749_));
 sky130_fd_sc_hd__nand2_1 _08596_ (.A(_02442_),
    .B(_02446_),
    .Y(_02750_));
 sky130_fd_sc_hd__nor2_1 _08597_ (.A(_02446_),
    .B(_02442_),
    .Y(_02751_));
 sky130_fd_sc_hd__a21oi_4 _08598_ (.A1(_02750_),
    .A2(_02517_),
    .B1(_02751_),
    .Y(_02752_));
 sky130_fd_sc_hd__inv_2 _08599_ (.A(_02752_),
    .Y(_02754_));
 sky130_fd_sc_hd__nand2_1 _08600_ (.A(_02749_),
    .B(_02754_),
    .Y(_02755_));
 sky130_fd_sc_hd__nand3_1 _08601_ (.A(_02752_),
    .B(_02747_),
    .C(_02748_),
    .Y(_02756_));
 sky130_fd_sc_hd__nand2_1 _08602_ (.A(_02755_),
    .B(_02756_),
    .Y(_02757_));
 sky130_fd_sc_hd__nand2_1 _08603_ (.A(_02505_),
    .B(_02509_),
    .Y(_02758_));
 sky130_fd_sc_hd__nor2_1 _08604_ (.A(_02509_),
    .B(_02505_),
    .Y(_02759_));
 sky130_fd_sc_hd__a21oi_2 _08605_ (.A1(_02758_),
    .A2(_02513_),
    .B1(_02759_),
    .Y(_02760_));
 sky130_fd_sc_hd__inv_2 _08606_ (.A(_02760_),
    .Y(_02761_));
 sky130_fd_sc_hd__and4_1 _08607_ (.A(net49),
    .B(net50),
    .C(_04911_),
    .D(_04895_),
    .X(_02762_));
 sky130_fd_sc_hd__inv_2 _08608_ (.A(_02762_),
    .Y(_02763_));
 sky130_fd_sc_hd__a22o_1 _08609_ (.A1(net49),
    .A2(_04991_),
    .B1(net50),
    .B2(_04895_),
    .X(_02765_));
 sky130_fd_sc_hd__nand2_1 _08610_ (.A(_02763_),
    .B(_02765_),
    .Y(_02766_));
 sky130_fd_sc_hd__o21ba_1 _08611_ (.A1(_02462_),
    .A2(_02469_),
    .B1_N(_02466_),
    .X(_02767_));
 sky130_fd_sc_hd__nor2_1 _08612_ (.A(_02766_),
    .B(_02767_),
    .Y(_02768_));
 sky130_fd_sc_hd__inv_2 _08613_ (.A(_02768_),
    .Y(_02769_));
 sky130_fd_sc_hd__nand2_1 _08614_ (.A(_02767_),
    .B(_02766_),
    .Y(_02770_));
 sky130_fd_sc_hd__nand2_1 _08615_ (.A(_02769_),
    .B(_02770_),
    .Y(_02771_));
 sky130_fd_sc_hd__a21oi_1 _08616_ (.A1(_02460_),
    .A2(_02473_),
    .B1(_02459_),
    .Y(_02772_));
 sky130_fd_sc_hd__or2_1 _08617_ (.A(_02771_),
    .B(_02772_),
    .X(_02773_));
 sky130_fd_sc_hd__nand2_1 _08618_ (.A(_02772_),
    .B(_02771_),
    .Y(_02774_));
 sky130_fd_sc_hd__nand2_1 _08619_ (.A(_02773_),
    .B(_02774_),
    .Y(_02776_));
 sky130_fd_sc_hd__nand2_1 _08620_ (.A(_02776_),
    .B(_02530_),
    .Y(_02777_));
 sky130_fd_sc_hd__nand3_2 _08621_ (.A(_02773_),
    .B(_02529_),
    .C(_02774_),
    .Y(_02778_));
 sky130_fd_sc_hd__nand2_1 _08622_ (.A(_02777_),
    .B(_02778_),
    .Y(_02779_));
 sky130_fd_sc_hd__nand2_1 _08623_ (.A(_02779_),
    .B(_02535_),
    .Y(_02780_));
 sky130_fd_sc_hd__nand3b_2 _08624_ (.A_N(_02535_),
    .B(_02777_),
    .C(_02778_),
    .Y(_02781_));
 sky130_fd_sc_hd__nand2_1 _08625_ (.A(_02780_),
    .B(_02781_),
    .Y(_02782_));
 sky130_fd_sc_hd__inv_2 _08626_ (.A(_02782_),
    .Y(_02783_));
 sky130_fd_sc_hd__nand2_1 _08627_ (.A(_02761_),
    .B(_02783_),
    .Y(_02784_));
 sky130_fd_sc_hd__nand2_1 _08628_ (.A(_02760_),
    .B(_02782_),
    .Y(_02785_));
 sky130_fd_sc_hd__nand2_1 _08629_ (.A(_02784_),
    .B(_02785_),
    .Y(_02787_));
 sky130_fd_sc_hd__nand2_1 _08630_ (.A(_02787_),
    .B(_02538_),
    .Y(_02788_));
 sky130_fd_sc_hd__nand3b_1 _08631_ (.A_N(_02538_),
    .B(_02784_),
    .C(_02785_),
    .Y(_02789_));
 sky130_fd_sc_hd__nand2_1 _08632_ (.A(_02788_),
    .B(_02789_),
    .Y(_02790_));
 sky130_fd_sc_hd__inv_2 _08633_ (.A(_02790_),
    .Y(_02791_));
 sky130_fd_sc_hd__nand2_1 _08634_ (.A(_02757_),
    .B(_02791_),
    .Y(_02792_));
 sky130_fd_sc_hd__nand3_1 _08635_ (.A(_02755_),
    .B(_02756_),
    .C(_02790_),
    .Y(_02793_));
 sky130_fd_sc_hd__nand2_1 _08636_ (.A(_02792_),
    .B(_02793_),
    .Y(_02794_));
 sky130_fd_sc_hd__nand2_1 _08637_ (.A(_02520_),
    .B(_02524_),
    .Y(_02795_));
 sky130_fd_sc_hd__nor2_1 _08638_ (.A(_02524_),
    .B(_02520_),
    .Y(_02796_));
 sky130_fd_sc_hd__a21oi_2 _08639_ (.A1(_02795_),
    .A2(_02545_),
    .B1(_02796_),
    .Y(_02798_));
 sky130_fd_sc_hd__inv_2 _08640_ (.A(_02798_),
    .Y(_02799_));
 sky130_fd_sc_hd__nand2_1 _08641_ (.A(_02794_),
    .B(_02799_),
    .Y(_02800_));
 sky130_fd_sc_hd__nand3_1 _08642_ (.A(_02798_),
    .B(_02792_),
    .C(_02793_),
    .Y(_02801_));
 sky130_fd_sc_hd__nand2_1 _08643_ (.A(_02800_),
    .B(_02801_),
    .Y(_02802_));
 sky130_fd_sc_hd__nand2_1 _08644_ (.A(_02802_),
    .B(_02542_),
    .Y(_02803_));
 sky130_fd_sc_hd__nand3b_1 _08645_ (.A_N(_02542_),
    .B(_02800_),
    .C(_02801_),
    .Y(_02804_));
 sky130_fd_sc_hd__nand3_1 _08646_ (.A(_02553_),
    .B(_02803_),
    .C(_02804_),
    .Y(_02805_));
 sky130_fd_sc_hd__nand2_1 _08647_ (.A(_02803_),
    .B(_02804_),
    .Y(_02806_));
 sky130_fd_sc_hd__a21oi_2 _08648_ (.A1(_02551_),
    .A2(_00578_),
    .B1(_02552_),
    .Y(_02807_));
 sky130_fd_sc_hd__nand2_1 _08649_ (.A(_02806_),
    .B(_02807_),
    .Y(_02809_));
 sky130_fd_sc_hd__nand2_1 _08650_ (.A(_02805_),
    .B(_02809_),
    .Y(_02810_));
 sky130_fd_sc_hd__nand2_1 _08651_ (.A(_02548_),
    .B(_02549_),
    .Y(_02811_));
 sky130_fd_sc_hd__nand3_1 _08652_ (.A(_02546_),
    .B(_02547_),
    .C(_02550_),
    .Y(_02812_));
 sky130_fd_sc_hd__nand2_1 _08653_ (.A(_02811_),
    .B(_02812_),
    .Y(_02813_));
 sky130_fd_sc_hd__nand2_1 _08654_ (.A(_02813_),
    .B(_00578_),
    .Y(_02814_));
 sky130_fd_sc_hd__or2_1 _08655_ (.A(_00371_),
    .B(_00591_),
    .X(_02815_));
 sky130_fd_sc_hd__nand2_2 _08656_ (.A(_00605_),
    .B(_02815_),
    .Y(_02816_));
 sky130_fd_sc_hd__nand3_1 _08657_ (.A(_02811_),
    .B(_02812_),
    .C(_00579_),
    .Y(_02817_));
 sky130_fd_sc_hd__nand3_2 _08658_ (.A(_02814_),
    .B(_02816_),
    .C(_02817_),
    .Y(_02818_));
 sky130_fd_sc_hd__nand2_1 _08659_ (.A(_02810_),
    .B(_02818_),
    .Y(_02820_));
 sky130_fd_sc_hd__nand3b_1 _08660_ (.A_N(_02818_),
    .B(_02805_),
    .C(_02809_),
    .Y(_02821_));
 sky130_fd_sc_hd__nand2_1 _08661_ (.A(_02820_),
    .B(_02821_),
    .Y(_02822_));
 sky130_fd_sc_hd__inv_2 _08662_ (.A(_02822_),
    .Y(_02823_));
 sky130_fd_sc_hd__nand2_1 _08663_ (.A(_02814_),
    .B(_02817_),
    .Y(_02824_));
 sky130_fd_sc_hd__inv_2 _08664_ (.A(_02816_),
    .Y(_02825_));
 sky130_fd_sc_hd__nand2_1 _08665_ (.A(_02824_),
    .B(_02825_),
    .Y(_02826_));
 sky130_fd_sc_hd__nand2_1 _08666_ (.A(_02826_),
    .B(_02818_),
    .Y(_02827_));
 sky130_fd_sc_hd__nand2_1 _08667_ (.A(_02827_),
    .B(_00602_),
    .Y(_02828_));
 sky130_fd_sc_hd__nand3b_1 _08668_ (.A_N(_00602_),
    .B(_02826_),
    .C(_02818_),
    .Y(_02829_));
 sky130_fd_sc_hd__nand2_1 _08669_ (.A(_02828_),
    .B(_02829_),
    .Y(_02831_));
 sky130_fd_sc_hd__inv_2 _08670_ (.A(_02831_),
    .Y(_02832_));
 sky130_fd_sc_hd__nand2_1 _08671_ (.A(_02823_),
    .B(_02832_),
    .Y(_02833_));
 sky130_fd_sc_hd__nand2_1 _08672_ (.A(_02662_),
    .B(_02618_),
    .Y(_02834_));
 sky130_fd_sc_hd__nand2_1 _08673_ (.A(_02613_),
    .B(_02587_),
    .Y(_02835_));
 sky130_fd_sc_hd__nand2_1 _08674_ (.A(_02564_),
    .B(_02561_),
    .Y(_02836_));
 sky130_fd_sc_hd__nand2_1 _08675_ (.A(_02357_),
    .B(net18),
    .Y(_02837_));
 sky130_fd_sc_hd__nand2_1 _08676_ (.A(_02379_),
    .B(net19),
    .Y(_02838_));
 sky130_fd_sc_hd__or2_1 _08677_ (.A(_02837_),
    .B(_02838_),
    .X(_02839_));
 sky130_fd_sc_hd__nand2_1 _08678_ (.A(_02837_),
    .B(_02838_),
    .Y(_02840_));
 sky130_fd_sc_hd__nand2_1 _08679_ (.A(_01535_),
    .B(net17),
    .Y(_02842_));
 sky130_fd_sc_hd__inv_2 _08680_ (.A(_02842_),
    .Y(_02843_));
 sky130_fd_sc_hd__a21o_1 _08681_ (.A1(_02839_),
    .A2(_02840_),
    .B1(_02843_),
    .X(_02844_));
 sky130_fd_sc_hd__nand3_1 _08682_ (.A(_02839_),
    .B(_02843_),
    .C(_02840_),
    .Y(_02845_));
 sky130_fd_sc_hd__nand3_1 _08683_ (.A(_02836_),
    .B(_02844_),
    .C(_02845_),
    .Y(_02846_));
 sky130_fd_sc_hd__nand2_1 _08684_ (.A(_02844_),
    .B(_02845_),
    .Y(_02847_));
 sky130_fd_sc_hd__o21a_1 _08685_ (.A1(_02556_),
    .A2(_02563_),
    .B1(_02561_),
    .X(_02848_));
 sky130_fd_sc_hd__nand2_1 _08686_ (.A(_02847_),
    .B(_02848_),
    .Y(_02849_));
 sky130_fd_sc_hd__nand2_1 _08687_ (.A(_02846_),
    .B(_02849_),
    .Y(_02850_));
 sky130_fd_sc_hd__nand2_1 _08688_ (.A(_01048_),
    .B(_05160_),
    .Y(_02851_));
 sky130_fd_sc_hd__nand2_1 _08689_ (.A(_01092_),
    .B(_00393_),
    .Y(_02853_));
 sky130_fd_sc_hd__or2_1 _08690_ (.A(_02851_),
    .B(_02853_),
    .X(_02854_));
 sky130_fd_sc_hd__nand2_1 _08691_ (.A(_02851_),
    .B(_02853_),
    .Y(_02855_));
 sky130_fd_sc_hd__nand2_1 _08692_ (.A(_01565_),
    .B(_04084_),
    .Y(_02856_));
 sky130_fd_sc_hd__inv_2 _08693_ (.A(_02856_),
    .Y(_02857_));
 sky130_fd_sc_hd__a21o_1 _08694_ (.A1(_02854_),
    .A2(_02855_),
    .B1(_02857_),
    .X(_02858_));
 sky130_fd_sc_hd__nand3_1 _08695_ (.A(_02854_),
    .B(_02857_),
    .C(_02855_),
    .Y(_02859_));
 sky130_fd_sc_hd__nand2_1 _08696_ (.A(_02858_),
    .B(_02859_),
    .Y(_02860_));
 sky130_fd_sc_hd__nand2_1 _08697_ (.A(_02850_),
    .B(_02860_),
    .Y(_02861_));
 sky130_fd_sc_hd__nand3b_1 _08698_ (.A_N(_02860_),
    .B(_02846_),
    .C(_02849_),
    .Y(_02862_));
 sky130_fd_sc_hd__nand2_1 _08699_ (.A(_02861_),
    .B(_02862_),
    .Y(_02864_));
 sky130_fd_sc_hd__nand2_1 _08700_ (.A(_02584_),
    .B(_02570_),
    .Y(_02865_));
 sky130_fd_sc_hd__inv_2 _08701_ (.A(_02865_),
    .Y(_02866_));
 sky130_fd_sc_hd__nand2_1 _08702_ (.A(_02864_),
    .B(_02866_),
    .Y(_02867_));
 sky130_fd_sc_hd__nand3_1 _08703_ (.A(_02865_),
    .B(_02861_),
    .C(_02862_),
    .Y(_02868_));
 sky130_fd_sc_hd__nand2_1 _08704_ (.A(_02867_),
    .B(_02868_),
    .Y(_02869_));
 sky130_fd_sc_hd__inv_2 _08705_ (.A(_01323_),
    .Y(_02870_));
 sky130_fd_sc_hd__nand2_1 _08706_ (.A(_00784_),
    .B(_00412_),
    .Y(_02871_));
 sky130_fd_sc_hd__or3_1 _08707_ (.A(_02870_),
    .B(_01937_),
    .C(_02871_),
    .X(_02872_));
 sky130_fd_sc_hd__o21ai_1 _08708_ (.A1(_02870_),
    .A2(_01937_),
    .B1(_02871_),
    .Y(_02873_));
 sky130_fd_sc_hd__nand2_1 _08709_ (.A(_02872_),
    .B(_02873_),
    .Y(_02875_));
 sky130_fd_sc_hd__nand2_1 _08710_ (.A(_00740_),
    .B(_00003_),
    .Y(_02876_));
 sky130_fd_sc_hd__nand2_1 _08711_ (.A(_02875_),
    .B(_02876_),
    .Y(_02877_));
 sky130_fd_sc_hd__nand3b_1 _08712_ (.A_N(_02876_),
    .B(_02872_),
    .C(_02873_),
    .Y(_02878_));
 sky130_fd_sc_hd__nand2_1 _08713_ (.A(_02877_),
    .B(_02878_),
    .Y(_02879_));
 sky130_fd_sc_hd__nand2_1 _08714_ (.A(_02580_),
    .B(_02574_),
    .Y(_02880_));
 sky130_fd_sc_hd__nand2_1 _08715_ (.A(_02879_),
    .B(_02880_),
    .Y(_02881_));
 sky130_fd_sc_hd__inv_2 _08716_ (.A(_02880_),
    .Y(_02882_));
 sky130_fd_sc_hd__nand3_1 _08717_ (.A(_02877_),
    .B(_02878_),
    .C(_02882_),
    .Y(_02883_));
 sky130_fd_sc_hd__nand2_1 _08718_ (.A(_02881_),
    .B(_02883_),
    .Y(_02884_));
 sky130_fd_sc_hd__nand2_1 _08719_ (.A(_02598_),
    .B(_02593_),
    .Y(_02886_));
 sky130_fd_sc_hd__nand2_1 _08720_ (.A(_02884_),
    .B(_02886_),
    .Y(_02887_));
 sky130_fd_sc_hd__nand3b_1 _08721_ (.A_N(_02886_),
    .B(_02881_),
    .C(_02883_),
    .Y(_02888_));
 sky130_fd_sc_hd__nand2_1 _08722_ (.A(_02887_),
    .B(_02888_),
    .Y(_02889_));
 sky130_fd_sc_hd__nand2_1 _08723_ (.A(_02869_),
    .B(_02889_),
    .Y(_02890_));
 sky130_fd_sc_hd__inv_2 _08724_ (.A(_02889_),
    .Y(_02891_));
 sky130_fd_sc_hd__nand3_2 _08725_ (.A(_02891_),
    .B(_02868_),
    .C(_02867_),
    .Y(_02892_));
 sky130_fd_sc_hd__nand3_2 _08726_ (.A(_02835_),
    .B(_02890_),
    .C(_02892_),
    .Y(_02893_));
 sky130_fd_sc_hd__inv_2 _08727_ (.A(net9),
    .Y(_02894_));
 sky130_fd_sc_hd__nand2_1 _08728_ (.A(_01081_),
    .B(_02995_),
    .Y(_02895_));
 sky130_fd_sc_hd__nor3_1 _08729_ (.A(_02894_),
    .B(_01957_),
    .C(_02895_),
    .Y(_02897_));
 sky130_fd_sc_hd__inv_2 _08730_ (.A(_02897_),
    .Y(_02898_));
 sky130_fd_sc_hd__o21ai_1 _08731_ (.A1(_02894_),
    .A2(_01957_),
    .B1(_02895_),
    .Y(_02899_));
 sky130_fd_sc_hd__nand2_1 _08732_ (.A(_03215_),
    .B(_01037_),
    .Y(_02900_));
 sky130_fd_sc_hd__inv_2 _08733_ (.A(_02900_),
    .Y(_02901_));
 sky130_fd_sc_hd__a21o_1 _08734_ (.A1(_02898_),
    .A2(_02899_),
    .B1(_02901_),
    .X(_02902_));
 sky130_fd_sc_hd__nand3_1 _08735_ (.A(_02898_),
    .B(_02901_),
    .C(_02899_),
    .Y(_02903_));
 sky130_fd_sc_hd__nand2_1 _08736_ (.A(_02902_),
    .B(_02903_),
    .Y(_02904_));
 sky130_fd_sc_hd__nand2_1 _08737_ (.A(_02628_),
    .B(_02623_),
    .Y(_02905_));
 sky130_fd_sc_hd__nand2_1 _08738_ (.A(_02904_),
    .B(_02905_),
    .Y(_02906_));
 sky130_fd_sc_hd__inv_2 _08739_ (.A(_02905_),
    .Y(_02908_));
 sky130_fd_sc_hd__nand3_1 _08740_ (.A(_02908_),
    .B(_02902_),
    .C(_02903_),
    .Y(_02909_));
 sky130_fd_sc_hd__nand2_1 _08741_ (.A(_02906_),
    .B(_02909_),
    .Y(_02910_));
 sky130_fd_sc_hd__nand2_1 _08742_ (.A(_03809_),
    .B(_01873_),
    .Y(_02911_));
 sky130_fd_sc_hd__inv_2 _08743_ (.A(_02911_),
    .Y(_02912_));
 sky130_fd_sc_hd__inv_2 _08744_ (.A(net6),
    .Y(_02913_));
 sky130_fd_sc_hd__nand2_1 _08745_ (.A(net37),
    .B(net5),
    .Y(_02914_));
 sky130_fd_sc_hd__nor3_1 _08746_ (.A(_01330_),
    .B(_02913_),
    .C(_02914_),
    .Y(_02915_));
 sky130_fd_sc_hd__o21ai_1 _08747_ (.A1(_01330_),
    .A2(_02913_),
    .B1(_02914_),
    .Y(_02916_));
 sky130_fd_sc_hd__nor2b_1 _08748_ (.A(_02915_),
    .B_N(_02916_),
    .Y(_02917_));
 sky130_fd_sc_hd__or2_1 _08749_ (.A(_02912_),
    .B(_02917_),
    .X(_02919_));
 sky130_fd_sc_hd__nand2_1 _08750_ (.A(_02917_),
    .B(_02912_),
    .Y(_02920_));
 sky130_fd_sc_hd__nand2_1 _08751_ (.A(_02919_),
    .B(_02920_),
    .Y(_02921_));
 sky130_fd_sc_hd__inv_2 _08752_ (.A(_02921_),
    .Y(_02922_));
 sky130_fd_sc_hd__nand2_1 _08753_ (.A(_02910_),
    .B(_02922_),
    .Y(_02923_));
 sky130_fd_sc_hd__nand3_1 _08754_ (.A(_02906_),
    .B(_02909_),
    .C(_02921_),
    .Y(_02924_));
 sky130_fd_sc_hd__nand2_1 _08755_ (.A(_02923_),
    .B(_02924_),
    .Y(_02925_));
 sky130_fd_sc_hd__nand2_1 _08756_ (.A(_02600_),
    .B(_02601_),
    .Y(_02926_));
 sky130_fd_sc_hd__nor2_1 _08757_ (.A(_02601_),
    .B(_02600_),
    .Y(_02927_));
 sky130_fd_sc_hd__a21oi_2 _08758_ (.A1(_02926_),
    .A2(_02605_),
    .B1(_02927_),
    .Y(_02928_));
 sky130_fd_sc_hd__inv_2 _08759_ (.A(_02928_),
    .Y(_02930_));
 sky130_fd_sc_hd__nand2_1 _08760_ (.A(_02925_),
    .B(_02930_),
    .Y(_02931_));
 sky130_fd_sc_hd__nand3_1 _08761_ (.A(_02923_),
    .B(_02924_),
    .C(_02928_),
    .Y(_02932_));
 sky130_fd_sc_hd__nand2_1 _08762_ (.A(_02931_),
    .B(_02932_),
    .Y(_02933_));
 sky130_fd_sc_hd__nand2_1 _08763_ (.A(_02646_),
    .B(_02634_),
    .Y(_02934_));
 sky130_fd_sc_hd__nand2_1 _08764_ (.A(_02933_),
    .B(_02934_),
    .Y(_02935_));
 sky130_fd_sc_hd__nand3b_1 _08765_ (.A_N(_02934_),
    .B(_02931_),
    .C(_02932_),
    .Y(_02936_));
 sky130_fd_sc_hd__nand2_1 _08766_ (.A(_02935_),
    .B(_02936_),
    .Y(_02937_));
 sky130_fd_sc_hd__inv_2 _08767_ (.A(_02937_),
    .Y(_02938_));
 sky130_fd_sc_hd__a21boi_1 _08768_ (.A1(_02612_),
    .A2(_02589_),
    .B1_N(_02587_),
    .Y(_02939_));
 sky130_fd_sc_hd__nand2_1 _08769_ (.A(_02892_),
    .B(_02890_),
    .Y(_02941_));
 sky130_fd_sc_hd__nand2_1 _08770_ (.A(_02939_),
    .B(_02941_),
    .Y(_02942_));
 sky130_fd_sc_hd__nand3_2 _08771_ (.A(_02893_),
    .B(_02938_),
    .C(_02942_),
    .Y(_02943_));
 sky130_fd_sc_hd__nand2_1 _08772_ (.A(_02893_),
    .B(_02942_),
    .Y(_02944_));
 sky130_fd_sc_hd__nand2_1 _08773_ (.A(_02944_),
    .B(_02937_),
    .Y(_02945_));
 sky130_fd_sc_hd__nand3_2 _08774_ (.A(_02834_),
    .B(_02943_),
    .C(_02945_),
    .Y(_02946_));
 sky130_fd_sc_hd__nand2_1 _08775_ (.A(_02945_),
    .B(_02943_),
    .Y(_02947_));
 sky130_fd_sc_hd__a21boi_1 _08776_ (.A1(_02617_),
    .A2(_02661_),
    .B1_N(_02618_),
    .Y(_02948_));
 sky130_fd_sc_hd__nand2_1 _08777_ (.A(_02947_),
    .B(_02948_),
    .Y(_02949_));
 sky130_fd_sc_hd__nand2_1 _08778_ (.A(_02946_),
    .B(_02949_),
    .Y(_02950_));
 sky130_fd_sc_hd__inv_2 _08779_ (.A(net3),
    .Y(_02952_));
 sky130_fd_sc_hd__nand2_1 _08780_ (.A(_04808_),
    .B(_02753_),
    .Y(_02953_));
 sky130_fd_sc_hd__or3_1 _08781_ (.A(_00263_),
    .B(_02952_),
    .C(_02953_),
    .X(_02954_));
 sky130_fd_sc_hd__o21ai_1 _08782_ (.A1(_00263_),
    .A2(_02952_),
    .B1(_02953_),
    .Y(_02955_));
 sky130_fd_sc_hd__nand2_1 _08783_ (.A(_02954_),
    .B(_02955_),
    .Y(_02956_));
 sky130_fd_sc_hd__nand2_1 _08784_ (.A(_04818_),
    .B(_03182_),
    .Y(_02957_));
 sky130_fd_sc_hd__nand2_1 _08785_ (.A(_02956_),
    .B(_02957_),
    .Y(_02958_));
 sky130_fd_sc_hd__nand3b_1 _08786_ (.A_N(_02957_),
    .B(_02954_),
    .C(_02955_),
    .Y(_02959_));
 sky130_fd_sc_hd__nand2_1 _08787_ (.A(_02958_),
    .B(_02959_),
    .Y(_02960_));
 sky130_fd_sc_hd__inv_2 _08788_ (.A(net5),
    .Y(_02961_));
 sky130_fd_sc_hd__o21ai_1 _08789_ (.A1(_01330_),
    .A2(_02961_),
    .B1(_02638_),
    .Y(_02963_));
 sky130_fd_sc_hd__nor3_1 _08790_ (.A(_01330_),
    .B(_02961_),
    .C(_02638_),
    .Y(_02964_));
 sky130_fd_sc_hd__a21oi_2 _08791_ (.A1(_02963_),
    .A2(_02637_),
    .B1(_02964_),
    .Y(_02965_));
 sky130_fd_sc_hd__inv_2 _08792_ (.A(_02965_),
    .Y(_02966_));
 sky130_fd_sc_hd__nand2_1 _08793_ (.A(_02960_),
    .B(_02966_),
    .Y(_02967_));
 sky130_fd_sc_hd__nand3_1 _08794_ (.A(_02958_),
    .B(_02959_),
    .C(_02965_),
    .Y(_02968_));
 sky130_fd_sc_hd__nand2_1 _08795_ (.A(_02967_),
    .B(_02968_),
    .Y(_02969_));
 sky130_fd_sc_hd__nand2_1 _08796_ (.A(_02679_),
    .B(_02673_),
    .Y(_02970_));
 sky130_fd_sc_hd__nand2_1 _08797_ (.A(_02969_),
    .B(_02970_),
    .Y(_02971_));
 sky130_fd_sc_hd__nand3b_1 _08798_ (.A_N(_02970_),
    .B(_02967_),
    .C(_02968_),
    .Y(_02972_));
 sky130_fd_sc_hd__nand2_1 _08799_ (.A(_02971_),
    .B(_02972_),
    .Y(_02974_));
 sky130_fd_sc_hd__nand2_1 _08800_ (.A(_02678_),
    .B(_02679_),
    .Y(_02975_));
 sky130_fd_sc_hd__nand2_1 _08801_ (.A(_02975_),
    .B(_02681_),
    .Y(_02976_));
 sky130_fd_sc_hd__nor2_1 _08802_ (.A(_02681_),
    .B(_02975_),
    .Y(_02977_));
 sky130_fd_sc_hd__a21oi_2 _08803_ (.A1(_02976_),
    .A2(_02685_),
    .B1(_02977_),
    .Y(_02978_));
 sky130_fd_sc_hd__inv_2 _08804_ (.A(_02978_),
    .Y(_02979_));
 sky130_fd_sc_hd__nand2_1 _08805_ (.A(_02974_),
    .B(_02979_),
    .Y(_02980_));
 sky130_fd_sc_hd__nand3_1 _08806_ (.A(_02971_),
    .B(_02972_),
    .C(_02978_),
    .Y(_02981_));
 sky130_fd_sc_hd__nand2_1 _08807_ (.A(_02980_),
    .B(_02981_),
    .Y(_02982_));
 sky130_fd_sc_hd__a21o_1 _08808_ (.A1(_02702_),
    .A2(_02706_),
    .B1(_02701_),
    .X(_02983_));
 sky130_fd_sc_hd__inv_2 _08809_ (.A(_02983_),
    .Y(_02985_));
 sky130_fd_sc_hd__nand2_1 _08810_ (.A(_04871_),
    .B(_03314_),
    .Y(_02986_));
 sky130_fd_sc_hd__or3_1 _08811_ (.A(_00110_),
    .B(_01596_),
    .C(_02986_),
    .X(_02987_));
 sky130_fd_sc_hd__o21ai_1 _08812_ (.A1(_00110_),
    .A2(_01596_),
    .B1(_02986_),
    .Y(_02988_));
 sky130_fd_sc_hd__nand2_1 _08813_ (.A(_02987_),
    .B(_02988_),
    .Y(_02989_));
 sky130_fd_sc_hd__nand2_1 _08814_ (.A(_04876_),
    .B(_03402_),
    .Y(_02990_));
 sky130_fd_sc_hd__nand2_1 _08815_ (.A(_02989_),
    .B(_02990_),
    .Y(_02991_));
 sky130_fd_sc_hd__nand3b_1 _08816_ (.A_N(_02990_),
    .B(_02987_),
    .C(_02988_),
    .Y(_02992_));
 sky130_fd_sc_hd__nand2_1 _08817_ (.A(_02991_),
    .B(_02992_),
    .Y(_02993_));
 sky130_fd_sc_hd__nor2_1 _08818_ (.A(_02985_),
    .B(_02993_),
    .Y(_02994_));
 sky130_fd_sc_hd__inv_2 _08819_ (.A(_02994_),
    .Y(_02996_));
 sky130_fd_sc_hd__nand2_1 _08820_ (.A(_02993_),
    .B(_02985_),
    .Y(_02997_));
 sky130_fd_sc_hd__nand2_1 _08821_ (.A(_02996_),
    .B(_02997_),
    .Y(_02998_));
 sky130_fd_sc_hd__nand2_1 _08822_ (.A(_00529_),
    .B(_04819_),
    .Y(_02999_));
 sky130_fd_sc_hd__inv_2 _08823_ (.A(_02999_),
    .Y(_03000_));
 sky130_fd_sc_hd__nand2_1 _08824_ (.A(_00124_),
    .B(_04809_),
    .Y(_03001_));
 sky130_fd_sc_hd__nand2_1 _08825_ (.A(net46),
    .B(_03820_),
    .Y(_03002_));
 sky130_fd_sc_hd__xor2_1 _08826_ (.A(_03001_),
    .B(_03002_),
    .X(_03003_));
 sky130_fd_sc_hd__or2_1 _08827_ (.A(_03000_),
    .B(_03003_),
    .X(_03004_));
 sky130_fd_sc_hd__nand2_1 _08828_ (.A(_03003_),
    .B(_03000_),
    .Y(_03005_));
 sky130_fd_sc_hd__nand2_1 _08829_ (.A(_03004_),
    .B(_03005_),
    .Y(_03007_));
 sky130_fd_sc_hd__nand2_1 _08830_ (.A(_02998_),
    .B(_03007_),
    .Y(_03008_));
 sky130_fd_sc_hd__inv_2 _08831_ (.A(_03007_),
    .Y(_03009_));
 sky130_fd_sc_hd__nand3_1 _08832_ (.A(_02996_),
    .B(_03009_),
    .C(_02997_),
    .Y(_03010_));
 sky130_fd_sc_hd__nand2_1 _08833_ (.A(_03008_),
    .B(_03010_),
    .Y(_03011_));
 sky130_fd_sc_hd__inv_2 _08834_ (.A(_03011_),
    .Y(_03012_));
 sky130_fd_sc_hd__nand2_1 _08835_ (.A(_02982_),
    .B(_03012_),
    .Y(_03013_));
 sky130_fd_sc_hd__nand3_1 _08836_ (.A(_02980_),
    .B(_03011_),
    .C(_02981_),
    .Y(_03014_));
 sky130_fd_sc_hd__nand2_1 _08837_ (.A(_03013_),
    .B(_03014_),
    .Y(_03015_));
 sky130_fd_sc_hd__nand2_1 _08838_ (.A(_02647_),
    .B(_02650_),
    .Y(_03016_));
 sky130_fd_sc_hd__nor2_1 _08839_ (.A(_02650_),
    .B(_02647_),
    .Y(_03018_));
 sky130_fd_sc_hd__a21oi_2 _08840_ (.A1(_03016_),
    .A2(_02657_),
    .B1(_03018_),
    .Y(_03019_));
 sky130_fd_sc_hd__inv_2 _08841_ (.A(_03019_),
    .Y(_03020_));
 sky130_fd_sc_hd__nand2_1 _08842_ (.A(_03015_),
    .B(_03020_),
    .Y(_03021_));
 sky130_fd_sc_hd__nand3_1 _08843_ (.A(_03019_),
    .B(_03013_),
    .C(_03014_),
    .Y(_03022_));
 sky130_fd_sc_hd__nand2_1 _08844_ (.A(_03021_),
    .B(_03022_),
    .Y(_03023_));
 sky130_fd_sc_hd__o21ai_1 _08845_ (.A1(_02693_),
    .A2(_02690_),
    .B1(_02730_),
    .Y(_03024_));
 sky130_fd_sc_hd__nand2_1 _08846_ (.A(_03023_),
    .B(_03024_),
    .Y(_03025_));
 sky130_fd_sc_hd__nand3b_1 _08847_ (.A_N(_03024_),
    .B(_03021_),
    .C(_03022_),
    .Y(_03026_));
 sky130_fd_sc_hd__nand2_1 _08848_ (.A(_03025_),
    .B(_03026_),
    .Y(_03027_));
 sky130_fd_sc_hd__nand2_1 _08849_ (.A(_02950_),
    .B(_03027_),
    .Y(_03029_));
 sky130_fd_sc_hd__inv_2 _08850_ (.A(_03027_),
    .Y(_03030_));
 sky130_fd_sc_hd__nand3_2 _08851_ (.A(_02946_),
    .B(_02949_),
    .C(_03030_),
    .Y(_03031_));
 sky130_fd_sc_hd__nand2_1 _08852_ (.A(_03029_),
    .B(_03031_),
    .Y(_03032_));
 sky130_fd_sc_hd__nand2_1 _08853_ (.A(_02667_),
    .B(_02554_),
    .Y(_03033_));
 sky130_fd_sc_hd__nor2_1 _08854_ (.A(_02554_),
    .B(_02667_),
    .Y(_03034_));
 sky130_fd_sc_hd__a21oi_4 _08855_ (.A1(_03033_),
    .A2(_02746_),
    .B1(_03034_),
    .Y(_03035_));
 sky130_fd_sc_hd__nand2_1 _08856_ (.A(_03032_),
    .B(_03035_),
    .Y(_03036_));
 sky130_fd_sc_hd__nand2_1 _08857_ (.A(_02733_),
    .B(_02736_),
    .Y(_03037_));
 sky130_fd_sc_hd__nor2_1 _08858_ (.A(_02736_),
    .B(_02733_),
    .Y(_03038_));
 sky130_fd_sc_hd__a21o_1 _08859_ (.A1(_03037_),
    .A2(_02741_),
    .B1(_03038_),
    .X(_03040_));
 sky130_fd_sc_hd__a21boi_1 _08860_ (.A1(_02726_),
    .A2(_02714_),
    .B1_N(_02713_),
    .Y(_03041_));
 sky130_fd_sc_hd__inv_2 _08861_ (.A(net49),
    .Y(_03042_));
 sky130_fd_sc_hd__nand2_1 _08862_ (.A(net50),
    .B(_04911_),
    .Y(_03043_));
 sky130_fd_sc_hd__or3_1 _08863_ (.A(_03042_),
    .B(_02085_),
    .C(_03043_),
    .X(_03044_));
 sky130_fd_sc_hd__o21ai_1 _08864_ (.A1(_03042_),
    .A2(_02085_),
    .B1(_03043_),
    .Y(_03045_));
 sky130_fd_sc_hd__nand2_1 _08865_ (.A(_03044_),
    .B(_03045_),
    .Y(_03046_));
 sky130_fd_sc_hd__nand2_1 _08866_ (.A(net51),
    .B(_04895_),
    .Y(_03047_));
 sky130_fd_sc_hd__nand2_1 _08867_ (.A(_03046_),
    .B(_03047_),
    .Y(_03048_));
 sky130_fd_sc_hd__nand3b_1 _08868_ (.A_N(_03047_),
    .B(_03044_),
    .C(_03045_),
    .Y(_03049_));
 sky130_fd_sc_hd__nand2_1 _08869_ (.A(_03048_),
    .B(_03049_),
    .Y(_03051_));
 sky130_fd_sc_hd__inv_2 _08870_ (.A(_02716_),
    .Y(_03052_));
 sky130_fd_sc_hd__a21oi_1 _08871_ (.A1(_02719_),
    .A2(_03052_),
    .B1(_02718_),
    .Y(_03053_));
 sky130_fd_sc_hd__nand2_1 _08872_ (.A(_03051_),
    .B(_03053_),
    .Y(_03054_));
 sky130_fd_sc_hd__nand3b_1 _08873_ (.A_N(_03053_),
    .B(_03048_),
    .C(_03049_),
    .Y(_03055_));
 sky130_fd_sc_hd__nand2_1 _08874_ (.A(_03054_),
    .B(_03055_),
    .Y(_03056_));
 sky130_fd_sc_hd__nand2_1 _08875_ (.A(_03056_),
    .B(_02763_),
    .Y(_03057_));
 sky130_fd_sc_hd__nand3_1 _08876_ (.A(_03054_),
    .B(_03055_),
    .C(_02762_),
    .Y(_03058_));
 sky130_fd_sc_hd__nand2_1 _08877_ (.A(_03057_),
    .B(_03058_),
    .Y(_03059_));
 sky130_fd_sc_hd__nor2_1 _08878_ (.A(_03041_),
    .B(_03059_),
    .Y(_03060_));
 sky130_fd_sc_hd__nand2_1 _08879_ (.A(_03059_),
    .B(_03041_),
    .Y(_03062_));
 sky130_fd_sc_hd__nand2b_1 _08880_ (.A_N(_03060_),
    .B(_03062_),
    .Y(_03063_));
 sky130_fd_sc_hd__nand2_1 _08881_ (.A(_03063_),
    .B(_02769_),
    .Y(_03064_));
 sky130_fd_sc_hd__nand3b_1 _08882_ (.A_N(_03060_),
    .B(_02768_),
    .C(_03062_),
    .Y(_03065_));
 sky130_fd_sc_hd__nand2_1 _08883_ (.A(_02778_),
    .B(_02773_),
    .Y(_03066_));
 sky130_fd_sc_hd__nand3_2 _08884_ (.A(_03064_),
    .B(_03065_),
    .C(_03066_),
    .Y(_03067_));
 sky130_fd_sc_hd__nand2_1 _08885_ (.A(_03064_),
    .B(_03065_),
    .Y(_03068_));
 sky130_fd_sc_hd__nand3_1 _08886_ (.A(_03068_),
    .B(_02773_),
    .C(_02778_),
    .Y(_03069_));
 sky130_fd_sc_hd__nand3_1 _08887_ (.A(_03040_),
    .B(_03067_),
    .C(_03069_),
    .Y(_03070_));
 sky130_fd_sc_hd__nand2_1 _08888_ (.A(_03069_),
    .B(_03067_),
    .Y(_03071_));
 sky130_fd_sc_hd__a21oi_1 _08889_ (.A1(_03037_),
    .A2(_02741_),
    .B1(_03038_),
    .Y(_03073_));
 sky130_fd_sc_hd__nand2_1 _08890_ (.A(_03071_),
    .B(_03073_),
    .Y(_03074_));
 sky130_fd_sc_hd__nand2_1 _08891_ (.A(_03070_),
    .B(_03074_),
    .Y(_03075_));
 sky130_fd_sc_hd__nand2_1 _08892_ (.A(_03075_),
    .B(_02781_),
    .Y(_03076_));
 sky130_fd_sc_hd__inv_2 _08893_ (.A(_02781_),
    .Y(_03077_));
 sky130_fd_sc_hd__nand3_1 _08894_ (.A(_03070_),
    .B(_03074_),
    .C(_03077_),
    .Y(_03078_));
 sky130_fd_sc_hd__nand2_1 _08895_ (.A(_03076_),
    .B(_03078_),
    .Y(_03079_));
 sky130_fd_sc_hd__inv_2 _08896_ (.A(_03079_),
    .Y(_03080_));
 sky130_fd_sc_hd__nor2_1 _08897_ (.A(_03035_),
    .B(_03032_),
    .Y(_03081_));
 sky130_fd_sc_hd__a21o_1 _08898_ (.A1(_03036_),
    .A2(_03080_),
    .B1(_03081_),
    .X(_03082_));
 sky130_fd_sc_hd__nand2_1 _08899_ (.A(_03031_),
    .B(_02946_),
    .Y(_03084_));
 sky130_fd_sc_hd__nand2_1 _08900_ (.A(_02943_),
    .B(_02893_),
    .Y(_03085_));
 sky130_fd_sc_hd__nand2_1 _08901_ (.A(_02892_),
    .B(_02868_),
    .Y(_03086_));
 sky130_fd_sc_hd__inv_2 _08902_ (.A(net20),
    .Y(_03087_));
 sky130_fd_sc_hd__nand2_1 _08903_ (.A(_02357_),
    .B(net19),
    .Y(_03088_));
 sky130_fd_sc_hd__nor3_1 _08904_ (.A(_01597_),
    .B(_03087_),
    .C(_03088_),
    .Y(_03089_));
 sky130_fd_sc_hd__inv_2 _08905_ (.A(_03089_),
    .Y(_03090_));
 sky130_fd_sc_hd__o21ai_1 _08906_ (.A1(_01597_),
    .A2(_03087_),
    .B1(_03088_),
    .Y(_03091_));
 sky130_fd_sc_hd__nand2_1 _08907_ (.A(_01535_),
    .B(net18),
    .Y(_03092_));
 sky130_fd_sc_hd__a21bo_1 _08908_ (.A1(_03090_),
    .A2(_03091_),
    .B1_N(_03092_),
    .X(_03093_));
 sky130_fd_sc_hd__nand3b_1 _08909_ (.A_N(_03092_),
    .B(_03090_),
    .C(_03091_),
    .Y(_03095_));
 sky130_fd_sc_hd__nand2_1 _08910_ (.A(_03093_),
    .B(_03095_),
    .Y(_03096_));
 sky130_fd_sc_hd__nand2_1 _08911_ (.A(_02845_),
    .B(_02839_),
    .Y(_03097_));
 sky130_fd_sc_hd__inv_2 _08912_ (.A(_03097_),
    .Y(_03098_));
 sky130_fd_sc_hd__nand2_1 _08913_ (.A(_03096_),
    .B(_03098_),
    .Y(_03099_));
 sky130_fd_sc_hd__nand3_1 _08914_ (.A(_03093_),
    .B(_03097_),
    .C(_03095_),
    .Y(_03100_));
 sky130_fd_sc_hd__nand2_1 _08915_ (.A(_03099_),
    .B(_03100_),
    .Y(_03101_));
 sky130_fd_sc_hd__nand2_1 _08916_ (.A(_01565_),
    .B(_05160_),
    .Y(_03102_));
 sky130_fd_sc_hd__inv_2 _08917_ (.A(_03102_),
    .Y(_03103_));
 sky130_fd_sc_hd__nand2_1 _08918_ (.A(_04260_),
    .B(_00393_),
    .Y(_03104_));
 sky130_fd_sc_hd__nand2_1 _08919_ (.A(_04293_),
    .B(net17),
    .Y(_03106_));
 sky130_fd_sc_hd__xor2_1 _08920_ (.A(_03104_),
    .B(_03106_),
    .X(_03107_));
 sky130_fd_sc_hd__or2_1 _08921_ (.A(_03103_),
    .B(_03107_),
    .X(_03108_));
 sky130_fd_sc_hd__nand2_1 _08922_ (.A(_03107_),
    .B(_03103_),
    .Y(_03109_));
 sky130_fd_sc_hd__nand2_1 _08923_ (.A(_03108_),
    .B(_03109_),
    .Y(_03110_));
 sky130_fd_sc_hd__nand2_1 _08924_ (.A(_03101_),
    .B(_03110_),
    .Y(_03111_));
 sky130_fd_sc_hd__nand3b_1 _08925_ (.A_N(_03110_),
    .B(_03099_),
    .C(_03100_),
    .Y(_03112_));
 sky130_fd_sc_hd__nand2_1 _08926_ (.A(_03111_),
    .B(_03112_),
    .Y(_03113_));
 sky130_fd_sc_hd__nand2_1 _08927_ (.A(_02862_),
    .B(_02846_),
    .Y(_03114_));
 sky130_fd_sc_hd__inv_2 _08928_ (.A(_03114_),
    .Y(_03115_));
 sky130_fd_sc_hd__nand2_1 _08929_ (.A(_03113_),
    .B(_03115_),
    .Y(_03117_));
 sky130_fd_sc_hd__nand3_1 _08930_ (.A(_03114_),
    .B(_03111_),
    .C(_03112_),
    .Y(_03118_));
 sky130_fd_sc_hd__nand2_1 _08931_ (.A(_03117_),
    .B(_03118_),
    .Y(_03119_));
 sky130_fd_sc_hd__and2_1 _08932_ (.A(_02878_),
    .B(_02872_),
    .X(_03120_));
 sky130_fd_sc_hd__nand2_2 _08933_ (.A(_02859_),
    .B(_02854_),
    .Y(_03121_));
 sky130_fd_sc_hd__inv_2 _08934_ (.A(_03121_),
    .Y(_03122_));
 sky130_fd_sc_hd__nand2_1 _08935_ (.A(_00784_),
    .B(_00003_),
    .Y(_03123_));
 sky130_fd_sc_hd__inv_2 _08936_ (.A(_03123_),
    .Y(_03124_));
 sky130_fd_sc_hd__nand2_1 _08937_ (.A(_01323_),
    .B(_00412_),
    .Y(_03125_));
 sky130_fd_sc_hd__nand2_1 _08938_ (.A(_00204_),
    .B(_04084_),
    .Y(_03126_));
 sky130_fd_sc_hd__xor2_1 _08939_ (.A(_03125_),
    .B(_03126_),
    .X(_03128_));
 sky130_fd_sc_hd__or2_1 _08940_ (.A(_03124_),
    .B(_03128_),
    .X(_03129_));
 sky130_fd_sc_hd__nand2_1 _08941_ (.A(_03128_),
    .B(_03124_),
    .Y(_03130_));
 sky130_fd_sc_hd__nand2_1 _08942_ (.A(_03129_),
    .B(_03130_),
    .Y(_03131_));
 sky130_fd_sc_hd__or2_1 _08943_ (.A(_03122_),
    .B(_03131_),
    .X(_03132_));
 sky130_fd_sc_hd__nand2_1 _08944_ (.A(_03131_),
    .B(_03122_),
    .Y(_03133_));
 sky130_fd_sc_hd__nand3b_1 _08945_ (.A_N(_03120_),
    .B(_03132_),
    .C(_03133_),
    .Y(_03134_));
 sky130_fd_sc_hd__nor2_1 _08946_ (.A(_03121_),
    .B(_03131_),
    .Y(_03135_));
 sky130_fd_sc_hd__nand2_1 _08947_ (.A(_03131_),
    .B(_03121_),
    .Y(_03136_));
 sky130_fd_sc_hd__nand3b_1 _08948_ (.A_N(_03135_),
    .B(_03120_),
    .C(_03136_),
    .Y(_03137_));
 sky130_fd_sc_hd__nand2_1 _08949_ (.A(_03134_),
    .B(_03137_),
    .Y(_03139_));
 sky130_fd_sc_hd__nand2_1 _08950_ (.A(_03119_),
    .B(_03139_),
    .Y(_03140_));
 sky130_fd_sc_hd__inv_2 _08951_ (.A(_03139_),
    .Y(_03141_));
 sky130_fd_sc_hd__nand3_1 _08952_ (.A(_03141_),
    .B(_03117_),
    .C(_03118_),
    .Y(_03142_));
 sky130_fd_sc_hd__nand3_2 _08953_ (.A(_03086_),
    .B(_03140_),
    .C(_03142_),
    .Y(_03143_));
 sky130_fd_sc_hd__inv_2 _08954_ (.A(_03086_),
    .Y(_03144_));
 sky130_fd_sc_hd__nand2_1 _08955_ (.A(_03140_),
    .B(_03142_),
    .Y(_03145_));
 sky130_fd_sc_hd__nand2_1 _08956_ (.A(_03144_),
    .B(_03145_),
    .Y(_03146_));
 sky130_fd_sc_hd__nand2_1 _08957_ (.A(_03143_),
    .B(_03146_),
    .Y(_03147_));
 sky130_fd_sc_hd__nand2_1 _08958_ (.A(_02879_),
    .B(_02882_),
    .Y(_03148_));
 sky130_fd_sc_hd__nor2_1 _08959_ (.A(_02882_),
    .B(_02879_),
    .Y(_03150_));
 sky130_fd_sc_hd__a21oi_1 _08960_ (.A1(_03148_),
    .A2(_02886_),
    .B1(_03150_),
    .Y(_03151_));
 sky130_fd_sc_hd__nand2_1 _08961_ (.A(_03809_),
    .B(_02544_),
    .Y(_03152_));
 sky130_fd_sc_hd__inv_2 _08962_ (.A(_03152_),
    .Y(_03153_));
 sky130_fd_sc_hd__nand2_1 _08963_ (.A(_04962_),
    .B(_01147_),
    .Y(_03154_));
 sky130_fd_sc_hd__nand2_1 _08964_ (.A(_04964_),
    .B(_01037_),
    .Y(_03155_));
 sky130_fd_sc_hd__xor2_1 _08965_ (.A(_03154_),
    .B(_03155_),
    .X(_03156_));
 sky130_fd_sc_hd__or2_1 _08966_ (.A(_03153_),
    .B(_03156_),
    .X(_03157_));
 sky130_fd_sc_hd__nand2_1 _08967_ (.A(_03156_),
    .B(_03153_),
    .Y(_03158_));
 sky130_fd_sc_hd__nand2_1 _08968_ (.A(_03157_),
    .B(_03158_),
    .Y(_03159_));
 sky130_fd_sc_hd__nand2_1 _08969_ (.A(_03215_),
    .B(_01081_),
    .Y(_03161_));
 sky130_fd_sc_hd__inv_2 _08970_ (.A(_03161_),
    .Y(_03162_));
 sky130_fd_sc_hd__nand2_1 _08971_ (.A(_00850_),
    .B(_05029_),
    .Y(_03163_));
 sky130_fd_sc_hd__nand2_1 _08972_ (.A(_00740_),
    .B(_05032_),
    .Y(_03164_));
 sky130_fd_sc_hd__xor2_1 _08973_ (.A(_03163_),
    .B(_03164_),
    .X(_03165_));
 sky130_fd_sc_hd__or2_1 _08974_ (.A(_03162_),
    .B(_03165_),
    .X(_03166_));
 sky130_fd_sc_hd__nand2_1 _08975_ (.A(_03165_),
    .B(_03162_),
    .Y(_03167_));
 sky130_fd_sc_hd__nand2_1 _08976_ (.A(_03166_),
    .B(_03167_),
    .Y(_03168_));
 sky130_fd_sc_hd__a21oi_1 _08977_ (.A1(_02899_),
    .A2(_02901_),
    .B1(_02897_),
    .Y(_03169_));
 sky130_fd_sc_hd__nand2_1 _08978_ (.A(_03168_),
    .B(_03169_),
    .Y(_03170_));
 sky130_fd_sc_hd__nand3b_1 _08979_ (.A_N(_03169_),
    .B(_03166_),
    .C(_03167_),
    .Y(_03172_));
 sky130_fd_sc_hd__nand3b_1 _08980_ (.A_N(_03159_),
    .B(_03170_),
    .C(_03172_),
    .Y(_03173_));
 sky130_fd_sc_hd__nand2_1 _08981_ (.A(_03170_),
    .B(_03172_),
    .Y(_03174_));
 sky130_fd_sc_hd__nand2_1 _08982_ (.A(_03174_),
    .B(_03159_),
    .Y(_03175_));
 sky130_fd_sc_hd__nand3_1 _08983_ (.A(_03151_),
    .B(_03173_),
    .C(_03175_),
    .Y(_03176_));
 sky130_fd_sc_hd__a21o_1 _08984_ (.A1(_03148_),
    .A2(_02886_),
    .B1(_03150_),
    .X(_03177_));
 sky130_fd_sc_hd__nand2_1 _08985_ (.A(_03175_),
    .B(_03173_),
    .Y(_03178_));
 sky130_fd_sc_hd__nand2_1 _08986_ (.A(_03177_),
    .B(_03178_),
    .Y(_03179_));
 sky130_fd_sc_hd__nand2_1 _08987_ (.A(_03176_),
    .B(_03179_),
    .Y(_03180_));
 sky130_fd_sc_hd__o21ai_1 _08988_ (.A1(_02908_),
    .A2(_02904_),
    .B1(_02923_),
    .Y(_03181_));
 sky130_fd_sc_hd__nand2_1 _08989_ (.A(_03180_),
    .B(_03181_),
    .Y(_03183_));
 sky130_fd_sc_hd__nand3b_1 _08990_ (.A_N(_03181_),
    .B(_03176_),
    .C(_03179_),
    .Y(_03184_));
 sky130_fd_sc_hd__nand2_1 _08991_ (.A(_03183_),
    .B(_03184_),
    .Y(_03185_));
 sky130_fd_sc_hd__nand2_1 _08992_ (.A(_03147_),
    .B(_03185_),
    .Y(_03186_));
 sky130_fd_sc_hd__nand3b_2 _08993_ (.A_N(_03185_),
    .B(_03143_),
    .C(_03146_),
    .Y(_03187_));
 sky130_fd_sc_hd__nand3_2 _08994_ (.A(_03085_),
    .B(_03186_),
    .C(_03187_),
    .Y(_03188_));
 sky130_fd_sc_hd__and2_1 _08995_ (.A(_02959_),
    .B(_02954_),
    .X(_03189_));
 sky130_fd_sc_hd__nand2_1 _08996_ (.A(_04818_),
    .B(_03160_),
    .Y(_03190_));
 sky130_fd_sc_hd__inv_2 _08997_ (.A(_03190_),
    .Y(_03191_));
 sky130_fd_sc_hd__nand2_1 _08998_ (.A(_04808_),
    .B(_02049_),
    .Y(_03192_));
 sky130_fd_sc_hd__nor3_1 _08999_ (.A(_00263_),
    .B(_02410_),
    .C(_03192_),
    .Y(_03194_));
 sky130_fd_sc_hd__o21ai_1 _09000_ (.A1(_00263_),
    .A2(_02410_),
    .B1(_03192_),
    .Y(_03195_));
 sky130_fd_sc_hd__nor2b_1 _09001_ (.A(_03194_),
    .B_N(_03195_),
    .Y(_03196_));
 sky130_fd_sc_hd__or2_1 _09002_ (.A(_03191_),
    .B(_03196_),
    .X(_03197_));
 sky130_fd_sc_hd__nand2_1 _09003_ (.A(_03196_),
    .B(_03191_),
    .Y(_03198_));
 sky130_fd_sc_hd__nand2_1 _09004_ (.A(_03197_),
    .B(_03198_),
    .Y(_03199_));
 sky130_fd_sc_hd__a21oi_1 _09005_ (.A1(_02916_),
    .A2(_02912_),
    .B1(_02915_),
    .Y(_03200_));
 sky130_fd_sc_hd__nand2_1 _09006_ (.A(_03199_),
    .B(_03200_),
    .Y(_03201_));
 sky130_fd_sc_hd__inv_2 _09007_ (.A(_03200_),
    .Y(_03202_));
 sky130_fd_sc_hd__nand3_1 _09008_ (.A(_03197_),
    .B(_03198_),
    .C(_03202_),
    .Y(_03203_));
 sky130_fd_sc_hd__nand3b_1 _09009_ (.A_N(_03189_),
    .B(_03201_),
    .C(_03203_),
    .Y(_03205_));
 sky130_fd_sc_hd__nand2_1 _09010_ (.A(_03201_),
    .B(_03203_),
    .Y(_03206_));
 sky130_fd_sc_hd__nand2_1 _09011_ (.A(_03206_),
    .B(_03189_),
    .Y(_03207_));
 sky130_fd_sc_hd__nand2_1 _09012_ (.A(_03205_),
    .B(_03207_),
    .Y(_03208_));
 sky130_fd_sc_hd__nand2_1 _09013_ (.A(_02960_),
    .B(_02965_),
    .Y(_03209_));
 sky130_fd_sc_hd__nor2_1 _09014_ (.A(_02965_),
    .B(_02960_),
    .Y(_03210_));
 sky130_fd_sc_hd__a21oi_2 _09015_ (.A1(_03209_),
    .A2(_02970_),
    .B1(_03210_),
    .Y(_03211_));
 sky130_fd_sc_hd__inv_2 _09016_ (.A(_03211_),
    .Y(_03212_));
 sky130_fd_sc_hd__nand2_1 _09017_ (.A(_03208_),
    .B(_03212_),
    .Y(_03213_));
 sky130_fd_sc_hd__nand3_1 _09018_ (.A(_03211_),
    .B(_03205_),
    .C(_03207_),
    .Y(_03214_));
 sky130_fd_sc_hd__nand2_1 _09019_ (.A(_03213_),
    .B(_03214_),
    .Y(_03216_));
 sky130_fd_sc_hd__nand2_1 _09020_ (.A(_04876_),
    .B(_05028_),
    .Y(_03217_));
 sky130_fd_sc_hd__inv_2 _09021_ (.A(_03217_),
    .Y(_03218_));
 sky130_fd_sc_hd__and4_1 _09022_ (.A(_04873_),
    .B(_04871_),
    .C(_03094_),
    .D(_03226_),
    .X(_03219_));
 sky130_fd_sc_hd__a22o_1 _09023_ (.A1(_04873_),
    .A2(_03182_),
    .B1(_04871_),
    .B2(_05031_),
    .X(_03220_));
 sky130_fd_sc_hd__nor2b_1 _09024_ (.A(_03219_),
    .B_N(_03220_),
    .Y(_03221_));
 sky130_fd_sc_hd__or2_1 _09025_ (.A(_03218_),
    .B(_03221_),
    .X(_03222_));
 sky130_fd_sc_hd__nand2_1 _09026_ (.A(_03221_),
    .B(_03218_),
    .Y(_03223_));
 sky130_fd_sc_hd__nand2_1 _09027_ (.A(_03222_),
    .B(_03223_),
    .Y(_03224_));
 sky130_fd_sc_hd__nand2_1 _09028_ (.A(_02992_),
    .B(_02987_),
    .Y(_03225_));
 sky130_fd_sc_hd__nand2_1 _09029_ (.A(_03224_),
    .B(_03225_),
    .Y(_03227_));
 sky130_fd_sc_hd__inv_2 _09030_ (.A(_03225_),
    .Y(_03228_));
 sky130_fd_sc_hd__nand3_1 _09031_ (.A(_03222_),
    .B(_03228_),
    .C(_03223_),
    .Y(_03229_));
 sky130_fd_sc_hd__nand2_1 _09032_ (.A(_03227_),
    .B(_03229_),
    .Y(_03230_));
 sky130_fd_sc_hd__nand2_1 _09033_ (.A(_00529_),
    .B(_00254_),
    .Y(_03231_));
 sky130_fd_sc_hd__nand2_1 _09034_ (.A(_00124_),
    .B(_00656_),
    .Y(_03232_));
 sky130_fd_sc_hd__nor3_1 _09035_ (.A(_02463_),
    .B(_02451_),
    .C(_03232_),
    .Y(_03233_));
 sky130_fd_sc_hd__o21ai_1 _09036_ (.A1(_02463_),
    .A2(_02451_),
    .B1(_03232_),
    .Y(_03234_));
 sky130_fd_sc_hd__inv_2 _09037_ (.A(_03234_),
    .Y(_03235_));
 sky130_fd_sc_hd__nor2_1 _09038_ (.A(_03233_),
    .B(_03235_),
    .Y(_03236_));
 sky130_fd_sc_hd__xor2_1 _09039_ (.A(_03231_),
    .B(_03236_),
    .X(_03238_));
 sky130_fd_sc_hd__inv_2 _09040_ (.A(_03238_),
    .Y(_03239_));
 sky130_fd_sc_hd__nand2_1 _09041_ (.A(_03230_),
    .B(_03239_),
    .Y(_03240_));
 sky130_fd_sc_hd__nand3_1 _09042_ (.A(_03227_),
    .B(_03229_),
    .C(_03238_),
    .Y(_03241_));
 sky130_fd_sc_hd__nand2_1 _09043_ (.A(_03240_),
    .B(_03241_),
    .Y(_03242_));
 sky130_fd_sc_hd__inv_2 _09044_ (.A(_03242_),
    .Y(_03243_));
 sky130_fd_sc_hd__nand2_1 _09045_ (.A(_03216_),
    .B(_03243_),
    .Y(_03244_));
 sky130_fd_sc_hd__nand3_1 _09046_ (.A(_03242_),
    .B(_03213_),
    .C(_03214_),
    .Y(_03245_));
 sky130_fd_sc_hd__nand2_1 _09047_ (.A(_03244_),
    .B(_03245_),
    .Y(_03246_));
 sky130_fd_sc_hd__nand2_1 _09048_ (.A(_02925_),
    .B(_02928_),
    .Y(_03247_));
 sky130_fd_sc_hd__nor2_1 _09049_ (.A(_02928_),
    .B(_02925_),
    .Y(_03249_));
 sky130_fd_sc_hd__a21oi_2 _09050_ (.A1(_03247_),
    .A2(_02934_),
    .B1(_03249_),
    .Y(_03250_));
 sky130_fd_sc_hd__inv_2 _09051_ (.A(_03250_),
    .Y(_03251_));
 sky130_fd_sc_hd__nand2_1 _09052_ (.A(_03246_),
    .B(_03251_),
    .Y(_03252_));
 sky130_fd_sc_hd__nand3_1 _09053_ (.A(_03244_),
    .B(_03245_),
    .C(_03250_),
    .Y(_03253_));
 sky130_fd_sc_hd__nand2_1 _09054_ (.A(_03252_),
    .B(_03253_),
    .Y(_03254_));
 sky130_fd_sc_hd__nor2_1 _09055_ (.A(_02978_),
    .B(_02974_),
    .Y(_03255_));
 sky130_fd_sc_hd__inv_2 _09056_ (.A(_03013_),
    .Y(_03256_));
 sky130_fd_sc_hd__nor2_1 _09057_ (.A(_03255_),
    .B(_03256_),
    .Y(_03257_));
 sky130_fd_sc_hd__inv_2 _09058_ (.A(_03257_),
    .Y(_03258_));
 sky130_fd_sc_hd__nand2_1 _09059_ (.A(_03254_),
    .B(_03258_),
    .Y(_03260_));
 sky130_fd_sc_hd__nand3_1 _09060_ (.A(_03252_),
    .B(_03253_),
    .C(_03257_),
    .Y(_03261_));
 sky130_fd_sc_hd__nand2_1 _09061_ (.A(_03260_),
    .B(_03261_),
    .Y(_03262_));
 sky130_fd_sc_hd__inv_2 _09062_ (.A(_03262_),
    .Y(_03263_));
 sky130_fd_sc_hd__nand2_1 _09063_ (.A(_03186_),
    .B(_03187_),
    .Y(_03264_));
 sky130_fd_sc_hd__a21boi_1 _09064_ (.A1(_02938_),
    .A2(_02942_),
    .B1_N(_02893_),
    .Y(_03265_));
 sky130_fd_sc_hd__nand2_1 _09065_ (.A(_03264_),
    .B(_03265_),
    .Y(_03266_));
 sky130_fd_sc_hd__nand3_2 _09066_ (.A(_03188_),
    .B(_03263_),
    .C(_03266_),
    .Y(_03267_));
 sky130_fd_sc_hd__nand2_1 _09067_ (.A(_03188_),
    .B(_03266_),
    .Y(_03268_));
 sky130_fd_sc_hd__nand2_1 _09068_ (.A(_03268_),
    .B(_03262_),
    .Y(_03269_));
 sky130_fd_sc_hd__nand3_2 _09069_ (.A(_03084_),
    .B(_03267_),
    .C(_03269_),
    .Y(_03271_));
 sky130_fd_sc_hd__a21o_1 _09070_ (.A1(_02997_),
    .A2(_03009_),
    .B1(_02994_),
    .X(_03272_));
 sky130_fd_sc_hd__and2_1 _09071_ (.A(_03049_),
    .B(_03044_),
    .X(_03273_));
 sky130_fd_sc_hd__nand2_1 _09072_ (.A(net51),
    .B(_04991_),
    .Y(_03274_));
 sky130_fd_sc_hd__inv_2 _09073_ (.A(_03274_),
    .Y(_03275_));
 sky130_fd_sc_hd__nand2_1 _09074_ (.A(net50),
    .B(_04828_),
    .Y(_03276_));
 sky130_fd_sc_hd__nor3_1 _09075_ (.A(_03042_),
    .B(_02464_),
    .C(_03276_),
    .Y(_03277_));
 sky130_fd_sc_hd__o21ai_1 _09076_ (.A1(_03042_),
    .A2(_02464_),
    .B1(_03276_),
    .Y(_03278_));
 sky130_fd_sc_hd__nor2b_1 _09077_ (.A(_03277_),
    .B_N(_03278_),
    .Y(_03279_));
 sky130_fd_sc_hd__or2_1 _09078_ (.A(_03275_),
    .B(_03279_),
    .X(_03280_));
 sky130_fd_sc_hd__nand2_1 _09079_ (.A(_03279_),
    .B(_03275_),
    .Y(_03282_));
 sky130_fd_sc_hd__nand2_1 _09080_ (.A(_03280_),
    .B(_03282_),
    .Y(_03283_));
 sky130_fd_sc_hd__inv_2 _09081_ (.A(_00656_),
    .Y(_03284_));
 sky130_fd_sc_hd__o21ai_1 _09082_ (.A1(_02463_),
    .A2(_03284_),
    .B1(_03001_),
    .Y(_03285_));
 sky130_fd_sc_hd__nor3_1 _09083_ (.A(_02463_),
    .B(_03284_),
    .C(_03001_),
    .Y(_03286_));
 sky130_fd_sc_hd__a21oi_1 _09084_ (.A1(_03285_),
    .A2(_03000_),
    .B1(_03286_),
    .Y(_03287_));
 sky130_fd_sc_hd__nand2_1 _09085_ (.A(_03283_),
    .B(_03287_),
    .Y(_03288_));
 sky130_fd_sc_hd__inv_2 _09086_ (.A(_03287_),
    .Y(_03289_));
 sky130_fd_sc_hd__nand3_1 _09087_ (.A(_03280_),
    .B(_03282_),
    .C(_03289_),
    .Y(_03290_));
 sky130_fd_sc_hd__nand3b_1 _09088_ (.A_N(_03273_),
    .B(_03288_),
    .C(_03290_),
    .Y(_03291_));
 sky130_fd_sc_hd__nand2_1 _09089_ (.A(_03288_),
    .B(_03290_),
    .Y(_03293_));
 sky130_fd_sc_hd__nand2_1 _09090_ (.A(_03293_),
    .B(_03273_),
    .Y(_03294_));
 sky130_fd_sc_hd__nand3_1 _09091_ (.A(_03272_),
    .B(_03291_),
    .C(_03294_),
    .Y(_03295_));
 sky130_fd_sc_hd__nand2_1 _09092_ (.A(_03291_),
    .B(_03294_),
    .Y(_03296_));
 sky130_fd_sc_hd__a21oi_1 _09093_ (.A1(_02997_),
    .A2(_03009_),
    .B1(_02994_),
    .Y(_03297_));
 sky130_fd_sc_hd__nand2_1 _09094_ (.A(_03296_),
    .B(_03297_),
    .Y(_03298_));
 sky130_fd_sc_hd__nand2_1 _09095_ (.A(_03295_),
    .B(_03298_),
    .Y(_03299_));
 sky130_fd_sc_hd__nand2_1 _09096_ (.A(_03058_),
    .B(_03055_),
    .Y(_03300_));
 sky130_fd_sc_hd__inv_2 _09097_ (.A(_03300_),
    .Y(_03301_));
 sky130_fd_sc_hd__nand2_1 _09098_ (.A(_03299_),
    .B(_03301_),
    .Y(_03302_));
 sky130_fd_sc_hd__nand3_1 _09099_ (.A(_03295_),
    .B(_03298_),
    .C(_03300_),
    .Y(_03304_));
 sky130_fd_sc_hd__nand2_1 _09100_ (.A(_03302_),
    .B(_03304_),
    .Y(_03305_));
 sky130_fd_sc_hd__a21oi_1 _09101_ (.A1(_03062_),
    .A2(_02768_),
    .B1(_03060_),
    .Y(_03306_));
 sky130_fd_sc_hd__nand2_1 _09102_ (.A(_03305_),
    .B(_03306_),
    .Y(_03307_));
 sky130_fd_sc_hd__a21o_1 _09103_ (.A1(_03062_),
    .A2(_02768_),
    .B1(_03060_),
    .X(_03308_));
 sky130_fd_sc_hd__nand3_1 _09104_ (.A(_03308_),
    .B(_03302_),
    .C(_03304_),
    .Y(_03309_));
 sky130_fd_sc_hd__nand2_1 _09105_ (.A(_03307_),
    .B(_03309_),
    .Y(_03310_));
 sky130_fd_sc_hd__nand2_1 _09106_ (.A(net52),
    .B(_04992_),
    .Y(_03311_));
 sky130_fd_sc_hd__nand2_1 _09107_ (.A(_03310_),
    .B(_03311_),
    .Y(_03312_));
 sky130_fd_sc_hd__nand3b_1 _09108_ (.A_N(_03311_),
    .B(_03307_),
    .C(_03309_),
    .Y(_03313_));
 sky130_fd_sc_hd__nand2_1 _09109_ (.A(_03312_),
    .B(_03313_),
    .Y(_03315_));
 sky130_fd_sc_hd__nand2_1 _09110_ (.A(_03015_),
    .B(_03019_),
    .Y(_03316_));
 sky130_fd_sc_hd__nor2_1 _09111_ (.A(_03019_),
    .B(_03015_),
    .Y(_03317_));
 sky130_fd_sc_hd__a21o_1 _09112_ (.A1(_03316_),
    .A2(_03024_),
    .B1(_03317_),
    .X(_03318_));
 sky130_fd_sc_hd__inv_2 _09113_ (.A(_03318_),
    .Y(_03319_));
 sky130_fd_sc_hd__nand2_1 _09114_ (.A(_03315_),
    .B(_03319_),
    .Y(_03320_));
 sky130_fd_sc_hd__nand3_1 _09115_ (.A(_03318_),
    .B(_03312_),
    .C(_03313_),
    .Y(_03321_));
 sky130_fd_sc_hd__nand2_1 _09116_ (.A(_03320_),
    .B(_03321_),
    .Y(_03322_));
 sky130_fd_sc_hd__nand2_1 _09117_ (.A(_03322_),
    .B(_03067_),
    .Y(_03323_));
 sky130_fd_sc_hd__inv_2 _09118_ (.A(_03067_),
    .Y(_03324_));
 sky130_fd_sc_hd__nand3_1 _09119_ (.A(_03320_),
    .B(_03321_),
    .C(_03324_),
    .Y(_03326_));
 sky130_fd_sc_hd__nand2_1 _09120_ (.A(_03323_),
    .B(_03326_),
    .Y(_03327_));
 sky130_fd_sc_hd__inv_2 _09121_ (.A(_03327_),
    .Y(_03328_));
 sky130_fd_sc_hd__nand2_1 _09122_ (.A(_03269_),
    .B(_03267_),
    .Y(_03329_));
 sky130_fd_sc_hd__a21boi_1 _09123_ (.A1(_03030_),
    .A2(_02949_),
    .B1_N(_02946_),
    .Y(_03330_));
 sky130_fd_sc_hd__nand2_1 _09124_ (.A(_03329_),
    .B(_03330_),
    .Y(_03331_));
 sky130_fd_sc_hd__nand3_1 _09125_ (.A(_03271_),
    .B(_03328_),
    .C(_03331_),
    .Y(_03332_));
 sky130_fd_sc_hd__nand2_1 _09126_ (.A(_03271_),
    .B(_03331_),
    .Y(_03333_));
 sky130_fd_sc_hd__nand2_1 _09127_ (.A(_03333_),
    .B(_03327_),
    .Y(_03334_));
 sky130_fd_sc_hd__nand3_1 _09128_ (.A(_03082_),
    .B(_03332_),
    .C(_03334_),
    .Y(_03335_));
 sky130_fd_sc_hd__nand2_1 _09129_ (.A(_03334_),
    .B(_03332_),
    .Y(_03337_));
 sky130_fd_sc_hd__a21oi_1 _09130_ (.A1(_03036_),
    .A2(_03080_),
    .B1(_03081_),
    .Y(_03338_));
 sky130_fd_sc_hd__nand2_1 _09131_ (.A(_03337_),
    .B(_03338_),
    .Y(_03339_));
 sky130_fd_sc_hd__nand2_1 _09132_ (.A(_03078_),
    .B(_03070_),
    .Y(_03340_));
 sky130_fd_sc_hd__inv_2 _09133_ (.A(_03340_),
    .Y(_03341_));
 sky130_fd_sc_hd__nand3_1 _09134_ (.A(_03335_),
    .B(_03339_),
    .C(_03341_),
    .Y(_03342_));
 sky130_fd_sc_hd__nand2_1 _09135_ (.A(_03337_),
    .B(_03082_),
    .Y(_03343_));
 sky130_fd_sc_hd__nand3_1 _09136_ (.A(_03338_),
    .B(_03334_),
    .C(_03332_),
    .Y(_03344_));
 sky130_fd_sc_hd__nand3_1 _09137_ (.A(_03343_),
    .B(_03344_),
    .C(_03340_),
    .Y(_03345_));
 sky130_fd_sc_hd__nand2_1 _09138_ (.A(_03342_),
    .B(_03345_),
    .Y(_03346_));
 sky130_fd_sc_hd__inv_2 _09139_ (.A(_03035_),
    .Y(_03348_));
 sky130_fd_sc_hd__nand2_1 _09140_ (.A(_03032_),
    .B(_03348_),
    .Y(_03349_));
 sky130_fd_sc_hd__nand3_1 _09141_ (.A(_03035_),
    .B(_03029_),
    .C(_03031_),
    .Y(_03350_));
 sky130_fd_sc_hd__nand2_1 _09142_ (.A(_03349_),
    .B(_03350_),
    .Y(_03351_));
 sky130_fd_sc_hd__nand2_1 _09143_ (.A(_03351_),
    .B(_03080_),
    .Y(_03352_));
 sky130_fd_sc_hd__nand3_1 _09144_ (.A(_03349_),
    .B(_03350_),
    .C(_03079_),
    .Y(_03353_));
 sky130_fd_sc_hd__nand2_1 _09145_ (.A(_03352_),
    .B(_03353_),
    .Y(_03354_));
 sky130_fd_sc_hd__nand2_1 _09146_ (.A(_02749_),
    .B(_02752_),
    .Y(_03355_));
 sky130_fd_sc_hd__nor2_1 _09147_ (.A(_02752_),
    .B(_02749_),
    .Y(_03356_));
 sky130_fd_sc_hd__a21oi_1 _09148_ (.A1(_03355_),
    .A2(_02791_),
    .B1(_03356_),
    .Y(_03357_));
 sky130_fd_sc_hd__nand2_1 _09149_ (.A(_03354_),
    .B(_03357_),
    .Y(_03359_));
 sky130_fd_sc_hd__nand2_2 _09150_ (.A(_02789_),
    .B(_02784_),
    .Y(_03360_));
 sky130_fd_sc_hd__nor2_1 _09151_ (.A(_03357_),
    .B(_03354_),
    .Y(_03361_));
 sky130_fd_sc_hd__a21oi_1 _09152_ (.A1(_03359_),
    .A2(_03360_),
    .B1(_03361_),
    .Y(_03362_));
 sky130_fd_sc_hd__inv_2 _09153_ (.A(_03362_),
    .Y(_03363_));
 sky130_fd_sc_hd__nand2_1 _09154_ (.A(_03346_),
    .B(_03363_),
    .Y(_03364_));
 sky130_fd_sc_hd__nand3_1 _09155_ (.A(_03362_),
    .B(_03342_),
    .C(_03345_),
    .Y(_03365_));
 sky130_fd_sc_hd__nand2_1 _09156_ (.A(_03364_),
    .B(_03365_),
    .Y(_03366_));
 sky130_fd_sc_hd__a21o_1 _09157_ (.A1(_03355_),
    .A2(_02791_),
    .B1(_03356_),
    .X(_03367_));
 sky130_fd_sc_hd__nand3_1 _09158_ (.A(_03367_),
    .B(_03352_),
    .C(_03353_),
    .Y(_03368_));
 sky130_fd_sc_hd__inv_2 _09159_ (.A(_03360_),
    .Y(_03370_));
 sky130_fd_sc_hd__nand3_1 _09160_ (.A(_03368_),
    .B(_03359_),
    .C(_03370_),
    .Y(_03371_));
 sky130_fd_sc_hd__nand2_1 _09161_ (.A(_03354_),
    .B(_03367_),
    .Y(_03372_));
 sky130_fd_sc_hd__nand3_1 _09162_ (.A(_03357_),
    .B(_03352_),
    .C(_03353_),
    .Y(_03373_));
 sky130_fd_sc_hd__nand3_1 _09163_ (.A(_03372_),
    .B(_03373_),
    .C(_03360_),
    .Y(_03374_));
 sky130_fd_sc_hd__nand2_1 _09164_ (.A(_03371_),
    .B(_03374_),
    .Y(_03375_));
 sky130_fd_sc_hd__nand2_1 _09165_ (.A(_02794_),
    .B(_02798_),
    .Y(_03376_));
 sky130_fd_sc_hd__nor2_1 _09166_ (.A(_02798_),
    .B(_02794_),
    .Y(_03377_));
 sky130_fd_sc_hd__a21oi_2 _09167_ (.A1(_03376_),
    .A2(_02542_),
    .B1(_03377_),
    .Y(_03378_));
 sky130_fd_sc_hd__inv_2 _09168_ (.A(_03378_),
    .Y(_03379_));
 sky130_fd_sc_hd__nand2_1 _09169_ (.A(_03375_),
    .B(_03379_),
    .Y(_03381_));
 sky130_fd_sc_hd__nand2_1 _09170_ (.A(_03366_),
    .B(_03381_),
    .Y(_03382_));
 sky130_fd_sc_hd__nand3_1 _09171_ (.A(_03368_),
    .B(_03359_),
    .C(_03360_),
    .Y(_03383_));
 sky130_fd_sc_hd__nand3_1 _09172_ (.A(_03372_),
    .B(_03373_),
    .C(_03370_),
    .Y(_03384_));
 sky130_fd_sc_hd__nand2_1 _09173_ (.A(_03383_),
    .B(_03384_),
    .Y(_03385_));
 sky130_fd_sc_hd__nor2_1 _09174_ (.A(_03378_),
    .B(_03385_),
    .Y(_03386_));
 sky130_fd_sc_hd__nand3_1 _09175_ (.A(_03364_),
    .B(_03386_),
    .C(_03365_),
    .Y(_03387_));
 sky130_fd_sc_hd__nand2_1 _09176_ (.A(_03382_),
    .B(_03387_),
    .Y(_03388_));
 sky130_fd_sc_hd__inv_4 _09177_ (.A(_03388_),
    .Y(_03389_));
 sky130_fd_sc_hd__nand2_1 _09178_ (.A(_03385_),
    .B(_03378_),
    .Y(_03390_));
 sky130_fd_sc_hd__nand2_1 _09179_ (.A(_03381_),
    .B(_03390_),
    .Y(_03392_));
 sky130_fd_sc_hd__nand2_1 _09180_ (.A(_03392_),
    .B(_02805_),
    .Y(_03393_));
 sky130_fd_sc_hd__nor2_1 _09181_ (.A(_02807_),
    .B(_02806_),
    .Y(_03394_));
 sky130_fd_sc_hd__nand3_2 _09182_ (.A(_03394_),
    .B(_03381_),
    .C(_03390_),
    .Y(_03395_));
 sky130_fd_sc_hd__nand2_1 _09183_ (.A(_03393_),
    .B(_03395_),
    .Y(_03396_));
 sky130_fd_sc_hd__inv_2 _09184_ (.A(_03396_),
    .Y(_03397_));
 sky130_fd_sc_hd__nand2_1 _09185_ (.A(_03389_),
    .B(_03397_),
    .Y(_03398_));
 sky130_fd_sc_hd__nor2_1 _09186_ (.A(_02833_),
    .B(_03398_),
    .Y(_03399_));
 sky130_fd_sc_hd__nand2_1 _09187_ (.A(_02327_),
    .B(_03399_),
    .Y(_03400_));
 sky130_fd_sc_hd__nor2_1 _09188_ (.A(_00602_),
    .B(_02827_),
    .Y(_03401_));
 sky130_fd_sc_hd__nand3_1 _09189_ (.A(_02820_),
    .B(_02821_),
    .C(_03401_),
    .Y(_03403_));
 sky130_fd_sc_hd__nand2_1 _09190_ (.A(_03403_),
    .B(_02821_),
    .Y(_03404_));
 sky130_fd_sc_hd__nor2_1 _09191_ (.A(_03396_),
    .B(_03388_),
    .Y(_03405_));
 sky130_fd_sc_hd__inv_2 _09192_ (.A(_03395_),
    .Y(_03406_));
 sky130_fd_sc_hd__nand3_1 _09193_ (.A(_03406_),
    .B(_03382_),
    .C(_03387_),
    .Y(_03407_));
 sky130_fd_sc_hd__nand2_1 _09194_ (.A(_03407_),
    .B(_03387_),
    .Y(_03408_));
 sky130_fd_sc_hd__a21oi_1 _09195_ (.A1(_03404_),
    .A2(_03405_),
    .B1(_03408_),
    .Y(_03409_));
 sky130_fd_sc_hd__nand2_1 _09196_ (.A(_03400_),
    .B(_03409_),
    .Y(_03410_));
 sky130_fd_sc_hd__a21oi_2 _09197_ (.A1(_03220_),
    .A2(_03218_),
    .B1(_03219_),
    .Y(_03411_));
 sky130_fd_sc_hd__nand2_1 _09198_ (.A(_04876_),
    .B(_05031_),
    .Y(_03412_));
 sky130_fd_sc_hd__and4_1 _09199_ (.A(_04873_),
    .B(_04871_),
    .C(_03160_),
    .D(_03182_),
    .X(_03414_));
 sky130_fd_sc_hd__inv_2 _09200_ (.A(_03414_),
    .Y(_03415_));
 sky130_fd_sc_hd__a22o_1 _09201_ (.A1(_04873_),
    .A2(_03160_),
    .B1(_04871_),
    .B2(_03182_),
    .X(_03416_));
 sky130_fd_sc_hd__nand2_1 _09202_ (.A(_03415_),
    .B(_03416_),
    .Y(_03417_));
 sky130_fd_sc_hd__or2_1 _09203_ (.A(_03412_),
    .B(_03417_),
    .X(_03418_));
 sky130_fd_sc_hd__nand2_1 _09204_ (.A(_03417_),
    .B(_03412_),
    .Y(_03419_));
 sky130_fd_sc_hd__nand2_1 _09205_ (.A(_03418_),
    .B(_03419_),
    .Y(_03420_));
 sky130_fd_sc_hd__inv_2 _09206_ (.A(_03420_),
    .Y(_03421_));
 sky130_fd_sc_hd__or2_1 _09207_ (.A(_03411_),
    .B(_03421_),
    .X(_03422_));
 sky130_fd_sc_hd__nand2_1 _09208_ (.A(_03421_),
    .B(_03411_),
    .Y(_03423_));
 sky130_fd_sc_hd__nand2_1 _09209_ (.A(_00529_),
    .B(_00656_),
    .Y(_03425_));
 sky130_fd_sc_hd__and4_1 _09210_ (.A(net46),
    .B(_00124_),
    .C(_05028_),
    .D(_04928_),
    .X(_03426_));
 sky130_fd_sc_hd__a22o_1 _09211_ (.A1(net46),
    .A2(_05028_),
    .B1(_00124_),
    .B2(_04928_),
    .X(_03427_));
 sky130_fd_sc_hd__and2b_1 _09212_ (.A_N(_03426_),
    .B(_03427_),
    .X(_03428_));
 sky130_fd_sc_hd__xor2_1 _09213_ (.A(_03425_),
    .B(_03428_),
    .X(_03429_));
 sky130_fd_sc_hd__a21o_1 _09214_ (.A1(_03422_),
    .A2(_03423_),
    .B1(_03429_),
    .X(_03430_));
 sky130_fd_sc_hd__nand3_1 _09215_ (.A(_03422_),
    .B(_03429_),
    .C(_03423_),
    .Y(_03431_));
 sky130_fd_sc_hd__nand2_1 _09216_ (.A(_03430_),
    .B(_03431_),
    .Y(_03432_));
 sky130_fd_sc_hd__nand2_1 _09217_ (.A(_03205_),
    .B(_03203_),
    .Y(_03433_));
 sky130_fd_sc_hd__inv_2 _09218_ (.A(_03433_),
    .Y(_03434_));
 sky130_fd_sc_hd__nand2_1 _09219_ (.A(_04818_),
    .B(_02049_),
    .Y(_03436_));
 sky130_fd_sc_hd__and4_1 _09220_ (.A(_04812_),
    .B(_04808_),
    .C(_02544_),
    .D(_01873_),
    .X(_03437_));
 sky130_fd_sc_hd__a22o_1 _09221_ (.A1(_04812_),
    .A2(_02544_),
    .B1(_04808_),
    .B2(_01873_),
    .X(_03438_));
 sky130_fd_sc_hd__nand2b_1 _09222_ (.A_N(_03437_),
    .B(_03438_),
    .Y(_03439_));
 sky130_fd_sc_hd__or2_1 _09223_ (.A(_03436_),
    .B(_03439_),
    .X(_03440_));
 sky130_fd_sc_hd__nand2_1 _09224_ (.A(_03439_),
    .B(_03436_),
    .Y(_03441_));
 sky130_fd_sc_hd__nand2_1 _09225_ (.A(_03440_),
    .B(_03441_),
    .Y(_03442_));
 sky130_fd_sc_hd__inv_2 _09226_ (.A(_01037_),
    .Y(_03443_));
 sky130_fd_sc_hd__nor3_1 _09227_ (.A(_01330_),
    .B(_03443_),
    .C(_03154_),
    .Y(_03444_));
 sky130_fd_sc_hd__inv_2 _09228_ (.A(_03444_),
    .Y(_03445_));
 sky130_fd_sc_hd__nand3_1 _09229_ (.A(_03442_),
    .B(_03445_),
    .C(_03158_),
    .Y(_03447_));
 sky130_fd_sc_hd__nand2_1 _09230_ (.A(_03158_),
    .B(_03445_),
    .Y(_03448_));
 sky130_fd_sc_hd__nand3_1 _09231_ (.A(_03440_),
    .B(_03441_),
    .C(_03448_),
    .Y(_03449_));
 sky130_fd_sc_hd__nand2_1 _09232_ (.A(_03447_),
    .B(_03449_),
    .Y(_03450_));
 sky130_fd_sc_hd__inv_2 _09233_ (.A(_03198_),
    .Y(_03451_));
 sky130_fd_sc_hd__nor2_1 _09234_ (.A(_03194_),
    .B(_03451_),
    .Y(_03452_));
 sky130_fd_sc_hd__nand2_1 _09235_ (.A(_03450_),
    .B(_03452_),
    .Y(_03453_));
 sky130_fd_sc_hd__nand3b_1 _09236_ (.A_N(_03452_),
    .B(_03447_),
    .C(_03449_),
    .Y(_03454_));
 sky130_fd_sc_hd__nand2_1 _09237_ (.A(_03453_),
    .B(_03454_),
    .Y(_03455_));
 sky130_fd_sc_hd__or2_1 _09238_ (.A(_03434_),
    .B(_03455_),
    .X(_03456_));
 sky130_fd_sc_hd__nand2_1 _09239_ (.A(_03455_),
    .B(_03434_),
    .Y(_03458_));
 sky130_fd_sc_hd__nand3b_1 _09240_ (.A_N(_03432_),
    .B(_03456_),
    .C(_03458_),
    .Y(_03459_));
 sky130_fd_sc_hd__or2_1 _09241_ (.A(_03433_),
    .B(_03455_),
    .X(_03460_));
 sky130_fd_sc_hd__nand2_1 _09242_ (.A(_03455_),
    .B(_03433_),
    .Y(_03461_));
 sky130_fd_sc_hd__nand3_1 _09243_ (.A(_03460_),
    .B(_03461_),
    .C(_03432_),
    .Y(_03462_));
 sky130_fd_sc_hd__nand2_1 _09244_ (.A(_03459_),
    .B(_03462_),
    .Y(_03463_));
 sky130_fd_sc_hd__o21a_2 _09245_ (.A1(_03178_),
    .A2(_03151_),
    .B1(_03183_),
    .X(_03464_));
 sky130_fd_sc_hd__inv_2 _09246_ (.A(_03464_),
    .Y(_03465_));
 sky130_fd_sc_hd__nand2_1 _09247_ (.A(_03463_),
    .B(_03465_),
    .Y(_03466_));
 sky130_fd_sc_hd__nand3_1 _09248_ (.A(_03459_),
    .B(_03462_),
    .C(_03464_),
    .Y(_03467_));
 sky130_fd_sc_hd__nand2_1 _09249_ (.A(_03466_),
    .B(_03467_),
    .Y(_03469_));
 sky130_fd_sc_hd__o21ai_2 _09250_ (.A1(_03211_),
    .A2(_03208_),
    .B1(_03244_),
    .Y(_03470_));
 sky130_fd_sc_hd__nand2_1 _09251_ (.A(_03469_),
    .B(_03470_),
    .Y(_03471_));
 sky130_fd_sc_hd__nand3b_1 _09252_ (.A_N(_03470_),
    .B(_03466_),
    .C(_03467_),
    .Y(_03472_));
 sky130_fd_sc_hd__nand2_1 _09253_ (.A(_03471_),
    .B(_03472_),
    .Y(_03473_));
 sky130_fd_sc_hd__inv_2 _09254_ (.A(_03473_),
    .Y(_03474_));
 sky130_fd_sc_hd__nand2_1 _09255_ (.A(_01535_),
    .B(net19),
    .Y(_03475_));
 sky130_fd_sc_hd__and4_1 _09256_ (.A(_02379_),
    .B(_02357_),
    .C(net20),
    .D(net21),
    .X(_03476_));
 sky130_fd_sc_hd__a22o_1 _09257_ (.A1(_02379_),
    .A2(net21),
    .B1(_02357_),
    .B2(net20),
    .X(_03477_));
 sky130_fd_sc_hd__nand2b_1 _09258_ (.A_N(_03476_),
    .B(_03477_),
    .Y(_03478_));
 sky130_fd_sc_hd__or2_1 _09259_ (.A(_03475_),
    .B(_03478_),
    .X(_03480_));
 sky130_fd_sc_hd__nand2_1 _09260_ (.A(_03478_),
    .B(_03475_),
    .Y(_03481_));
 sky130_fd_sc_hd__nand2_1 _09261_ (.A(_03480_),
    .B(_03481_),
    .Y(_03482_));
 sky130_fd_sc_hd__nand2_1 _09262_ (.A(_03095_),
    .B(_03090_),
    .Y(_03483_));
 sky130_fd_sc_hd__inv_2 _09263_ (.A(_03483_),
    .Y(_03484_));
 sky130_fd_sc_hd__nand2_1 _09264_ (.A(_03482_),
    .B(_03484_),
    .Y(_03485_));
 sky130_fd_sc_hd__nand3_2 _09265_ (.A(_03480_),
    .B(_03483_),
    .C(_03481_),
    .Y(_03486_));
 sky130_fd_sc_hd__nand2_1 _09266_ (.A(_03485_),
    .B(_03486_),
    .Y(_03487_));
 sky130_fd_sc_hd__nand2_1 _09267_ (.A(_01565_),
    .B(_00393_),
    .Y(_03488_));
 sky130_fd_sc_hd__inv_2 _09268_ (.A(net18),
    .Y(_03489_));
 sky130_fd_sc_hd__nand2_1 _09269_ (.A(_04260_),
    .B(net17),
    .Y(_03491_));
 sky130_fd_sc_hd__nor3_1 _09270_ (.A(_02086_),
    .B(_03489_),
    .C(_03491_),
    .Y(_03492_));
 sky130_fd_sc_hd__o21ai_1 _09271_ (.A1(_02086_),
    .A2(_03489_),
    .B1(_03491_),
    .Y(_03493_));
 sky130_fd_sc_hd__and2b_1 _09272_ (.A_N(_03492_),
    .B(_03493_),
    .X(_03494_));
 sky130_fd_sc_hd__xor2_1 _09273_ (.A(_03488_),
    .B(_03494_),
    .X(_03495_));
 sky130_fd_sc_hd__nand2_1 _09274_ (.A(_03487_),
    .B(_03495_),
    .Y(_03496_));
 sky130_fd_sc_hd__nand3b_1 _09275_ (.A_N(_03495_),
    .B(_03485_),
    .C(_03486_),
    .Y(_03497_));
 sky130_fd_sc_hd__nand2_1 _09276_ (.A(_03496_),
    .B(_03497_),
    .Y(_03498_));
 sky130_fd_sc_hd__nand2_1 _09277_ (.A(_03112_),
    .B(_03100_),
    .Y(_03499_));
 sky130_fd_sc_hd__nand2b_1 _09278_ (.A_N(_03498_),
    .B(_03499_),
    .Y(_03500_));
 sky130_fd_sc_hd__nand2b_1 _09279_ (.A_N(_03499_),
    .B(_03498_),
    .Y(_03502_));
 sky130_fd_sc_hd__nand2_1 _09280_ (.A(_03500_),
    .B(_03502_),
    .Y(_03503_));
 sky130_fd_sc_hd__nand2_1 _09281_ (.A(_01323_),
    .B(_00003_),
    .Y(_03504_));
 sky130_fd_sc_hd__and4_1 _09282_ (.A(_00204_),
    .B(_00412_),
    .C(_04084_),
    .D(_05160_),
    .X(_03505_));
 sky130_fd_sc_hd__a22o_1 _09283_ (.A1(_00204_),
    .A2(_05160_),
    .B1(_00412_),
    .B2(_04084_),
    .X(_03506_));
 sky130_fd_sc_hd__nand2b_1 _09284_ (.A_N(_03505_),
    .B(_03506_),
    .Y(_03507_));
 sky130_fd_sc_hd__or2_1 _09285_ (.A(_03504_),
    .B(_03507_),
    .X(_03508_));
 sky130_fd_sc_hd__nand2_1 _09286_ (.A(_03507_),
    .B(_03504_),
    .Y(_03509_));
 sky130_fd_sc_hd__nand2_1 _09287_ (.A(_03508_),
    .B(_03509_),
    .Y(_03510_));
 sky130_fd_sc_hd__inv_2 _09288_ (.A(net17),
    .Y(_03511_));
 sky130_fd_sc_hd__nor3_1 _09289_ (.A(_02086_),
    .B(_03511_),
    .C(_03104_),
    .Y(_03513_));
 sky130_fd_sc_hd__inv_2 _09290_ (.A(_03513_),
    .Y(_03514_));
 sky130_fd_sc_hd__nand2_1 _09291_ (.A(_03109_),
    .B(_03514_),
    .Y(_03515_));
 sky130_fd_sc_hd__nand2_1 _09292_ (.A(_03510_),
    .B(_03515_),
    .Y(_03516_));
 sky130_fd_sc_hd__inv_2 _09293_ (.A(_03515_),
    .Y(_03517_));
 sky130_fd_sc_hd__nand3_1 _09294_ (.A(_03508_),
    .B(_03509_),
    .C(_03517_),
    .Y(_03518_));
 sky130_fd_sc_hd__inv_2 _09295_ (.A(_04084_),
    .Y(_03519_));
 sky130_fd_sc_hd__nor3_1 _09296_ (.A(_01937_),
    .B(_03519_),
    .C(_03125_),
    .Y(_03520_));
 sky130_fd_sc_hd__inv_2 _09297_ (.A(_03130_),
    .Y(_03521_));
 sky130_fd_sc_hd__nor2_1 _09298_ (.A(_03520_),
    .B(_03521_),
    .Y(_03522_));
 sky130_fd_sc_hd__a21o_1 _09299_ (.A1(_03516_),
    .A2(_03518_),
    .B1(_03522_),
    .X(_03524_));
 sky130_fd_sc_hd__nand3_1 _09300_ (.A(_03516_),
    .B(_03522_),
    .C(_03518_),
    .Y(_03525_));
 sky130_fd_sc_hd__nand2_1 _09301_ (.A(_03524_),
    .B(_03525_),
    .Y(_03526_));
 sky130_fd_sc_hd__nand2_1 _09302_ (.A(_03503_),
    .B(_03526_),
    .Y(_03527_));
 sky130_fd_sc_hd__inv_2 _09303_ (.A(_03526_),
    .Y(_03528_));
 sky130_fd_sc_hd__nand3_1 _09304_ (.A(_03500_),
    .B(_03502_),
    .C(_03528_),
    .Y(_03529_));
 sky130_fd_sc_hd__nand2_1 _09305_ (.A(_03527_),
    .B(_03529_),
    .Y(_03530_));
 sky130_fd_sc_hd__and2_1 _09306_ (.A(_03142_),
    .B(_03118_),
    .X(_03531_));
 sky130_fd_sc_hd__nand2_1 _09307_ (.A(_03530_),
    .B(_03531_),
    .Y(_03532_));
 sky130_fd_sc_hd__nand3b_2 _09308_ (.A_N(_03531_),
    .B(_03527_),
    .C(_03529_),
    .Y(_03533_));
 sky130_fd_sc_hd__nand2_1 _09309_ (.A(_03532_),
    .B(_03533_),
    .Y(_03535_));
 sky130_fd_sc_hd__o21a_1 _09310_ (.A1(_03163_),
    .A2(_03164_),
    .B1(_03167_),
    .X(_03536_));
 sky130_fd_sc_hd__nand2_1 _09311_ (.A(_03215_),
    .B(_00850_),
    .Y(_03537_));
 sky130_fd_sc_hd__inv_2 _09312_ (.A(_03537_),
    .Y(_03538_));
 sky130_fd_sc_hd__and4_1 _09313_ (.A(_00784_),
    .B(_00740_),
    .C(_05032_),
    .D(_02995_),
    .X(_03539_));
 sky130_fd_sc_hd__inv_2 _09314_ (.A(_03539_),
    .Y(_03540_));
 sky130_fd_sc_hd__a22o_1 _09315_ (.A1(_00784_),
    .A2(_05032_),
    .B1(_00740_),
    .B2(_05029_),
    .X(_03541_));
 sky130_fd_sc_hd__and2_1 _09316_ (.A(_03540_),
    .B(_03541_),
    .X(_03542_));
 sky130_fd_sc_hd__or2_1 _09317_ (.A(_03538_),
    .B(_03542_),
    .X(_03543_));
 sky130_fd_sc_hd__nand2_1 _09318_ (.A(_03542_),
    .B(_03538_),
    .Y(_03544_));
 sky130_fd_sc_hd__nand2_1 _09319_ (.A(_03543_),
    .B(_03544_),
    .Y(_03546_));
 sky130_fd_sc_hd__nor2_1 _09320_ (.A(_03536_),
    .B(_03546_),
    .Y(_03547_));
 sky130_fd_sc_hd__nand2_1 _09321_ (.A(_03546_),
    .B(_03536_),
    .Y(_03548_));
 sky130_fd_sc_hd__inv_2 _09322_ (.A(_03548_),
    .Y(_03549_));
 sky130_fd_sc_hd__nand2_1 _09323_ (.A(_03809_),
    .B(_01147_),
    .Y(_03550_));
 sky130_fd_sc_hd__and4_1 _09324_ (.A(_04964_),
    .B(_04962_),
    .C(_01081_),
    .D(_01037_),
    .X(_03551_));
 sky130_fd_sc_hd__a22o_1 _09325_ (.A1(_04964_),
    .A2(_01081_),
    .B1(_04962_),
    .B2(_01037_),
    .X(_03552_));
 sky130_fd_sc_hd__and2b_1 _09326_ (.A_N(_03551_),
    .B(_03552_),
    .X(_03553_));
 sky130_fd_sc_hd__xor2_1 _09327_ (.A(_03550_),
    .B(_03553_),
    .X(_03554_));
 sky130_fd_sc_hd__o21ai_1 _09328_ (.A1(_03547_),
    .A2(_03549_),
    .B1(_03554_),
    .Y(_03555_));
 sky130_fd_sc_hd__inv_2 _09329_ (.A(_03554_),
    .Y(_03557_));
 sky130_fd_sc_hd__nand3b_1 _09330_ (.A_N(_03547_),
    .B(_03557_),
    .C(_03548_),
    .Y(_03558_));
 sky130_fd_sc_hd__nand2_1 _09331_ (.A(_03555_),
    .B(_03558_),
    .Y(_03559_));
 sky130_fd_sc_hd__nand2_1 _09332_ (.A(_03134_),
    .B(_03132_),
    .Y(_03560_));
 sky130_fd_sc_hd__nand2_1 _09333_ (.A(_03559_),
    .B(_03560_),
    .Y(_03561_));
 sky130_fd_sc_hd__inv_2 _09334_ (.A(_03560_),
    .Y(_03562_));
 sky130_fd_sc_hd__nand3_1 _09335_ (.A(_03555_),
    .B(_03558_),
    .C(_03562_),
    .Y(_03563_));
 sky130_fd_sc_hd__nand2_1 _09336_ (.A(_03561_),
    .B(_03563_),
    .Y(_03564_));
 sky130_fd_sc_hd__nand2_1 _09337_ (.A(_03173_),
    .B(_03172_),
    .Y(_03565_));
 sky130_fd_sc_hd__nand2_1 _09338_ (.A(_03564_),
    .B(_03565_),
    .Y(_03566_));
 sky130_fd_sc_hd__nand3b_1 _09339_ (.A_N(_03565_),
    .B(_03561_),
    .C(_03563_),
    .Y(_03568_));
 sky130_fd_sc_hd__nand2_1 _09340_ (.A(_03566_),
    .B(_03568_),
    .Y(_03569_));
 sky130_fd_sc_hd__nand2_1 _09341_ (.A(_03535_),
    .B(_03569_),
    .Y(_03570_));
 sky130_fd_sc_hd__inv_2 _09342_ (.A(_03569_),
    .Y(_03571_));
 sky130_fd_sc_hd__nand3_2 _09343_ (.A(_03571_),
    .B(_03532_),
    .C(_03533_),
    .Y(_03572_));
 sky130_fd_sc_hd__nand2_1 _09344_ (.A(_03570_),
    .B(_03572_),
    .Y(_03573_));
 sky130_fd_sc_hd__and2_1 _09345_ (.A(_03187_),
    .B(_03143_),
    .X(_03574_));
 sky130_fd_sc_hd__nand2_1 _09346_ (.A(_03573_),
    .B(_03574_),
    .Y(_03575_));
 sky130_fd_sc_hd__nand3b_2 _09347_ (.A_N(_03574_),
    .B(_03570_),
    .C(_03572_),
    .Y(_03576_));
 sky130_fd_sc_hd__nand3_1 _09348_ (.A(_03474_),
    .B(_03575_),
    .C(_03576_),
    .Y(_03577_));
 sky130_fd_sc_hd__nand2_1 _09349_ (.A(_03575_),
    .B(_03576_),
    .Y(_03579_));
 sky130_fd_sc_hd__nand2_1 _09350_ (.A(_03579_),
    .B(_03473_),
    .Y(_03580_));
 sky130_fd_sc_hd__nand2_1 _09351_ (.A(_03577_),
    .B(_03580_),
    .Y(_03581_));
 sky130_fd_sc_hd__and2_1 _09352_ (.A(_03267_),
    .B(_03188_),
    .X(_03582_));
 sky130_fd_sc_hd__nand2_1 _09353_ (.A(_03581_),
    .B(_03582_),
    .Y(_03583_));
 sky130_fd_sc_hd__nand3b_2 _09354_ (.A_N(_03582_),
    .B(_03577_),
    .C(_03580_),
    .Y(_03584_));
 sky130_fd_sc_hd__nand2_1 _09355_ (.A(_03583_),
    .B(_03584_),
    .Y(_03585_));
 sky130_fd_sc_hd__nor2_1 _09356_ (.A(_03228_),
    .B(_03224_),
    .Y(_03586_));
 sky130_fd_sc_hd__inv_2 _09357_ (.A(_03240_),
    .Y(_03587_));
 sky130_fd_sc_hd__inv_2 _09358_ (.A(_03233_),
    .Y(_03588_));
 sky130_fd_sc_hd__o21a_1 _09359_ (.A1(_03231_),
    .A2(_03235_),
    .B1(_03588_),
    .X(_03590_));
 sky130_fd_sc_hd__inv_2 _09360_ (.A(_03590_),
    .Y(_03591_));
 sky130_fd_sc_hd__and4_1 _09361_ (.A(net49),
    .B(net50),
    .C(_04809_),
    .D(_04819_),
    .X(_03592_));
 sky130_fd_sc_hd__inv_2 _09362_ (.A(_03592_),
    .Y(_03593_));
 sky130_fd_sc_hd__a22o_1 _09363_ (.A1(net49),
    .A2(_00254_),
    .B1(net50),
    .B2(_00522_),
    .X(_03594_));
 sky130_fd_sc_hd__nand2_1 _09364_ (.A(_03593_),
    .B(_03594_),
    .Y(_03595_));
 sky130_fd_sc_hd__inv_2 _09365_ (.A(_03595_),
    .Y(_03596_));
 sky130_fd_sc_hd__nand2_1 _09366_ (.A(net51),
    .B(_04828_),
    .Y(_03597_));
 sky130_fd_sc_hd__inv_2 _09367_ (.A(_03597_),
    .Y(_03598_));
 sky130_fd_sc_hd__nand2_1 _09368_ (.A(_03596_),
    .B(_03598_),
    .Y(_03599_));
 sky130_fd_sc_hd__nand2_1 _09369_ (.A(_03595_),
    .B(_03597_),
    .Y(_03601_));
 sky130_fd_sc_hd__nand2_1 _09370_ (.A(_03599_),
    .B(_03601_),
    .Y(_03602_));
 sky130_fd_sc_hd__or2_1 _09371_ (.A(_03591_),
    .B(_03602_),
    .X(_03603_));
 sky130_fd_sc_hd__nand2_1 _09372_ (.A(_03602_),
    .B(_03591_),
    .Y(_03604_));
 sky130_fd_sc_hd__a21oi_1 _09373_ (.A1(_03278_),
    .A2(_03275_),
    .B1(_03277_),
    .Y(_03605_));
 sky130_fd_sc_hd__a21o_1 _09374_ (.A1(_03603_),
    .A2(_03604_),
    .B1(_03605_),
    .X(_03606_));
 sky130_fd_sc_hd__nand3_1 _09375_ (.A(_03603_),
    .B(_03605_),
    .C(_03604_),
    .Y(_03607_));
 sky130_fd_sc_hd__nand2_1 _09376_ (.A(_03606_),
    .B(_03607_),
    .Y(_03608_));
 sky130_fd_sc_hd__o21ai_1 _09377_ (.A1(_03586_),
    .A2(_03587_),
    .B1(_03608_),
    .Y(_03609_));
 sky130_fd_sc_hd__nor2_1 _09378_ (.A(_03586_),
    .B(_03587_),
    .Y(_03610_));
 sky130_fd_sc_hd__nand3_1 _09379_ (.A(_03610_),
    .B(_03606_),
    .C(_03607_),
    .Y(_03612_));
 sky130_fd_sc_hd__nand2_1 _09380_ (.A(_03609_),
    .B(_03612_),
    .Y(_03613_));
 sky130_fd_sc_hd__nand2_1 _09381_ (.A(_03291_),
    .B(_03290_),
    .Y(_03614_));
 sky130_fd_sc_hd__nand2_1 _09382_ (.A(_03613_),
    .B(_03614_),
    .Y(_03615_));
 sky130_fd_sc_hd__nand3b_1 _09383_ (.A_N(_03614_),
    .B(_03609_),
    .C(_03612_),
    .Y(_03616_));
 sky130_fd_sc_hd__nand2_1 _09384_ (.A(_03615_),
    .B(_03616_),
    .Y(_03617_));
 sky130_fd_sc_hd__nand2_1 _09385_ (.A(_03304_),
    .B(_03295_),
    .Y(_03618_));
 sky130_fd_sc_hd__nand2_1 _09386_ (.A(_03617_),
    .B(_03618_),
    .Y(_03619_));
 sky130_fd_sc_hd__inv_2 _09387_ (.A(_03618_),
    .Y(_03620_));
 sky130_fd_sc_hd__nand3_1 _09388_ (.A(_03615_),
    .B(_03616_),
    .C(_03620_),
    .Y(_03621_));
 sky130_fd_sc_hd__nand2_1 _09389_ (.A(_03619_),
    .B(_03621_),
    .Y(_03623_));
 sky130_fd_sc_hd__inv_2 _09390_ (.A(net52),
    .Y(_03624_));
 sky130_fd_sc_hd__inv_2 _09391_ (.A(net53),
    .Y(_03625_));
 sky130_fd_sc_hd__or4_2 _09392_ (.A(_03624_),
    .B(_03625_),
    .C(_00264_),
    .D(_01956_),
    .X(_03626_));
 sky130_fd_sc_hd__a22o_1 _09393_ (.A1(net52),
    .A2(_04991_),
    .B1(net53),
    .B2(_04992_),
    .X(_03627_));
 sky130_fd_sc_hd__nand2_1 _09394_ (.A(_03626_),
    .B(_03627_),
    .Y(_03628_));
 sky130_fd_sc_hd__inv_2 _09395_ (.A(_03628_),
    .Y(_03629_));
 sky130_fd_sc_hd__nand2_1 _09396_ (.A(_03623_),
    .B(_03629_),
    .Y(_03630_));
 sky130_fd_sc_hd__nand3_1 _09397_ (.A(_03619_),
    .B(_03621_),
    .C(_03628_),
    .Y(_03631_));
 sky130_fd_sc_hd__nand2_1 _09398_ (.A(_03630_),
    .B(_03631_),
    .Y(_03632_));
 sky130_fd_sc_hd__nor2_1 _09399_ (.A(_03250_),
    .B(_03246_),
    .Y(_03634_));
 sky130_fd_sc_hd__inv_2 _09400_ (.A(_03260_),
    .Y(_03635_));
 sky130_fd_sc_hd__nor2_2 _09401_ (.A(_03634_),
    .B(_03635_),
    .Y(_03636_));
 sky130_fd_sc_hd__inv_2 _09402_ (.A(_03636_),
    .Y(_03637_));
 sky130_fd_sc_hd__nand2_1 _09403_ (.A(_03632_),
    .B(_03637_),
    .Y(_03638_));
 sky130_fd_sc_hd__nand3_1 _09404_ (.A(_03630_),
    .B(_03631_),
    .C(_03636_),
    .Y(_03639_));
 sky130_fd_sc_hd__nand2_1 _09405_ (.A(_03638_),
    .B(_03639_),
    .Y(_03640_));
 sky130_fd_sc_hd__nand2_1 _09406_ (.A(_03313_),
    .B(_03309_),
    .Y(_03641_));
 sky130_fd_sc_hd__nand2_1 _09407_ (.A(_03640_),
    .B(_03641_),
    .Y(_03642_));
 sky130_fd_sc_hd__nand3b_1 _09408_ (.A_N(_03641_),
    .B(_03638_),
    .C(_03639_),
    .Y(_03643_));
 sky130_fd_sc_hd__nand2_1 _09409_ (.A(_03642_),
    .B(_03643_),
    .Y(_03645_));
 sky130_fd_sc_hd__nand2_1 _09410_ (.A(_03585_),
    .B(_03645_),
    .Y(_03646_));
 sky130_fd_sc_hd__inv_2 _09411_ (.A(_03645_),
    .Y(_03647_));
 sky130_fd_sc_hd__nand3_2 _09412_ (.A(_03647_),
    .B(_03583_),
    .C(_03584_),
    .Y(_03648_));
 sky130_fd_sc_hd__nand2_1 _09413_ (.A(_03646_),
    .B(_03648_),
    .Y(_03649_));
 sky130_fd_sc_hd__and2_1 _09414_ (.A(_03332_),
    .B(_03271_),
    .X(_03650_));
 sky130_fd_sc_hd__nand2_1 _09415_ (.A(_03649_),
    .B(_03650_),
    .Y(_03651_));
 sky130_fd_sc_hd__nand3b_1 _09416_ (.A_N(_03650_),
    .B(_03646_),
    .C(_03648_),
    .Y(_03652_));
 sky130_fd_sc_hd__nand2_1 _09417_ (.A(_03651_),
    .B(_03652_),
    .Y(_03653_));
 sky130_fd_sc_hd__nand2_1 _09418_ (.A(_03326_),
    .B(_03321_),
    .Y(_03654_));
 sky130_fd_sc_hd__inv_2 _09419_ (.A(_03654_),
    .Y(_03656_));
 sky130_fd_sc_hd__nand2_1 _09420_ (.A(_03653_),
    .B(_03656_),
    .Y(_03657_));
 sky130_fd_sc_hd__nand3_1 _09421_ (.A(_03651_),
    .B(_03652_),
    .C(_03654_),
    .Y(_03658_));
 sky130_fd_sc_hd__nand2_1 _09422_ (.A(_03657_),
    .B(_03658_),
    .Y(_03659_));
 sky130_fd_sc_hd__a21o_1 _09423_ (.A1(_03343_),
    .A2(_03344_),
    .B1(_03341_),
    .X(_03660_));
 sky130_fd_sc_hd__nand2_1 _09424_ (.A(_03660_),
    .B(_03335_),
    .Y(_03661_));
 sky130_fd_sc_hd__inv_2 _09425_ (.A(_03661_),
    .Y(_03662_));
 sky130_fd_sc_hd__nand2_1 _09426_ (.A(_03659_),
    .B(_03662_),
    .Y(_03663_));
 sky130_fd_sc_hd__nand3_1 _09427_ (.A(_03657_),
    .B(_03658_),
    .C(_03661_),
    .Y(_03664_));
 sky130_fd_sc_hd__nand2_1 _09428_ (.A(_03663_),
    .B(_03664_),
    .Y(_03665_));
 sky130_fd_sc_hd__nand2_1 _09429_ (.A(_03665_),
    .B(_03364_),
    .Y(_03667_));
 sky130_fd_sc_hd__inv_2 _09430_ (.A(_03364_),
    .Y(_03668_));
 sky130_fd_sc_hd__nand3_1 _09431_ (.A(_03663_),
    .B(_03668_),
    .C(_03664_),
    .Y(_03669_));
 sky130_fd_sc_hd__nand2_1 _09432_ (.A(_03667_),
    .B(_03669_),
    .Y(_03670_));
 sky130_fd_sc_hd__nand2_1 _09433_ (.A(_03577_),
    .B(_03576_),
    .Y(_03671_));
 sky130_fd_sc_hd__inv_2 _09434_ (.A(_03488_),
    .Y(_03672_));
 sky130_fd_sc_hd__a21oi_1 _09435_ (.A1(_03493_),
    .A2(_03672_),
    .B1(_03492_),
    .Y(_03673_));
 sky130_fd_sc_hd__inv_2 _09436_ (.A(_03673_),
    .Y(_03674_));
 sky130_fd_sc_hd__nand2_1 _09437_ (.A(_00003_),
    .B(_04084_),
    .Y(_03675_));
 sky130_fd_sc_hd__and4_1 _09438_ (.A(_00204_),
    .B(_00412_),
    .C(_05160_),
    .D(_00393_),
    .X(_03676_));
 sky130_fd_sc_hd__inv_2 _09439_ (.A(_03676_),
    .Y(_03678_));
 sky130_fd_sc_hd__a22o_1 _09440_ (.A1(_00204_),
    .A2(_00393_),
    .B1(_00412_),
    .B2(_05160_),
    .X(_03679_));
 sky130_fd_sc_hd__nand2_1 _09441_ (.A(_03678_),
    .B(_03679_),
    .Y(_03680_));
 sky130_fd_sc_hd__or2_1 _09442_ (.A(_03675_),
    .B(_03680_),
    .X(_03681_));
 sky130_fd_sc_hd__nand2_1 _09443_ (.A(_03680_),
    .B(_03675_),
    .Y(_03682_));
 sky130_fd_sc_hd__nand2_1 _09444_ (.A(_03681_),
    .B(_03682_),
    .Y(_03683_));
 sky130_fd_sc_hd__or2_1 _09445_ (.A(_03674_),
    .B(_03683_),
    .X(_03684_));
 sky130_fd_sc_hd__nand2_1 _09446_ (.A(_03683_),
    .B(_03674_),
    .Y(_03685_));
 sky130_fd_sc_hd__inv_2 _09447_ (.A(_03508_),
    .Y(_03686_));
 sky130_fd_sc_hd__nor2_1 _09448_ (.A(_03505_),
    .B(_03686_),
    .Y(_03687_));
 sky130_fd_sc_hd__a21oi_1 _09449_ (.A1(_03684_),
    .A2(_03685_),
    .B1(_03687_),
    .Y(_03689_));
 sky130_fd_sc_hd__inv_2 _09450_ (.A(_03689_),
    .Y(_03690_));
 sky130_fd_sc_hd__nand3_1 _09451_ (.A(_03684_),
    .B(_03687_),
    .C(_03685_),
    .Y(_03691_));
 sky130_fd_sc_hd__nand2_1 _09452_ (.A(_03690_),
    .B(_03691_),
    .Y(_03692_));
 sky130_fd_sc_hd__nand2_1 _09453_ (.A(_01535_),
    .B(net20),
    .Y(_03693_));
 sky130_fd_sc_hd__and4_1 _09454_ (.A(_02379_),
    .B(_02357_),
    .C(net21),
    .D(net22),
    .X(_03694_));
 sky130_fd_sc_hd__a22o_1 _09455_ (.A1(_02379_),
    .A2(net22),
    .B1(_02357_),
    .B2(net21),
    .X(_03695_));
 sky130_fd_sc_hd__nand2b_1 _09456_ (.A_N(_03694_),
    .B(_03695_),
    .Y(_03696_));
 sky130_fd_sc_hd__or2_1 _09457_ (.A(_03693_),
    .B(_03696_),
    .X(_03697_));
 sky130_fd_sc_hd__nand2_1 _09458_ (.A(_03696_),
    .B(_03693_),
    .Y(_03698_));
 sky130_fd_sc_hd__a31o_1 _09459_ (.A1(_03477_),
    .A2(_01535_),
    .A3(net19),
    .B1(_03476_),
    .X(_03700_));
 sky130_fd_sc_hd__a21o_1 _09460_ (.A1(_03697_),
    .A2(_03698_),
    .B1(_03700_),
    .X(_03701_));
 sky130_fd_sc_hd__nand3_2 _09461_ (.A(_03697_),
    .B(_03700_),
    .C(_03698_),
    .Y(_03702_));
 sky130_fd_sc_hd__nand2_1 _09462_ (.A(_03701_),
    .B(_03702_),
    .Y(_03703_));
 sky130_fd_sc_hd__nand2_1 _09463_ (.A(_01565_),
    .B(net17),
    .Y(_03704_));
 sky130_fd_sc_hd__and4_1 _09464_ (.A(_04293_),
    .B(_04260_),
    .C(net18),
    .D(net19),
    .X(_03705_));
 sky130_fd_sc_hd__inv_2 _09465_ (.A(_03705_),
    .Y(_03706_));
 sky130_fd_sc_hd__a22o_1 _09466_ (.A1(_04293_),
    .A2(net19),
    .B1(_04260_),
    .B2(net18),
    .X(_03707_));
 sky130_fd_sc_hd__nand2_1 _09467_ (.A(_03706_),
    .B(_03707_),
    .Y(_03708_));
 sky130_fd_sc_hd__xnor2_1 _09468_ (.A(_03704_),
    .B(_03708_),
    .Y(_03709_));
 sky130_fd_sc_hd__nand2_1 _09469_ (.A(_03703_),
    .B(_03709_),
    .Y(_03711_));
 sky130_fd_sc_hd__nand3b_2 _09470_ (.A_N(_03709_),
    .B(_03701_),
    .C(_03702_),
    .Y(_03712_));
 sky130_fd_sc_hd__nand2_1 _09471_ (.A(_03711_),
    .B(_03712_),
    .Y(_03713_));
 sky130_fd_sc_hd__nand3_1 _09472_ (.A(_03713_),
    .B(_03486_),
    .C(_03497_),
    .Y(_03714_));
 sky130_fd_sc_hd__nand2_1 _09473_ (.A(_03497_),
    .B(_03486_),
    .Y(_03715_));
 sky130_fd_sc_hd__nand3_2 _09474_ (.A(_03711_),
    .B(_03715_),
    .C(_03712_),
    .Y(_03716_));
 sky130_fd_sc_hd__nand3b_2 _09475_ (.A_N(_03692_),
    .B(_03714_),
    .C(_03716_),
    .Y(_03717_));
 sky130_fd_sc_hd__nand2_1 _09476_ (.A(_03714_),
    .B(_03716_),
    .Y(_03718_));
 sky130_fd_sc_hd__nand2_1 _09477_ (.A(_03718_),
    .B(_03692_),
    .Y(_03719_));
 sky130_fd_sc_hd__nand2_1 _09478_ (.A(_03717_),
    .B(_03719_),
    .Y(_03720_));
 sky130_fd_sc_hd__nand2_1 _09479_ (.A(_03529_),
    .B(_03500_),
    .Y(_03722_));
 sky130_fd_sc_hd__inv_2 _09480_ (.A(_03722_),
    .Y(_03723_));
 sky130_fd_sc_hd__nand2_1 _09481_ (.A(_03720_),
    .B(_03723_),
    .Y(_03724_));
 sky130_fd_sc_hd__nand3_2 _09482_ (.A(_03722_),
    .B(_03717_),
    .C(_03719_),
    .Y(_03725_));
 sky130_fd_sc_hd__nand2_1 _09483_ (.A(_03724_),
    .B(_03725_),
    .Y(_03726_));
 sky130_fd_sc_hd__nand2_1 _09484_ (.A(_03544_),
    .B(_03540_),
    .Y(_03727_));
 sky130_fd_sc_hd__and4_1 _09485_ (.A(_01323_),
    .B(_00784_),
    .C(_05032_),
    .D(_05029_),
    .X(_03728_));
 sky130_fd_sc_hd__inv_2 _09486_ (.A(_03728_),
    .Y(_03729_));
 sky130_fd_sc_hd__a22o_1 _09487_ (.A1(_01323_),
    .A2(_05032_),
    .B1(_00784_),
    .B2(_05029_),
    .X(_03730_));
 sky130_fd_sc_hd__nand2_1 _09488_ (.A(_03729_),
    .B(_03730_),
    .Y(_03731_));
 sky130_fd_sc_hd__nand2_1 _09489_ (.A(_03215_),
    .B(_00740_),
    .Y(_03733_));
 sky130_fd_sc_hd__inv_2 _09490_ (.A(_03733_),
    .Y(_03734_));
 sky130_fd_sc_hd__or2b_1 _09491_ (.A(_03731_),
    .B_N(_03734_),
    .X(_03735_));
 sky130_fd_sc_hd__nand2_1 _09492_ (.A(_03731_),
    .B(_03733_),
    .Y(_03736_));
 sky130_fd_sc_hd__nand2_1 _09493_ (.A(_03735_),
    .B(_03736_),
    .Y(_03737_));
 sky130_fd_sc_hd__or2_1 _09494_ (.A(_03727_),
    .B(_03737_),
    .X(_03738_));
 sky130_fd_sc_hd__nand2_1 _09495_ (.A(_03737_),
    .B(_03727_),
    .Y(_03739_));
 sky130_fd_sc_hd__nand2_1 _09496_ (.A(_03809_),
    .B(_01037_),
    .Y(_03740_));
 sky130_fd_sc_hd__and4_1 _09497_ (.A(_04964_),
    .B(_04962_),
    .C(_00850_),
    .D(_01081_),
    .X(_03741_));
 sky130_fd_sc_hd__inv_2 _09498_ (.A(_03741_),
    .Y(_03742_));
 sky130_fd_sc_hd__a22o_1 _09499_ (.A1(_04964_),
    .A2(_00850_),
    .B1(_04962_),
    .B2(_01081_),
    .X(_03744_));
 sky130_fd_sc_hd__nand2_1 _09500_ (.A(_03742_),
    .B(_03744_),
    .Y(_03745_));
 sky130_fd_sc_hd__xnor2_1 _09501_ (.A(_03740_),
    .B(_03745_),
    .Y(_03746_));
 sky130_fd_sc_hd__a21o_1 _09502_ (.A1(_03738_),
    .A2(_03739_),
    .B1(_03746_),
    .X(_03747_));
 sky130_fd_sc_hd__nand3_1 _09503_ (.A(_03738_),
    .B(_03746_),
    .C(_03739_),
    .Y(_03748_));
 sky130_fd_sc_hd__nand2_1 _09504_ (.A(_03747_),
    .B(_03748_),
    .Y(_03749_));
 sky130_fd_sc_hd__nand2_1 _09505_ (.A(_03510_),
    .B(_03517_),
    .Y(_03750_));
 sky130_fd_sc_hd__inv_2 _09506_ (.A(_03522_),
    .Y(_03751_));
 sky130_fd_sc_hd__nor2_1 _09507_ (.A(_03517_),
    .B(_03510_),
    .Y(_03752_));
 sky130_fd_sc_hd__a21oi_2 _09508_ (.A1(_03750_),
    .A2(_03751_),
    .B1(_03752_),
    .Y(_03753_));
 sky130_fd_sc_hd__inv_2 _09509_ (.A(_03753_),
    .Y(_03755_));
 sky130_fd_sc_hd__nand2_1 _09510_ (.A(_03749_),
    .B(_03755_),
    .Y(_03756_));
 sky130_fd_sc_hd__nand3_1 _09511_ (.A(_03747_),
    .B(_03748_),
    .C(_03753_),
    .Y(_03757_));
 sky130_fd_sc_hd__nand2_1 _09512_ (.A(_03756_),
    .B(_03757_),
    .Y(_03758_));
 sky130_fd_sc_hd__a21o_1 _09513_ (.A1(_03548_),
    .A2(_03557_),
    .B1(_03547_),
    .X(_03759_));
 sky130_fd_sc_hd__nand2_1 _09514_ (.A(_03758_),
    .B(_03759_),
    .Y(_03760_));
 sky130_fd_sc_hd__nand3b_1 _09515_ (.A_N(_03759_),
    .B(_03756_),
    .C(_03757_),
    .Y(_03761_));
 sky130_fd_sc_hd__nand2_1 _09516_ (.A(_03760_),
    .B(_03761_),
    .Y(_03762_));
 sky130_fd_sc_hd__nand2_1 _09517_ (.A(_03726_),
    .B(_03762_),
    .Y(_03763_));
 sky130_fd_sc_hd__nand3b_2 _09518_ (.A_N(_03762_),
    .B(_03724_),
    .C(_03725_),
    .Y(_03764_));
 sky130_fd_sc_hd__nand2_1 _09519_ (.A(_03763_),
    .B(_03764_),
    .Y(_03766_));
 sky130_fd_sc_hd__nand2_1 _09520_ (.A(_03572_),
    .B(_03533_),
    .Y(_03767_));
 sky130_fd_sc_hd__inv_2 _09521_ (.A(_03767_),
    .Y(_03768_));
 sky130_fd_sc_hd__nand2_1 _09522_ (.A(_03766_),
    .B(_03768_),
    .Y(_03769_));
 sky130_fd_sc_hd__nand3_2 _09523_ (.A(_03767_),
    .B(_03763_),
    .C(_03764_),
    .Y(_03770_));
 sky130_fd_sc_hd__nand2_1 _09524_ (.A(_03769_),
    .B(_03770_),
    .Y(_03771_));
 sky130_fd_sc_hd__inv_2 _09525_ (.A(_03440_),
    .Y(_03772_));
 sky130_fd_sc_hd__nor2_1 _09526_ (.A(_03437_),
    .B(_03772_),
    .Y(_03773_));
 sky130_fd_sc_hd__a31o_1 _09527_ (.A1(_03552_),
    .A2(_03809_),
    .A3(_01147_),
    .B1(_03551_),
    .X(_03774_));
 sky130_fd_sc_hd__and4_1 _09528_ (.A(_04812_),
    .B(_04808_),
    .C(_01147_),
    .D(_02544_),
    .X(_03775_));
 sky130_fd_sc_hd__inv_2 _09529_ (.A(_03775_),
    .Y(_03777_));
 sky130_fd_sc_hd__a22o_1 _09530_ (.A1(_04812_),
    .A2(_01147_),
    .B1(_04808_),
    .B2(_02544_),
    .X(_03778_));
 sky130_fd_sc_hd__nand2_1 _09531_ (.A(_03777_),
    .B(_03778_),
    .Y(_03779_));
 sky130_fd_sc_hd__inv_2 _09532_ (.A(_03779_),
    .Y(_03780_));
 sky130_fd_sc_hd__nand2_1 _09533_ (.A(_04818_),
    .B(_01873_),
    .Y(_03781_));
 sky130_fd_sc_hd__inv_2 _09534_ (.A(_03781_),
    .Y(_03782_));
 sky130_fd_sc_hd__nand2_1 _09535_ (.A(_03780_),
    .B(_03782_),
    .Y(_03783_));
 sky130_fd_sc_hd__nand2_1 _09536_ (.A(_03779_),
    .B(_03781_),
    .Y(_03784_));
 sky130_fd_sc_hd__nand2_1 _09537_ (.A(_03783_),
    .B(_03784_),
    .Y(_03785_));
 sky130_fd_sc_hd__or2_1 _09538_ (.A(_03774_),
    .B(_03785_),
    .X(_03786_));
 sky130_fd_sc_hd__nand2_1 _09539_ (.A(_03785_),
    .B(_03774_),
    .Y(_03788_));
 sky130_fd_sc_hd__nand2_1 _09540_ (.A(_03786_),
    .B(_03788_),
    .Y(_03789_));
 sky130_fd_sc_hd__xor2_1 _09541_ (.A(_03773_),
    .B(_03789_),
    .X(_03790_));
 sky130_fd_sc_hd__nand2_1 _09542_ (.A(_03454_),
    .B(_03449_),
    .Y(_03791_));
 sky130_fd_sc_hd__inv_2 _09543_ (.A(_03791_),
    .Y(_03792_));
 sky130_fd_sc_hd__nand2b_1 _09544_ (.A_N(_03790_),
    .B(_03792_),
    .Y(_03793_));
 sky130_fd_sc_hd__nand2_1 _09545_ (.A(_03790_),
    .B(_03791_),
    .Y(_03794_));
 sky130_fd_sc_hd__nand2_1 _09546_ (.A(_03793_),
    .B(_03794_),
    .Y(_03795_));
 sky130_fd_sc_hd__nand2_1 _09547_ (.A(_04876_),
    .B(_03182_),
    .Y(_03796_));
 sky130_fd_sc_hd__inv_2 _09548_ (.A(_04871_),
    .Y(_03797_));
 sky130_fd_sc_hd__or4b_1 _09549_ (.A(_00110_),
    .B(_03797_),
    .C(_02952_),
    .D_N(_03160_),
    .X(_03799_));
 sky130_fd_sc_hd__a22o_1 _09550_ (.A1(_04873_),
    .A2(_02049_),
    .B1(_04871_),
    .B2(_03160_),
    .X(_03800_));
 sky130_fd_sc_hd__nand2_1 _09551_ (.A(_03799_),
    .B(_03800_),
    .Y(_03801_));
 sky130_fd_sc_hd__or2_1 _09552_ (.A(_03796_),
    .B(_03801_),
    .X(_03802_));
 sky130_fd_sc_hd__nand2_1 _09553_ (.A(_03801_),
    .B(_03796_),
    .Y(_03803_));
 sky130_fd_sc_hd__nand2_1 _09554_ (.A(_03802_),
    .B(_03803_),
    .Y(_03804_));
 sky130_fd_sc_hd__nand2_1 _09555_ (.A(_03418_),
    .B(_03415_),
    .Y(_03805_));
 sky130_fd_sc_hd__nand2_1 _09556_ (.A(_03804_),
    .B(_03805_),
    .Y(_03806_));
 sky130_fd_sc_hd__inv_2 _09557_ (.A(_03805_),
    .Y(_03807_));
 sky130_fd_sc_hd__nand3_1 _09558_ (.A(_03802_),
    .B(_03807_),
    .C(_03803_),
    .Y(_03808_));
 sky130_fd_sc_hd__nand2_1 _09559_ (.A(_03806_),
    .B(_03808_),
    .Y(_03810_));
 sky130_fd_sc_hd__nand2_1 _09560_ (.A(_00529_),
    .B(_04928_),
    .Y(_03811_));
 sky130_fd_sc_hd__inv_2 _09561_ (.A(_03811_),
    .Y(_03812_));
 sky130_fd_sc_hd__and4_1 _09562_ (.A(net46),
    .B(_00124_),
    .C(_05031_),
    .D(_05028_),
    .X(_03813_));
 sky130_fd_sc_hd__a22o_1 _09563_ (.A1(net46),
    .A2(_05031_),
    .B1(_00124_),
    .B2(_05028_),
    .X(_03814_));
 sky130_fd_sc_hd__or2b_1 _09564_ (.A(_03813_),
    .B_N(_03814_),
    .X(_03815_));
 sky130_fd_sc_hd__xor2_1 _09565_ (.A(_03812_),
    .B(_03815_),
    .X(_03816_));
 sky130_fd_sc_hd__inv_2 _09566_ (.A(_03816_),
    .Y(_03817_));
 sky130_fd_sc_hd__nand2_1 _09567_ (.A(_03810_),
    .B(_03817_),
    .Y(_03818_));
 sky130_fd_sc_hd__nand3_1 _09568_ (.A(_03806_),
    .B(_03816_),
    .C(_03808_),
    .Y(_03819_));
 sky130_fd_sc_hd__nand2_1 _09569_ (.A(_03818_),
    .B(_03819_),
    .Y(_03821_));
 sky130_fd_sc_hd__inv_2 _09570_ (.A(_03821_),
    .Y(_03822_));
 sky130_fd_sc_hd__nand2_1 _09571_ (.A(_03795_),
    .B(_03822_),
    .Y(_03823_));
 sky130_fd_sc_hd__nand3_1 _09572_ (.A(_03793_),
    .B(_03821_),
    .C(_03794_),
    .Y(_03824_));
 sky130_fd_sc_hd__nand2_1 _09573_ (.A(_03823_),
    .B(_03824_),
    .Y(_03825_));
 sky130_fd_sc_hd__nand2_1 _09574_ (.A(_03559_),
    .B(_03562_),
    .Y(_03826_));
 sky130_fd_sc_hd__nor2_1 _09575_ (.A(_03562_),
    .B(_03559_),
    .Y(_03827_));
 sky130_fd_sc_hd__a21oi_2 _09576_ (.A1(_03826_),
    .A2(_03565_),
    .B1(_03827_),
    .Y(_03828_));
 sky130_fd_sc_hd__inv_2 _09577_ (.A(_03828_),
    .Y(_03829_));
 sky130_fd_sc_hd__nand2_1 _09578_ (.A(_03825_),
    .B(_03829_),
    .Y(_03830_));
 sky130_fd_sc_hd__nand3_1 _09579_ (.A(_03823_),
    .B(_03824_),
    .C(_03828_),
    .Y(_03832_));
 sky130_fd_sc_hd__nand2_1 _09580_ (.A(_03830_),
    .B(_03832_),
    .Y(_03833_));
 sky130_fd_sc_hd__nand2_1 _09581_ (.A(_03459_),
    .B(_03456_),
    .Y(_03834_));
 sky130_fd_sc_hd__nand2_1 _09582_ (.A(_03833_),
    .B(_03834_),
    .Y(_03835_));
 sky130_fd_sc_hd__nand3b_1 _09583_ (.A_N(_03834_),
    .B(_03830_),
    .C(_03832_),
    .Y(_03836_));
 sky130_fd_sc_hd__nand2_1 _09584_ (.A(_03835_),
    .B(_03836_),
    .Y(_03837_));
 sky130_fd_sc_hd__nand2_1 _09585_ (.A(_03771_),
    .B(_03837_),
    .Y(_03838_));
 sky130_fd_sc_hd__inv_2 _09586_ (.A(_03837_),
    .Y(_03839_));
 sky130_fd_sc_hd__nand3_2 _09587_ (.A(_03839_),
    .B(_03769_),
    .C(_03770_),
    .Y(_03840_));
 sky130_fd_sc_hd__nand3_2 _09588_ (.A(_03671_),
    .B(_03838_),
    .C(_03840_),
    .Y(_03841_));
 sky130_fd_sc_hd__nand2_1 _09589_ (.A(_03838_),
    .B(_03840_),
    .Y(_03843_));
 sky130_fd_sc_hd__a21boi_1 _09590_ (.A1(_03474_),
    .A2(_03575_),
    .B1_N(_03576_),
    .Y(_03844_));
 sky130_fd_sc_hd__nand2_1 _09591_ (.A(_03843_),
    .B(_03844_),
    .Y(_03845_));
 sky130_fd_sc_hd__nand2_1 _09592_ (.A(_03841_),
    .B(_03845_),
    .Y(_03846_));
 sky130_fd_sc_hd__and2_1 _09593_ (.A(_03420_),
    .B(_03411_),
    .X(_03847_));
 sky130_fd_sc_hd__nor2_1 _09594_ (.A(_03411_),
    .B(_03420_),
    .Y(_03848_));
 sky130_fd_sc_hd__o21ba_1 _09595_ (.A1(_03429_),
    .A2(_03847_),
    .B1_N(_03848_),
    .X(_03849_));
 sky130_fd_sc_hd__a31o_1 _09596_ (.A1(_03427_),
    .A2(_00529_),
    .A3(_00656_),
    .B1(_03426_),
    .X(_03850_));
 sky130_fd_sc_hd__and4_1 _09597_ (.A(net49),
    .B(net50),
    .C(_00656_),
    .D(_00254_),
    .X(_03851_));
 sky130_fd_sc_hd__inv_2 _09598_ (.A(_03851_),
    .Y(_03852_));
 sky130_fd_sc_hd__a22o_1 _09599_ (.A1(net49),
    .A2(_00656_),
    .B1(net50),
    .B2(_00254_),
    .X(_03854_));
 sky130_fd_sc_hd__nand2_1 _09600_ (.A(_03852_),
    .B(_03854_),
    .Y(_03855_));
 sky130_fd_sc_hd__nand2_1 _09601_ (.A(net51),
    .B(_00522_),
    .Y(_03856_));
 sky130_fd_sc_hd__inv_2 _09602_ (.A(_03856_),
    .Y(_03857_));
 sky130_fd_sc_hd__or2b_1 _09603_ (.A(_03855_),
    .B_N(_03857_),
    .X(_03858_));
 sky130_fd_sc_hd__nand2_1 _09604_ (.A(_03855_),
    .B(_03856_),
    .Y(_03859_));
 sky130_fd_sc_hd__nand2_1 _09605_ (.A(_03858_),
    .B(_03859_),
    .Y(_03860_));
 sky130_fd_sc_hd__or2_1 _09606_ (.A(_03850_),
    .B(_03860_),
    .X(_03861_));
 sky130_fd_sc_hd__nand2_1 _09607_ (.A(_03860_),
    .B(_03850_),
    .Y(_03862_));
 sky130_fd_sc_hd__nand2_1 _09608_ (.A(_03599_),
    .B(_03593_),
    .Y(_03863_));
 sky130_fd_sc_hd__inv_2 _09609_ (.A(_03863_),
    .Y(_03865_));
 sky130_fd_sc_hd__a21o_1 _09610_ (.A1(_03861_),
    .A2(_03862_),
    .B1(_03865_),
    .X(_03866_));
 sky130_fd_sc_hd__nand3_1 _09611_ (.A(_03861_),
    .B(_03865_),
    .C(_03862_),
    .Y(_03867_));
 sky130_fd_sc_hd__nand2_1 _09612_ (.A(_03866_),
    .B(_03867_),
    .Y(_03868_));
 sky130_fd_sc_hd__nor2_1 _09613_ (.A(_03849_),
    .B(_03868_),
    .Y(_03869_));
 sky130_fd_sc_hd__o21ai_2 _09614_ (.A1(_03602_),
    .A2(_03590_),
    .B1(_03606_),
    .Y(_03870_));
 sky130_fd_sc_hd__nand2_1 _09615_ (.A(_03868_),
    .B(_03849_),
    .Y(_03871_));
 sky130_fd_sc_hd__nand3b_1 _09616_ (.A_N(_03869_),
    .B(_03870_),
    .C(_03871_),
    .Y(_03872_));
 sky130_fd_sc_hd__or2b_1 _09617_ (.A(_03868_),
    .B_N(_03849_),
    .X(_03873_));
 sky130_fd_sc_hd__a21o_1 _09618_ (.A1(_03866_),
    .A2(_03867_),
    .B1(_03849_),
    .X(_03874_));
 sky130_fd_sc_hd__nand3b_1 _09619_ (.A_N(_03870_),
    .B(_03873_),
    .C(_03874_),
    .Y(_03876_));
 sky130_fd_sc_hd__nand2_1 _09620_ (.A(_03872_),
    .B(_03876_),
    .Y(_03877_));
 sky130_fd_sc_hd__nand2_1 _09621_ (.A(_03608_),
    .B(_03610_),
    .Y(_03878_));
 sky130_fd_sc_hd__nor2_1 _09622_ (.A(_03610_),
    .B(_03608_),
    .Y(_03879_));
 sky130_fd_sc_hd__a21oi_2 _09623_ (.A1(_03878_),
    .A2(_03614_),
    .B1(_03879_),
    .Y(_03880_));
 sky130_fd_sc_hd__inv_2 _09624_ (.A(_03880_),
    .Y(_03881_));
 sky130_fd_sc_hd__nand2_1 _09625_ (.A(_03877_),
    .B(_03881_),
    .Y(_03882_));
 sky130_fd_sc_hd__nand3_1 _09626_ (.A(_03872_),
    .B(_03876_),
    .C(_03880_),
    .Y(_03883_));
 sky130_fd_sc_hd__nand2_1 _09627_ (.A(_03882_),
    .B(_03883_),
    .Y(_03884_));
 sky130_fd_sc_hd__nand2_1 _09628_ (.A(net54),
    .B(_04992_),
    .Y(_03885_));
 sky130_fd_sc_hd__and4_1 _09629_ (.A(net52),
    .B(net53),
    .C(_04828_),
    .D(_04991_),
    .X(_03887_));
 sky130_fd_sc_hd__a22o_1 _09630_ (.A1(net52),
    .A2(_04828_),
    .B1(net53),
    .B2(_04991_),
    .X(_03888_));
 sky130_fd_sc_hd__and2b_1 _09631_ (.A_N(_03887_),
    .B(_03888_),
    .X(_03889_));
 sky130_fd_sc_hd__xor2_1 _09632_ (.A(_03885_),
    .B(_03889_),
    .X(_03890_));
 sky130_fd_sc_hd__or2_1 _09633_ (.A(_03626_),
    .B(_03890_),
    .X(_03891_));
 sky130_fd_sc_hd__nand2_1 _09634_ (.A(_03890_),
    .B(_03626_),
    .Y(_03892_));
 sky130_fd_sc_hd__nand2_1 _09635_ (.A(_03891_),
    .B(_03892_),
    .Y(_03893_));
 sky130_fd_sc_hd__inv_2 _09636_ (.A(_03893_),
    .Y(_03894_));
 sky130_fd_sc_hd__nand2_1 _09637_ (.A(_03884_),
    .B(_03894_),
    .Y(_03895_));
 sky130_fd_sc_hd__nand3_1 _09638_ (.A(_03882_),
    .B(_03883_),
    .C(_03893_),
    .Y(_03896_));
 sky130_fd_sc_hd__nand2_1 _09639_ (.A(_03895_),
    .B(_03896_),
    .Y(_03898_));
 sky130_fd_sc_hd__nand2_1 _09640_ (.A(_03463_),
    .B(_03464_),
    .Y(_03899_));
 sky130_fd_sc_hd__nor2_1 _09641_ (.A(_03464_),
    .B(_03463_),
    .Y(_03900_));
 sky130_fd_sc_hd__a21oi_2 _09642_ (.A1(_03899_),
    .A2(_03470_),
    .B1(_03900_),
    .Y(_03901_));
 sky130_fd_sc_hd__inv_2 _09643_ (.A(_03901_),
    .Y(_03902_));
 sky130_fd_sc_hd__nand2_1 _09644_ (.A(_03898_),
    .B(_03902_),
    .Y(_03903_));
 sky130_fd_sc_hd__nand3_1 _09645_ (.A(_03895_),
    .B(_03901_),
    .C(_03896_),
    .Y(_03904_));
 sky130_fd_sc_hd__nand2_1 _09646_ (.A(_03903_),
    .B(_03904_),
    .Y(_03905_));
 sky130_fd_sc_hd__nor2_1 _09647_ (.A(_03620_),
    .B(_03617_),
    .Y(_03906_));
 sky130_fd_sc_hd__inv_2 _09648_ (.A(_03630_),
    .Y(_03907_));
 sky130_fd_sc_hd__nor2_1 _09649_ (.A(_03906_),
    .B(_03907_),
    .Y(_03909_));
 sky130_fd_sc_hd__inv_2 _09650_ (.A(_03909_),
    .Y(_03910_));
 sky130_fd_sc_hd__nand2_1 _09651_ (.A(_03905_),
    .B(_03910_),
    .Y(_03911_));
 sky130_fd_sc_hd__nand3_1 _09652_ (.A(_03903_),
    .B(_03904_),
    .C(_03909_),
    .Y(_03912_));
 sky130_fd_sc_hd__nand2_1 _09653_ (.A(_03911_),
    .B(_03912_),
    .Y(_03913_));
 sky130_fd_sc_hd__nand2_1 _09654_ (.A(_03846_),
    .B(_03913_),
    .Y(_03914_));
 sky130_fd_sc_hd__inv_2 _09655_ (.A(_03913_),
    .Y(_03915_));
 sky130_fd_sc_hd__nand3_2 _09656_ (.A(_03915_),
    .B(_03841_),
    .C(_03845_),
    .Y(_03916_));
 sky130_fd_sc_hd__nand2_1 _09657_ (.A(_03914_),
    .B(_03916_),
    .Y(_03917_));
 sky130_fd_sc_hd__nand2_1 _09658_ (.A(_03648_),
    .B(_03584_),
    .Y(_03918_));
 sky130_fd_sc_hd__inv_2 _09659_ (.A(_03918_),
    .Y(_03920_));
 sky130_fd_sc_hd__nand2_1 _09660_ (.A(_03917_),
    .B(_03920_),
    .Y(_03921_));
 sky130_fd_sc_hd__nand3_1 _09661_ (.A(_03918_),
    .B(_03914_),
    .C(_03916_),
    .Y(_03922_));
 sky130_fd_sc_hd__nand2_1 _09662_ (.A(_03921_),
    .B(_03922_),
    .Y(_03923_));
 sky130_fd_sc_hd__nor2_1 _09663_ (.A(_03636_),
    .B(_03632_),
    .Y(_03924_));
 sky130_fd_sc_hd__inv_2 _09664_ (.A(_03642_),
    .Y(_03925_));
 sky130_fd_sc_hd__nor2_1 _09665_ (.A(_03924_),
    .B(_03925_),
    .Y(_03926_));
 sky130_fd_sc_hd__nand2_1 _09666_ (.A(_03923_),
    .B(_03926_),
    .Y(_03927_));
 sky130_fd_sc_hd__nand3b_2 _09667_ (.A_N(_03926_),
    .B(_03921_),
    .C(_03922_),
    .Y(_03928_));
 sky130_fd_sc_hd__nand2_1 _09668_ (.A(_03927_),
    .B(_03928_),
    .Y(_03929_));
 sky130_fd_sc_hd__nand2_1 _09669_ (.A(_03658_),
    .B(_03652_),
    .Y(_03931_));
 sky130_fd_sc_hd__inv_2 _09670_ (.A(_03931_),
    .Y(_03932_));
 sky130_fd_sc_hd__nand2_1 _09671_ (.A(_03929_),
    .B(_03932_),
    .Y(_03933_));
 sky130_fd_sc_hd__nand3_2 _09672_ (.A(_03931_),
    .B(_03927_),
    .C(_03928_),
    .Y(_03934_));
 sky130_fd_sc_hd__nand2_1 _09673_ (.A(_03933_),
    .B(_03934_),
    .Y(_03935_));
 sky130_fd_sc_hd__nand2_1 _09674_ (.A(_03935_),
    .B(_03664_),
    .Y(_03936_));
 sky130_fd_sc_hd__nand3b_1 _09675_ (.A_N(_03664_),
    .B(_03933_),
    .C(_03934_),
    .Y(_03937_));
 sky130_fd_sc_hd__nand2_1 _09676_ (.A(_03936_),
    .B(_03937_),
    .Y(_03938_));
 sky130_fd_sc_hd__nor2_1 _09677_ (.A(_03670_),
    .B(_03938_),
    .Y(_03939_));
 sky130_fd_sc_hd__nand2_1 _09678_ (.A(_03410_),
    .B(_03939_),
    .Y(_03940_));
 sky130_fd_sc_hd__inv_2 _09679_ (.A(_03669_),
    .Y(_03942_));
 sky130_fd_sc_hd__a21boi_1 _09680_ (.A1(_03936_),
    .A2(_03942_),
    .B1_N(_03937_),
    .Y(_03943_));
 sky130_fd_sc_hd__nand2_1 _09681_ (.A(_03940_),
    .B(_03943_),
    .Y(_03944_));
 sky130_fd_sc_hd__and2_1 _09682_ (.A(_03928_),
    .B(_03922_),
    .X(_03945_));
 sky130_fd_sc_hd__and2_1 _09683_ (.A(_03916_),
    .B(_03841_),
    .X(_03946_));
 sky130_fd_sc_hd__nand2_1 _09684_ (.A(_04818_),
    .B(_02544_),
    .Y(_03947_));
 sky130_fd_sc_hd__inv_2 _09685_ (.A(_04808_),
    .Y(_03948_));
 sky130_fd_sc_hd__or4_1 _09686_ (.A(_00263_),
    .B(_03948_),
    .C(_03443_),
    .D(_02913_),
    .X(_03949_));
 sky130_fd_sc_hd__a22o_1 _09687_ (.A1(_04812_),
    .A2(_01037_),
    .B1(_04808_),
    .B2(_01147_),
    .X(_03950_));
 sky130_fd_sc_hd__nand2_1 _09688_ (.A(_03949_),
    .B(_03950_),
    .Y(_03951_));
 sky130_fd_sc_hd__or2_1 _09689_ (.A(_03947_),
    .B(_03951_),
    .X(_03953_));
 sky130_fd_sc_hd__nand2_1 _09690_ (.A(_03951_),
    .B(_03947_),
    .Y(_03954_));
 sky130_fd_sc_hd__nand2_1 _09691_ (.A(_03953_),
    .B(_03954_),
    .Y(_03955_));
 sky130_fd_sc_hd__inv_2 _09692_ (.A(_03744_),
    .Y(_03956_));
 sky130_fd_sc_hd__o21a_1 _09693_ (.A1(_03740_),
    .A2(_03956_),
    .B1(_03742_),
    .X(_03957_));
 sky130_fd_sc_hd__inv_2 _09694_ (.A(_03957_),
    .Y(_03958_));
 sky130_fd_sc_hd__nand2_1 _09695_ (.A(_03955_),
    .B(_03958_),
    .Y(_03959_));
 sky130_fd_sc_hd__nand3_1 _09696_ (.A(_03953_),
    .B(_03957_),
    .C(_03954_),
    .Y(_03960_));
 sky130_fd_sc_hd__nand2_1 _09697_ (.A(_03959_),
    .B(_03960_),
    .Y(_03961_));
 sky130_fd_sc_hd__nand2_1 _09698_ (.A(_03783_),
    .B(_03777_),
    .Y(_03962_));
 sky130_fd_sc_hd__nand2_1 _09699_ (.A(_03961_),
    .B(_03962_),
    .Y(_03964_));
 sky130_fd_sc_hd__nand3b_1 _09700_ (.A_N(_03962_),
    .B(_03959_),
    .C(_03960_),
    .Y(_03965_));
 sky130_fd_sc_hd__nand2_1 _09701_ (.A(_03964_),
    .B(_03965_),
    .Y(_03966_));
 sky130_fd_sc_hd__inv_2 _09702_ (.A(_03774_),
    .Y(_03967_));
 sky130_fd_sc_hd__nor2_1 _09703_ (.A(_03785_),
    .B(_03967_),
    .Y(_03968_));
 sky130_fd_sc_hd__a21oi_1 _09704_ (.A1(_03786_),
    .A2(_03788_),
    .B1(_03773_),
    .Y(_03969_));
 sky130_fd_sc_hd__nor2_1 _09705_ (.A(_03968_),
    .B(_03969_),
    .Y(_03970_));
 sky130_fd_sc_hd__nand2b_1 _09706_ (.A_N(_03966_),
    .B(_03970_),
    .Y(_03971_));
 sky130_fd_sc_hd__o21ai_1 _09707_ (.A1(_03968_),
    .A2(_03969_),
    .B1(_03966_),
    .Y(_03972_));
 sky130_fd_sc_hd__nand2_1 _09708_ (.A(_03971_),
    .B(_03972_),
    .Y(_03973_));
 sky130_fd_sc_hd__nand2_1 _09709_ (.A(_04876_),
    .B(_03160_),
    .Y(_03975_));
 sky130_fd_sc_hd__or4_1 _09710_ (.A(_00110_),
    .B(_03797_),
    .C(_02410_),
    .D(_02952_),
    .X(_03976_));
 sky130_fd_sc_hd__a22o_1 _09711_ (.A1(_04873_),
    .A2(_01873_),
    .B1(_04871_),
    .B2(_02049_),
    .X(_03977_));
 sky130_fd_sc_hd__nand2_1 _09712_ (.A(_03976_),
    .B(_03977_),
    .Y(_03978_));
 sky130_fd_sc_hd__or2_1 _09713_ (.A(_03975_),
    .B(_03978_),
    .X(_03979_));
 sky130_fd_sc_hd__nand2_1 _09714_ (.A(_03978_),
    .B(_03975_),
    .Y(_03980_));
 sky130_fd_sc_hd__nand2_1 _09715_ (.A(_03979_),
    .B(_03980_),
    .Y(_03981_));
 sky130_fd_sc_hd__nand2_1 _09716_ (.A(_03802_),
    .B(_03799_),
    .Y(_03982_));
 sky130_fd_sc_hd__inv_2 _09717_ (.A(_03982_),
    .Y(_03983_));
 sky130_fd_sc_hd__nor2_1 _09718_ (.A(_03981_),
    .B(_03983_),
    .Y(_03984_));
 sky130_fd_sc_hd__and2_1 _09719_ (.A(_03983_),
    .B(_03981_),
    .X(_03986_));
 sky130_fd_sc_hd__nand2_1 _09720_ (.A(_00529_),
    .B(_05028_),
    .Y(_03987_));
 sky130_fd_sc_hd__inv_2 _09721_ (.A(_03987_),
    .Y(_03988_));
 sky130_fd_sc_hd__and4_1 _09722_ (.A(net46),
    .B(_00124_),
    .C(_03182_),
    .D(_05031_),
    .X(_03989_));
 sky130_fd_sc_hd__a22o_1 _09723_ (.A1(net46),
    .A2(_03182_),
    .B1(_00124_),
    .B2(_05031_),
    .X(_03990_));
 sky130_fd_sc_hd__or2b_1 _09724_ (.A(_03989_),
    .B_N(_03990_),
    .X(_03991_));
 sky130_fd_sc_hd__xor2_1 _09725_ (.A(_03988_),
    .B(_03991_),
    .X(_03992_));
 sky130_fd_sc_hd__o21ai_1 _09726_ (.A1(_03984_),
    .A2(_03986_),
    .B1(_03992_),
    .Y(_03993_));
 sky130_fd_sc_hd__inv_2 _09727_ (.A(_03992_),
    .Y(_03994_));
 sky130_fd_sc_hd__nand2_1 _09728_ (.A(_03983_),
    .B(_03981_),
    .Y(_03995_));
 sky130_fd_sc_hd__nand3b_1 _09729_ (.A_N(_03984_),
    .B(_03994_),
    .C(_03995_),
    .Y(_03997_));
 sky130_fd_sc_hd__nand2_1 _09730_ (.A(_03993_),
    .B(_03997_),
    .Y(_03998_));
 sky130_fd_sc_hd__inv_2 _09731_ (.A(_03998_),
    .Y(_03999_));
 sky130_fd_sc_hd__nand2_1 _09732_ (.A(_03973_),
    .B(_03999_),
    .Y(_04000_));
 sky130_fd_sc_hd__nand3_1 _09733_ (.A(_03971_),
    .B(_03998_),
    .C(_03972_),
    .Y(_04001_));
 sky130_fd_sc_hd__nand2_1 _09734_ (.A(_04000_),
    .B(_04001_),
    .Y(_04002_));
 sky130_fd_sc_hd__o21a_1 _09735_ (.A1(_03749_),
    .A2(_03753_),
    .B1(_03760_),
    .X(_04003_));
 sky130_fd_sc_hd__inv_2 _09736_ (.A(_04003_),
    .Y(_04004_));
 sky130_fd_sc_hd__nand2_1 _09737_ (.A(_04002_),
    .B(_04004_),
    .Y(_04005_));
 sky130_fd_sc_hd__nand3_1 _09738_ (.A(_04000_),
    .B(_04001_),
    .C(_04003_),
    .Y(_04006_));
 sky130_fd_sc_hd__nand2_1 _09739_ (.A(_04005_),
    .B(_04006_),
    .Y(_04008_));
 sky130_fd_sc_hd__nor2_1 _09740_ (.A(_03792_),
    .B(_03790_),
    .Y(_04009_));
 sky130_fd_sc_hd__inv_2 _09741_ (.A(_03823_),
    .Y(_04010_));
 sky130_fd_sc_hd__nor2_1 _09742_ (.A(_04009_),
    .B(_04010_),
    .Y(_04011_));
 sky130_fd_sc_hd__inv_2 _09743_ (.A(_04011_),
    .Y(_04012_));
 sky130_fd_sc_hd__nand2_1 _09744_ (.A(_04008_),
    .B(_04012_),
    .Y(_04013_));
 sky130_fd_sc_hd__nand3_1 _09745_ (.A(_04005_),
    .B(_04006_),
    .C(_04011_),
    .Y(_04014_));
 sky130_fd_sc_hd__nand2_1 _09746_ (.A(_04013_),
    .B(_04014_),
    .Y(_04015_));
 sky130_fd_sc_hd__inv_2 _09747_ (.A(_04015_),
    .Y(_04016_));
 sky130_fd_sc_hd__nand2_1 _09748_ (.A(_01535_),
    .B(net21),
    .Y(_04017_));
 sky130_fd_sc_hd__inv_2 _09749_ (.A(net24),
    .Y(_04019_));
 sky130_fd_sc_hd__nand2_1 _09750_ (.A(_02357_),
    .B(net22),
    .Y(_04020_));
 sky130_fd_sc_hd__nor3_1 _09751_ (.A(_01597_),
    .B(_04019_),
    .C(_04020_),
    .Y(_04021_));
 sky130_fd_sc_hd__o21ai_1 _09752_ (.A1(_01597_),
    .A2(_04019_),
    .B1(_04020_),
    .Y(_04022_));
 sky130_fd_sc_hd__and2b_1 _09753_ (.A_N(_04021_),
    .B(_04022_),
    .X(_04023_));
 sky130_fd_sc_hd__xor2_1 _09754_ (.A(_04017_),
    .B(_04023_),
    .X(_04024_));
 sky130_fd_sc_hd__a31o_1 _09755_ (.A1(_03695_),
    .A2(_01535_),
    .A3(net20),
    .B1(_03694_),
    .X(_04025_));
 sky130_fd_sc_hd__inv_2 _09756_ (.A(_04025_),
    .Y(_04026_));
 sky130_fd_sc_hd__nor2_1 _09757_ (.A(_04024_),
    .B(_04026_),
    .Y(_04027_));
 sky130_fd_sc_hd__inv_2 _09758_ (.A(_04027_),
    .Y(_04028_));
 sky130_fd_sc_hd__nand2_1 _09759_ (.A(_04026_),
    .B(_04024_),
    .Y(_04030_));
 sky130_fd_sc_hd__nand2_1 _09760_ (.A(_01565_),
    .B(net18),
    .Y(_04031_));
 sky130_fd_sc_hd__nand2_1 _09761_ (.A(_04260_),
    .B(net19),
    .Y(_04032_));
 sky130_fd_sc_hd__nor3_1 _09762_ (.A(_02086_),
    .B(_03087_),
    .C(_04032_),
    .Y(_04033_));
 sky130_fd_sc_hd__o21ai_1 _09763_ (.A1(_02086_),
    .A2(_03087_),
    .B1(_04032_),
    .Y(_04034_));
 sky130_fd_sc_hd__and2b_1 _09764_ (.A_N(_04033_),
    .B(_04034_),
    .X(_04035_));
 sky130_fd_sc_hd__xor2_1 _09765_ (.A(_04031_),
    .B(_04035_),
    .X(_04036_));
 sky130_fd_sc_hd__inv_2 _09766_ (.A(_04036_),
    .Y(_04037_));
 sky130_fd_sc_hd__a21o_1 _09767_ (.A1(_04028_),
    .A2(_04030_),
    .B1(_04037_),
    .X(_04038_));
 sky130_fd_sc_hd__nand3_1 _09768_ (.A(_04028_),
    .B(_04037_),
    .C(_04030_),
    .Y(_04039_));
 sky130_fd_sc_hd__nand2_1 _09769_ (.A(_04038_),
    .B(_04039_),
    .Y(_04041_));
 sky130_fd_sc_hd__and2_1 _09770_ (.A(_03712_),
    .B(_03702_),
    .X(_04042_));
 sky130_fd_sc_hd__nor2_1 _09771_ (.A(_04041_),
    .B(_04042_),
    .Y(_04043_));
 sky130_fd_sc_hd__inv_2 _09772_ (.A(_04043_),
    .Y(_04044_));
 sky130_fd_sc_hd__nand2_1 _09773_ (.A(_04042_),
    .B(_04041_),
    .Y(_04045_));
 sky130_fd_sc_hd__nand2_1 _09774_ (.A(_04044_),
    .B(_04045_),
    .Y(_04046_));
 sky130_fd_sc_hd__nand2_1 _09775_ (.A(_00003_),
    .B(_05160_),
    .Y(_04047_));
 sky130_fd_sc_hd__nand2_1 _09776_ (.A(_00412_),
    .B(_00393_),
    .Y(_04048_));
 sky130_fd_sc_hd__nor3_1 _09777_ (.A(_01937_),
    .B(_03511_),
    .C(_04048_),
    .Y(_04049_));
 sky130_fd_sc_hd__inv_2 _09778_ (.A(_04049_),
    .Y(_04050_));
 sky130_fd_sc_hd__o21ai_1 _09779_ (.A1(_01937_),
    .A2(_03511_),
    .B1(_04048_),
    .Y(_04052_));
 sky130_fd_sc_hd__nand2_1 _09780_ (.A(_04050_),
    .B(_04052_),
    .Y(_04053_));
 sky130_fd_sc_hd__or2_1 _09781_ (.A(_04047_),
    .B(_04053_),
    .X(_04054_));
 sky130_fd_sc_hd__nand2_1 _09782_ (.A(_04053_),
    .B(_04047_),
    .Y(_04055_));
 sky130_fd_sc_hd__nand2_1 _09783_ (.A(_04054_),
    .B(_04055_),
    .Y(_04056_));
 sky130_fd_sc_hd__inv_2 _09784_ (.A(_03707_),
    .Y(_04057_));
 sky130_fd_sc_hd__o21a_1 _09785_ (.A1(_03704_),
    .A2(_04057_),
    .B1(_03706_),
    .X(_04058_));
 sky130_fd_sc_hd__inv_2 _09786_ (.A(_04058_),
    .Y(_04059_));
 sky130_fd_sc_hd__or2_1 _09787_ (.A(_04056_),
    .B(_04059_),
    .X(_04060_));
 sky130_fd_sc_hd__nand2_1 _09788_ (.A(_04059_),
    .B(_04056_),
    .Y(_04061_));
 sky130_fd_sc_hd__nand2_1 _09789_ (.A(_03681_),
    .B(_03678_),
    .Y(_04063_));
 sky130_fd_sc_hd__inv_2 _09790_ (.A(_04063_),
    .Y(_04064_));
 sky130_fd_sc_hd__a21o_1 _09791_ (.A1(_04060_),
    .A2(_04061_),
    .B1(_04064_),
    .X(_04065_));
 sky130_fd_sc_hd__nand3_1 _09792_ (.A(_04060_),
    .B(_04064_),
    .C(_04061_),
    .Y(_04066_));
 sky130_fd_sc_hd__nand2_1 _09793_ (.A(_04065_),
    .B(_04066_),
    .Y(_04067_));
 sky130_fd_sc_hd__nand2_1 _09794_ (.A(_04046_),
    .B(_04067_),
    .Y(_04068_));
 sky130_fd_sc_hd__inv_2 _09795_ (.A(_04067_),
    .Y(_04069_));
 sky130_fd_sc_hd__nand3_1 _09796_ (.A(_04044_),
    .B(_04069_),
    .C(_04045_),
    .Y(_04070_));
 sky130_fd_sc_hd__nand2_1 _09797_ (.A(_04068_),
    .B(_04070_),
    .Y(_04071_));
 sky130_fd_sc_hd__nand3_2 _09798_ (.A(_04071_),
    .B(_03716_),
    .C(_03717_),
    .Y(_04072_));
 sky130_fd_sc_hd__nand2_1 _09799_ (.A(_03717_),
    .B(_03716_),
    .Y(_04074_));
 sky130_fd_sc_hd__nand3_2 _09800_ (.A(_04074_),
    .B(_04068_),
    .C(_04070_),
    .Y(_04075_));
 sky130_fd_sc_hd__nand2_1 _09801_ (.A(_04072_),
    .B(_04075_),
    .Y(_04076_));
 sky130_fd_sc_hd__nor2_1 _09802_ (.A(_03673_),
    .B(_03683_),
    .Y(_04077_));
 sky130_fd_sc_hd__nand2_1 _09803_ (.A(_03215_),
    .B(_00784_),
    .Y(_04078_));
 sky130_fd_sc_hd__inv_2 _09804_ (.A(_05029_),
    .Y(_04079_));
 sky130_fd_sc_hd__or4_1 _09805_ (.A(_02870_),
    .B(_01957_),
    .C(_04079_),
    .D(_03519_),
    .X(_04080_));
 sky130_fd_sc_hd__a22o_1 _09806_ (.A1(_01323_),
    .A2(_05029_),
    .B1(_05032_),
    .B2(_04084_),
    .X(_04081_));
 sky130_fd_sc_hd__nand2_1 _09807_ (.A(_04080_),
    .B(_04081_),
    .Y(_04082_));
 sky130_fd_sc_hd__or2_1 _09808_ (.A(_04078_),
    .B(_04082_),
    .X(_04083_));
 sky130_fd_sc_hd__nand2_1 _09809_ (.A(_04082_),
    .B(_04078_),
    .Y(_04085_));
 sky130_fd_sc_hd__nand2_1 _09810_ (.A(_04083_),
    .B(_04085_),
    .Y(_04086_));
 sky130_fd_sc_hd__nand2_1 _09811_ (.A(_03735_),
    .B(_03729_),
    .Y(_04087_));
 sky130_fd_sc_hd__inv_2 _09812_ (.A(_04087_),
    .Y(_04088_));
 sky130_fd_sc_hd__nand2_1 _09813_ (.A(_04086_),
    .B(_04088_),
    .Y(_04089_));
 sky130_fd_sc_hd__nand3_1 _09814_ (.A(_04083_),
    .B(_04087_),
    .C(_04085_),
    .Y(_04090_));
 sky130_fd_sc_hd__nand2_1 _09815_ (.A(_04089_),
    .B(_04090_),
    .Y(_04091_));
 sky130_fd_sc_hd__nand2_1 _09816_ (.A(_03809_),
    .B(_01081_),
    .Y(_04092_));
 sky130_fd_sc_hd__and4_1 _09817_ (.A(_04964_),
    .B(_04962_),
    .C(_00740_),
    .D(_00850_),
    .X(_04093_));
 sky130_fd_sc_hd__a22o_1 _09818_ (.A1(_04964_),
    .A2(_00740_),
    .B1(_04962_),
    .B2(_00850_),
    .X(_04094_));
 sky130_fd_sc_hd__and2b_1 _09819_ (.A_N(_04093_),
    .B(_04094_),
    .X(_04096_));
 sky130_fd_sc_hd__xor2_1 _09820_ (.A(_04092_),
    .B(_04096_),
    .X(_04097_));
 sky130_fd_sc_hd__nand2_1 _09821_ (.A(_04091_),
    .B(_04097_),
    .Y(_04098_));
 sky130_fd_sc_hd__nand3b_1 _09822_ (.A_N(_04097_),
    .B(_04089_),
    .C(_04090_),
    .Y(_04099_));
 sky130_fd_sc_hd__nand2_1 _09823_ (.A(_04098_),
    .B(_04099_),
    .Y(_04100_));
 sky130_fd_sc_hd__o21ai_1 _09824_ (.A1(_04077_),
    .A2(_03689_),
    .B1(_04100_),
    .Y(_04101_));
 sky130_fd_sc_hd__nor2_1 _09825_ (.A(_04077_),
    .B(_03689_),
    .Y(_04102_));
 sky130_fd_sc_hd__nand3_1 _09826_ (.A(_04098_),
    .B(_04099_),
    .C(_04102_),
    .Y(_04103_));
 sky130_fd_sc_hd__nand2_1 _09827_ (.A(_04101_),
    .B(_04103_),
    .Y(_04104_));
 sky130_fd_sc_hd__or2b_1 _09828_ (.A(_03737_),
    .B_N(_03727_),
    .X(_04105_));
 sky130_fd_sc_hd__nand2_1 _09829_ (.A(_03747_),
    .B(_04105_),
    .Y(_04107_));
 sky130_fd_sc_hd__nand2_1 _09830_ (.A(_04104_),
    .B(_04107_),
    .Y(_04108_));
 sky130_fd_sc_hd__nand3b_1 _09831_ (.A_N(_04107_),
    .B(_04101_),
    .C(_04103_),
    .Y(_04109_));
 sky130_fd_sc_hd__nand2_1 _09832_ (.A(_04108_),
    .B(_04109_),
    .Y(_04110_));
 sky130_fd_sc_hd__nand2_1 _09833_ (.A(_04076_),
    .B(_04110_),
    .Y(_04111_));
 sky130_fd_sc_hd__inv_2 _09834_ (.A(_04110_),
    .Y(_04112_));
 sky130_fd_sc_hd__nand3_2 _09835_ (.A(_04112_),
    .B(_04072_),
    .C(_04075_),
    .Y(_04113_));
 sky130_fd_sc_hd__nand2_1 _09836_ (.A(_04111_),
    .B(_04113_),
    .Y(_04114_));
 sky130_fd_sc_hd__nand2_1 _09837_ (.A(_03764_),
    .B(_03725_),
    .Y(_04115_));
 sky130_fd_sc_hd__inv_2 _09838_ (.A(_04115_),
    .Y(_04116_));
 sky130_fd_sc_hd__nand2_1 _09839_ (.A(_04114_),
    .B(_04116_),
    .Y(_04118_));
 sky130_fd_sc_hd__nand3_2 _09840_ (.A(_04111_),
    .B(_04113_),
    .C(_04115_),
    .Y(_04119_));
 sky130_fd_sc_hd__nand3_1 _09841_ (.A(_04016_),
    .B(_04118_),
    .C(_04119_),
    .Y(_04120_));
 sky130_fd_sc_hd__nand2_1 _09842_ (.A(_04118_),
    .B(_04119_),
    .Y(_04121_));
 sky130_fd_sc_hd__nand2_1 _09843_ (.A(_04121_),
    .B(_04015_),
    .Y(_04122_));
 sky130_fd_sc_hd__nand2_1 _09844_ (.A(_04120_),
    .B(_04122_),
    .Y(_04123_));
 sky130_fd_sc_hd__nand2_1 _09845_ (.A(_03840_),
    .B(_03770_),
    .Y(_04124_));
 sky130_fd_sc_hd__inv_2 _09846_ (.A(_04124_),
    .Y(_04125_));
 sky130_fd_sc_hd__nand2_1 _09847_ (.A(_04123_),
    .B(_04125_),
    .Y(_04126_));
 sky130_fd_sc_hd__nand3_1 _09848_ (.A(_04120_),
    .B(_04122_),
    .C(_04124_),
    .Y(_04127_));
 sky130_fd_sc_hd__nand2_1 _09849_ (.A(_04126_),
    .B(_04127_),
    .Y(_04129_));
 sky130_fd_sc_hd__nand2_1 _09850_ (.A(_03804_),
    .B(_03807_),
    .Y(_04130_));
 sky130_fd_sc_hd__nor2_1 _09851_ (.A(_03807_),
    .B(_03804_),
    .Y(_04131_));
 sky130_fd_sc_hd__a21oi_2 _09852_ (.A1(_04130_),
    .A2(_03817_),
    .B1(_04131_),
    .Y(_04132_));
 sky130_fd_sc_hd__nand2_1 _09853_ (.A(_03858_),
    .B(_03852_),
    .Y(_04133_));
 sky130_fd_sc_hd__nand2_1 _09854_ (.A(net51),
    .B(_00254_),
    .Y(_04134_));
 sky130_fd_sc_hd__inv_2 _09855_ (.A(net50),
    .Y(_04135_));
 sky130_fd_sc_hd__or4_1 _09856_ (.A(_03042_),
    .B(_04135_),
    .C(_02451_),
    .D(_03284_),
    .X(_04136_));
 sky130_fd_sc_hd__a22o_1 _09857_ (.A1(net49),
    .A2(_04928_),
    .B1(net50),
    .B2(_00656_),
    .X(_04137_));
 sky130_fd_sc_hd__nand2_1 _09858_ (.A(_04136_),
    .B(_04137_),
    .Y(_04138_));
 sky130_fd_sc_hd__or2_1 _09859_ (.A(_04134_),
    .B(_04138_),
    .X(_04140_));
 sky130_fd_sc_hd__nand2_1 _09860_ (.A(_04138_),
    .B(_04134_),
    .Y(_04141_));
 sky130_fd_sc_hd__nand2_1 _09861_ (.A(_04140_),
    .B(_04141_),
    .Y(_04142_));
 sky130_fd_sc_hd__a21oi_2 _09862_ (.A1(_03814_),
    .A2(_03812_),
    .B1(_03813_),
    .Y(_04143_));
 sky130_fd_sc_hd__inv_2 _09863_ (.A(_04143_),
    .Y(_04144_));
 sky130_fd_sc_hd__nand2_1 _09864_ (.A(_04142_),
    .B(_04144_),
    .Y(_04145_));
 sky130_fd_sc_hd__nand3_1 _09865_ (.A(_04140_),
    .B(_04143_),
    .C(_04141_),
    .Y(_04146_));
 sky130_fd_sc_hd__nand3b_1 _09866_ (.A_N(_04133_),
    .B(_04145_),
    .C(_04146_),
    .Y(_04147_));
 sky130_fd_sc_hd__nand2_1 _09867_ (.A(_04142_),
    .B(_04143_),
    .Y(_04148_));
 sky130_fd_sc_hd__nand3_1 _09868_ (.A(_04140_),
    .B(_04141_),
    .C(_04144_),
    .Y(_04149_));
 sky130_fd_sc_hd__nand3_1 _09869_ (.A(_04148_),
    .B(_04133_),
    .C(_04149_),
    .Y(_04151_));
 sky130_fd_sc_hd__nand2_1 _09870_ (.A(_04147_),
    .B(_04151_),
    .Y(_04152_));
 sky130_fd_sc_hd__nor2_1 _09871_ (.A(_04132_),
    .B(_04152_),
    .Y(_04153_));
 sky130_fd_sc_hd__inv_2 _09872_ (.A(_04153_),
    .Y(_04154_));
 sky130_fd_sc_hd__and3_1 _09873_ (.A(_03850_),
    .B(_03859_),
    .C(_03858_),
    .X(_04155_));
 sky130_fd_sc_hd__or2b_1 _09874_ (.A(_04155_),
    .B_N(_03866_),
    .X(_04156_));
 sky130_fd_sc_hd__nand2_1 _09875_ (.A(_04152_),
    .B(_04132_),
    .Y(_04157_));
 sky130_fd_sc_hd__nand3_1 _09876_ (.A(_04154_),
    .B(_04156_),
    .C(_04157_),
    .Y(_04158_));
 sky130_fd_sc_hd__nand3_1 _09877_ (.A(_04132_),
    .B(_04151_),
    .C(_04147_),
    .Y(_04159_));
 sky130_fd_sc_hd__inv_2 _09878_ (.A(_04132_),
    .Y(_04160_));
 sky130_fd_sc_hd__nand2_1 _09879_ (.A(_04160_),
    .B(_04152_),
    .Y(_04162_));
 sky130_fd_sc_hd__nand3b_1 _09880_ (.A_N(_04156_),
    .B(_04159_),
    .C(_04162_),
    .Y(_04163_));
 sky130_fd_sc_hd__nand2_1 _09881_ (.A(_04158_),
    .B(_04163_),
    .Y(_04164_));
 sky130_fd_sc_hd__a21oi_2 _09882_ (.A1(_03871_),
    .A2(_03870_),
    .B1(_03869_),
    .Y(_04165_));
 sky130_fd_sc_hd__inv_2 _09883_ (.A(_04165_),
    .Y(_04166_));
 sky130_fd_sc_hd__nand2_1 _09884_ (.A(_04164_),
    .B(_04166_),
    .Y(_04167_));
 sky130_fd_sc_hd__nand3_1 _09885_ (.A(_04158_),
    .B(_04163_),
    .C(_04165_),
    .Y(_04168_));
 sky130_fd_sc_hd__nand2_1 _09886_ (.A(_04167_),
    .B(_04168_),
    .Y(_04169_));
 sky130_fd_sc_hd__nand2_1 _09887_ (.A(net56),
    .B(_04992_),
    .Y(_04170_));
 sky130_fd_sc_hd__a31o_1 _09888_ (.A1(_03888_),
    .A2(net54),
    .A3(_04992_),
    .B1(_03887_),
    .X(_04171_));
 sky130_fd_sc_hd__nand2_1 _09889_ (.A(net54),
    .B(_04991_),
    .Y(_04173_));
 sky130_fd_sc_hd__or4_1 _09890_ (.A(_03624_),
    .B(_03625_),
    .C(_02464_),
    .D(_02085_),
    .X(_04174_));
 sky130_fd_sc_hd__a22o_1 _09891_ (.A1(net52),
    .A2(_00522_),
    .B1(net53),
    .B2(_04828_),
    .X(_04175_));
 sky130_fd_sc_hd__nand2_1 _09892_ (.A(_04174_),
    .B(_04175_),
    .Y(_04176_));
 sky130_fd_sc_hd__or2_1 _09893_ (.A(_04173_),
    .B(_04176_),
    .X(_04177_));
 sky130_fd_sc_hd__nand2_1 _09894_ (.A(_04176_),
    .B(_04173_),
    .Y(_04178_));
 sky130_fd_sc_hd__nand2_1 _09895_ (.A(_04177_),
    .B(_04178_),
    .Y(_04179_));
 sky130_fd_sc_hd__inv_2 _09896_ (.A(_04179_),
    .Y(_04180_));
 sky130_fd_sc_hd__nor2_1 _09897_ (.A(_04171_),
    .B(_04180_),
    .Y(_04181_));
 sky130_fd_sc_hd__nand2_1 _09898_ (.A(_04180_),
    .B(_04171_),
    .Y(_04182_));
 sky130_fd_sc_hd__nand2b_1 _09899_ (.A_N(_04181_),
    .B(_04182_),
    .Y(_04184_));
 sky130_fd_sc_hd__or2_1 _09900_ (.A(_04170_),
    .B(_04184_),
    .X(_04185_));
 sky130_fd_sc_hd__nand2_1 _09901_ (.A(_04184_),
    .B(_04170_),
    .Y(_04186_));
 sky130_fd_sc_hd__nand2_1 _09902_ (.A(_04185_),
    .B(_04186_),
    .Y(_04187_));
 sky130_fd_sc_hd__nand2_1 _09903_ (.A(_04187_),
    .B(_03891_),
    .Y(_04188_));
 sky130_fd_sc_hd__nand3b_2 _09904_ (.A_N(_03891_),
    .B(_04185_),
    .C(_04186_),
    .Y(_04189_));
 sky130_fd_sc_hd__nand2_1 _09905_ (.A(_04188_),
    .B(_04189_),
    .Y(_04190_));
 sky130_fd_sc_hd__inv_2 _09906_ (.A(_04190_),
    .Y(_04191_));
 sky130_fd_sc_hd__nand2_1 _09907_ (.A(_04169_),
    .B(_04191_),
    .Y(_04192_));
 sky130_fd_sc_hd__nand3_1 _09908_ (.A(_04167_),
    .B(_04190_),
    .C(_04168_),
    .Y(_04193_));
 sky130_fd_sc_hd__nand2_1 _09909_ (.A(_04192_),
    .B(_04193_),
    .Y(_04195_));
 sky130_fd_sc_hd__or2_1 _09910_ (.A(_03828_),
    .B(_03825_),
    .X(_04196_));
 sky130_fd_sc_hd__nand2_1 _09911_ (.A(_03835_),
    .B(_04196_),
    .Y(_04197_));
 sky130_fd_sc_hd__nand2_1 _09912_ (.A(_04195_),
    .B(_04197_),
    .Y(_04198_));
 sky130_fd_sc_hd__inv_2 _09913_ (.A(_04197_),
    .Y(_04199_));
 sky130_fd_sc_hd__nand3_1 _09914_ (.A(_04199_),
    .B(_04192_),
    .C(_04193_),
    .Y(_04200_));
 sky130_fd_sc_hd__nand2_1 _09915_ (.A(_04198_),
    .B(_04200_),
    .Y(_04201_));
 sky130_fd_sc_hd__nor2_1 _09916_ (.A(_03880_),
    .B(_03877_),
    .Y(_04202_));
 sky130_fd_sc_hd__inv_2 _09917_ (.A(_03895_),
    .Y(_04203_));
 sky130_fd_sc_hd__nor2_1 _09918_ (.A(_04202_),
    .B(_04203_),
    .Y(_04204_));
 sky130_fd_sc_hd__inv_2 _09919_ (.A(_04204_),
    .Y(_04206_));
 sky130_fd_sc_hd__nand2_1 _09920_ (.A(_04201_),
    .B(_04206_),
    .Y(_04207_));
 sky130_fd_sc_hd__nand3_1 _09921_ (.A(_04198_),
    .B(_04200_),
    .C(_04204_),
    .Y(_04208_));
 sky130_fd_sc_hd__nand2_1 _09922_ (.A(_04207_),
    .B(_04208_),
    .Y(_04209_));
 sky130_fd_sc_hd__nand2_1 _09923_ (.A(_04129_),
    .B(_04209_),
    .Y(_04210_));
 sky130_fd_sc_hd__inv_2 _09924_ (.A(_04209_),
    .Y(_04211_));
 sky130_fd_sc_hd__nand3_1 _09925_ (.A(_04126_),
    .B(_04211_),
    .C(_04127_),
    .Y(_04212_));
 sky130_fd_sc_hd__nand2_1 _09926_ (.A(_04210_),
    .B(_04212_),
    .Y(_04213_));
 sky130_fd_sc_hd__nor2_1 _09927_ (.A(_03946_),
    .B(_04213_),
    .Y(_04214_));
 sky130_fd_sc_hd__inv_2 _09928_ (.A(_04214_),
    .Y(_04215_));
 sky130_fd_sc_hd__nand2_1 _09929_ (.A(_04213_),
    .B(_03946_),
    .Y(_04217_));
 sky130_fd_sc_hd__nand2_1 _09930_ (.A(_04215_),
    .B(_04217_),
    .Y(_04218_));
 sky130_fd_sc_hd__nor2_1 _09931_ (.A(_03901_),
    .B(_03898_),
    .Y(_04219_));
 sky130_fd_sc_hd__inv_2 _09932_ (.A(_03911_),
    .Y(_04220_));
 sky130_fd_sc_hd__nor2_1 _09933_ (.A(_04219_),
    .B(_04220_),
    .Y(_04221_));
 sky130_fd_sc_hd__nand2_1 _09934_ (.A(_04218_),
    .B(_04221_),
    .Y(_04222_));
 sky130_fd_sc_hd__inv_2 _09935_ (.A(_04221_),
    .Y(_04223_));
 sky130_fd_sc_hd__nand3_2 _09936_ (.A(_04215_),
    .B(_04223_),
    .C(_04217_),
    .Y(_04224_));
 sky130_fd_sc_hd__nand3b_4 _09937_ (.A_N(_03945_),
    .B(_04222_),
    .C(_04224_),
    .Y(_04225_));
 sky130_fd_sc_hd__nand2_1 _09938_ (.A(_04222_),
    .B(_04224_),
    .Y(_04226_));
 sky130_fd_sc_hd__nand2_1 _09939_ (.A(_04226_),
    .B(_03945_),
    .Y(_04228_));
 sky130_fd_sc_hd__nand2_1 _09940_ (.A(_04225_),
    .B(_04228_),
    .Y(_04229_));
 sky130_fd_sc_hd__nand2_1 _09941_ (.A(_04229_),
    .B(_03934_),
    .Y(_04230_));
 sky130_fd_sc_hd__nand3b_1 _09942_ (.A_N(_03934_),
    .B(_04225_),
    .C(_04228_),
    .Y(_04231_));
 sky130_fd_sc_hd__nand2_1 _09943_ (.A(_04230_),
    .B(_04231_),
    .Y(_04232_));
 sky130_fd_sc_hd__inv_2 _09944_ (.A(_04232_),
    .Y(_04233_));
 sky130_fd_sc_hd__nand2_1 _09945_ (.A(_03944_),
    .B(_04233_),
    .Y(_04234_));
 sky130_fd_sc_hd__nand2_1 _09946_ (.A(_04234_),
    .B(_04231_),
    .Y(_04235_));
 sky130_fd_sc_hd__a21boi_1 _09947_ (.A1(_04016_),
    .A2(_04118_),
    .B1_N(_04119_),
    .Y(_04236_));
 sky130_fd_sc_hd__a21boi_1 _09948_ (.A1(_04112_),
    .A2(_04072_),
    .B1_N(_04075_),
    .Y(_04237_));
 sky130_fd_sc_hd__nor2_1 _09949_ (.A(_04058_),
    .B(_04056_),
    .Y(_04239_));
 sky130_fd_sc_hd__a21oi_1 _09950_ (.A1(_04060_),
    .A2(_04061_),
    .B1(_04064_),
    .Y(_04240_));
 sky130_fd_sc_hd__nand2_1 _09951_ (.A(_03215_),
    .B(_01323_),
    .Y(_04241_));
 sky130_fd_sc_hd__inv_2 _09952_ (.A(_04241_),
    .Y(_04242_));
 sky130_fd_sc_hd__or4b_1 _09953_ (.A(_01957_),
    .B(_04079_),
    .C(_03519_),
    .D_N(_05160_),
    .X(_04243_));
 sky130_fd_sc_hd__a22o_1 _09954_ (.A1(_05032_),
    .A2(_05160_),
    .B1(_05029_),
    .B2(_04084_),
    .X(_04244_));
 sky130_fd_sc_hd__nand2_1 _09955_ (.A(_04243_),
    .B(_04244_),
    .Y(_04245_));
 sky130_fd_sc_hd__xor2_1 _09956_ (.A(_04242_),
    .B(_04245_),
    .X(_04246_));
 sky130_fd_sc_hd__nand2_1 _09957_ (.A(_04083_),
    .B(_04080_),
    .Y(_04247_));
 sky130_fd_sc_hd__nor2_1 _09958_ (.A(_04246_),
    .B(_04247_),
    .Y(_04248_));
 sky130_fd_sc_hd__and2_1 _09959_ (.A(_04247_),
    .B(_04246_),
    .X(_04250_));
 sky130_fd_sc_hd__nand2_1 _09960_ (.A(_03809_),
    .B(_00850_),
    .Y(_04251_));
 sky130_fd_sc_hd__inv_2 _09961_ (.A(_04251_),
    .Y(_04252_));
 sky130_fd_sc_hd__nand2_1 _09962_ (.A(_04962_),
    .B(_00740_),
    .Y(_04253_));
 sky130_fd_sc_hd__nand2_1 _09963_ (.A(_04964_),
    .B(_00784_),
    .Y(_04254_));
 sky130_fd_sc_hd__xnor2_1 _09964_ (.A(_04253_),
    .B(_04254_),
    .Y(_04255_));
 sky130_fd_sc_hd__xor2_1 _09965_ (.A(_04252_),
    .B(_04255_),
    .X(_04256_));
 sky130_fd_sc_hd__o21bai_1 _09966_ (.A1(_04248_),
    .A2(_04250_),
    .B1_N(_04256_),
    .Y(_04257_));
 sky130_fd_sc_hd__nand2_1 _09967_ (.A(_04247_),
    .B(_04246_),
    .Y(_04258_));
 sky130_fd_sc_hd__nand3b_1 _09968_ (.A_N(_04248_),
    .B(_04256_),
    .C(_04258_),
    .Y(_04259_));
 sky130_fd_sc_hd__nand2_1 _09969_ (.A(_04257_),
    .B(_04259_),
    .Y(_04261_));
 sky130_fd_sc_hd__o21ai_1 _09970_ (.A1(_04239_),
    .A2(_04240_),
    .B1(_04261_),
    .Y(_04262_));
 sky130_fd_sc_hd__nand2_1 _09971_ (.A(_04056_),
    .B(_04058_),
    .Y(_04263_));
 sky130_fd_sc_hd__a21oi_1 _09972_ (.A1(_04063_),
    .A2(_04263_),
    .B1(_04239_),
    .Y(_04264_));
 sky130_fd_sc_hd__nand3_1 _09973_ (.A(_04257_),
    .B(_04259_),
    .C(_04264_),
    .Y(_04265_));
 sky130_fd_sc_hd__nand2_1 _09974_ (.A(_04262_),
    .B(_04265_),
    .Y(_04266_));
 sky130_fd_sc_hd__nand2_1 _09975_ (.A(_04099_),
    .B(_04090_),
    .Y(_04267_));
 sky130_fd_sc_hd__nand2_1 _09976_ (.A(_04266_),
    .B(_04267_),
    .Y(_04268_));
 sky130_fd_sc_hd__nand3b_1 _09977_ (.A_N(_04267_),
    .B(_04262_),
    .C(_04265_),
    .Y(_04269_));
 sky130_fd_sc_hd__nand2_1 _09978_ (.A(_04268_),
    .B(_04269_),
    .Y(_04270_));
 sky130_fd_sc_hd__inv_2 _09979_ (.A(_04270_),
    .Y(_04272_));
 sky130_fd_sc_hd__nand2_1 _09980_ (.A(_01565_),
    .B(net19),
    .Y(_04273_));
 sky130_fd_sc_hd__and4_1 _09981_ (.A(_04293_),
    .B(_04260_),
    .C(net20),
    .D(net21),
    .X(_04274_));
 sky130_fd_sc_hd__a22o_1 _09982_ (.A1(_04293_),
    .A2(net21),
    .B1(_04260_),
    .B2(net20),
    .X(_04275_));
 sky130_fd_sc_hd__and2b_1 _09983_ (.A_N(_04274_),
    .B(_04275_),
    .X(_04276_));
 sky130_fd_sc_hd__xor2_1 _09984_ (.A(_04273_),
    .B(_04276_),
    .X(_04277_));
 sky130_fd_sc_hd__a31oi_1 _09985_ (.A1(_04022_),
    .A2(_01535_),
    .A3(net21),
    .B1(_04021_),
    .Y(_04278_));
 sky130_fd_sc_hd__nand2_1 _09986_ (.A(_01535_),
    .B(net22),
    .Y(_04279_));
 sky130_fd_sc_hd__nand2_1 _09987_ (.A(_02357_),
    .B(net24),
    .Y(_04280_));
 sky130_fd_sc_hd__nand2_1 _09988_ (.A(_02379_),
    .B(net25),
    .Y(_04281_));
 sky130_fd_sc_hd__xnor2_1 _09989_ (.A(_04280_),
    .B(_04281_),
    .Y(_04283_));
 sky130_fd_sc_hd__xor2_1 _09990_ (.A(_04279_),
    .B(_04283_),
    .X(_04284_));
 sky130_fd_sc_hd__xor2_1 _09991_ (.A(_04278_),
    .B(_04284_),
    .X(_04285_));
 sky130_fd_sc_hd__xor2_1 _09992_ (.A(_04277_),
    .B(_04285_),
    .X(_04286_));
 sky130_fd_sc_hd__nand2_1 _09993_ (.A(_04039_),
    .B(_04028_),
    .Y(_04287_));
 sky130_fd_sc_hd__or2_1 _09994_ (.A(_04286_),
    .B(_04287_),
    .X(_04288_));
 sky130_fd_sc_hd__nand2_1 _09995_ (.A(_04287_),
    .B(_04286_),
    .Y(_04289_));
 sky130_fd_sc_hd__nand2_1 _09996_ (.A(_04054_),
    .B(_04050_),
    .Y(_04290_));
 sky130_fd_sc_hd__inv_2 _09997_ (.A(_04290_),
    .Y(_04291_));
 sky130_fd_sc_hd__nand2_1 _09998_ (.A(_00003_),
    .B(_00393_),
    .Y(_04292_));
 sky130_fd_sc_hd__nand2_1 _09999_ (.A(_00412_),
    .B(net17),
    .Y(_04294_));
 sky130_fd_sc_hd__nand2_1 _10000_ (.A(_00204_),
    .B(net18),
    .Y(_04295_));
 sky130_fd_sc_hd__xnor2_1 _10001_ (.A(_04294_),
    .B(_04295_),
    .Y(_04296_));
 sky130_fd_sc_hd__xnor2_1 _10002_ (.A(_04292_),
    .B(_04296_),
    .Y(_04297_));
 sky130_fd_sc_hd__a31oi_1 _10003_ (.A1(_04034_),
    .A2(_01565_),
    .A3(net18),
    .B1(_04033_),
    .Y(_04298_));
 sky130_fd_sc_hd__inv_2 _10004_ (.A(_04298_),
    .Y(_04299_));
 sky130_fd_sc_hd__or2_1 _10005_ (.A(_04297_),
    .B(_04299_),
    .X(_04300_));
 sky130_fd_sc_hd__nand2_1 _10006_ (.A(_04299_),
    .B(_04297_),
    .Y(_04301_));
 sky130_fd_sc_hd__nand2_1 _10007_ (.A(_04300_),
    .B(_04301_),
    .Y(_04302_));
 sky130_fd_sc_hd__xor2_1 _10008_ (.A(_04291_),
    .B(_04302_),
    .X(_04303_));
 sky130_fd_sc_hd__a21o_1 _10009_ (.A1(_04288_),
    .A2(_04289_),
    .B1(_04303_),
    .X(_04305_));
 sky130_fd_sc_hd__nand3_1 _10010_ (.A(_04288_),
    .B(_04303_),
    .C(_04289_),
    .Y(_04306_));
 sky130_fd_sc_hd__a21oi_1 _10011_ (.A1(_04045_),
    .A2(_04069_),
    .B1(_04043_),
    .Y(_04307_));
 sky130_fd_sc_hd__a21o_1 _10012_ (.A1(_04305_),
    .A2(_04306_),
    .B1(_04307_),
    .X(_04308_));
 sky130_fd_sc_hd__nand3_1 _10013_ (.A(_04305_),
    .B(_04307_),
    .C(_04306_),
    .Y(_04309_));
 sky130_fd_sc_hd__nand2_1 _10014_ (.A(_04308_),
    .B(_04309_),
    .Y(_04310_));
 sky130_fd_sc_hd__nand2_1 _10015_ (.A(_04272_),
    .B(_04310_),
    .Y(_04311_));
 sky130_fd_sc_hd__nand3_1 _10016_ (.A(_04270_),
    .B(_04308_),
    .C(_04309_),
    .Y(_04312_));
 sky130_fd_sc_hd__nand3_1 _10017_ (.A(_04237_),
    .B(_04311_),
    .C(_04312_),
    .Y(_04313_));
 sky130_fd_sc_hd__nand2_1 _10018_ (.A(_04312_),
    .B(_04311_),
    .Y(_04314_));
 sky130_fd_sc_hd__nand2_1 _10019_ (.A(_04113_),
    .B(_04075_),
    .Y(_04316_));
 sky130_fd_sc_hd__nand2_1 _10020_ (.A(_04314_),
    .B(_04316_),
    .Y(_04317_));
 sky130_fd_sc_hd__nand2_1 _10021_ (.A(_04313_),
    .B(_04317_),
    .Y(_04318_));
 sky130_fd_sc_hd__nor2_1 _10022_ (.A(_03957_),
    .B(_03955_),
    .Y(_04319_));
 sky130_fd_sc_hd__and2_1 _10023_ (.A(_03961_),
    .B(_03962_),
    .X(_04320_));
 sky130_fd_sc_hd__a31oi_1 _10024_ (.A1(_04094_),
    .A2(_03809_),
    .A3(_01081_),
    .B1(_04093_),
    .Y(_04321_));
 sky130_fd_sc_hd__inv_2 _10025_ (.A(_04321_),
    .Y(_04322_));
 sky130_fd_sc_hd__nand2_1 _10026_ (.A(_04818_),
    .B(_01147_),
    .Y(_04323_));
 sky130_fd_sc_hd__or4_1 _10027_ (.A(_00263_),
    .B(_02619_),
    .C(_03948_),
    .D(_03443_),
    .X(_04324_));
 sky130_fd_sc_hd__a22o_1 _10028_ (.A1(_04812_),
    .A2(_01081_),
    .B1(_04808_),
    .B2(_01037_),
    .X(_04325_));
 sky130_fd_sc_hd__nand2_1 _10029_ (.A(_04324_),
    .B(_04325_),
    .Y(_04327_));
 sky130_fd_sc_hd__xnor2_1 _10030_ (.A(_04323_),
    .B(_04327_),
    .Y(_04328_));
 sky130_fd_sc_hd__or2_1 _10031_ (.A(_04322_),
    .B(_04328_),
    .X(_04329_));
 sky130_fd_sc_hd__nand2_1 _10032_ (.A(_04328_),
    .B(_04322_),
    .Y(_04330_));
 sky130_fd_sc_hd__nand2_1 _10033_ (.A(_04329_),
    .B(_04330_),
    .Y(_04331_));
 sky130_fd_sc_hd__nand2_1 _10034_ (.A(_03953_),
    .B(_03949_),
    .Y(_04332_));
 sky130_fd_sc_hd__nand2_1 _10035_ (.A(_04331_),
    .B(_04332_),
    .Y(_04333_));
 sky130_fd_sc_hd__nand3b_1 _10036_ (.A_N(_04332_),
    .B(_04329_),
    .C(_04330_),
    .Y(_04334_));
 sky130_fd_sc_hd__nand2_1 _10037_ (.A(_04333_),
    .B(_04334_),
    .Y(_04335_));
 sky130_fd_sc_hd__o21ai_1 _10038_ (.A1(_04319_),
    .A2(_04320_),
    .B1(_04335_),
    .Y(_04336_));
 sky130_fd_sc_hd__nand2_1 _10039_ (.A(_03955_),
    .B(_03957_),
    .Y(_04338_));
 sky130_fd_sc_hd__a21oi_1 _10040_ (.A1(_04338_),
    .A2(_03962_),
    .B1(_04319_),
    .Y(_04339_));
 sky130_fd_sc_hd__nand3_1 _10041_ (.A(_04333_),
    .B(_04334_),
    .C(_04339_),
    .Y(_04340_));
 sky130_fd_sc_hd__nand2_1 _10042_ (.A(_04336_),
    .B(_04340_),
    .Y(_04341_));
 sky130_fd_sc_hd__nand2_1 _10043_ (.A(_04876_),
    .B(_02049_),
    .Y(_04342_));
 sky130_fd_sc_hd__or4_1 _10044_ (.A(_00110_),
    .B(_02961_),
    .C(_03797_),
    .D(_02410_),
    .X(_04343_));
 sky130_fd_sc_hd__a22o_1 _10045_ (.A1(_04873_),
    .A2(_02544_),
    .B1(_04871_),
    .B2(_01873_),
    .X(_04344_));
 sky130_fd_sc_hd__nand2_1 _10046_ (.A(_04343_),
    .B(_04344_),
    .Y(_04345_));
 sky130_fd_sc_hd__xnor2_1 _10047_ (.A(_04342_),
    .B(_04345_),
    .Y(_04346_));
 sky130_fd_sc_hd__nand2_1 _10048_ (.A(_03979_),
    .B(_03976_),
    .Y(_04347_));
 sky130_fd_sc_hd__xnor2_1 _10049_ (.A(_04346_),
    .B(_04347_),
    .Y(_04349_));
 sky130_fd_sc_hd__nand2_1 _10050_ (.A(_00529_),
    .B(_05031_),
    .Y(_04350_));
 sky130_fd_sc_hd__nand2_1 _10051_ (.A(_00124_),
    .B(_03182_),
    .Y(_04351_));
 sky130_fd_sc_hd__nand2_1 _10052_ (.A(_03160_),
    .B(net46),
    .Y(_04352_));
 sky130_fd_sc_hd__xnor2_1 _10053_ (.A(_04351_),
    .B(_04352_),
    .Y(_04353_));
 sky130_fd_sc_hd__xnor2_1 _10054_ (.A(_04350_),
    .B(_04353_),
    .Y(_04354_));
 sky130_fd_sc_hd__or2b_1 _10055_ (.A(_04349_),
    .B_N(_04354_),
    .X(_04355_));
 sky130_fd_sc_hd__or2b_1 _10056_ (.A(_04354_),
    .B_N(_04349_),
    .X(_04356_));
 sky130_fd_sc_hd__nand2_1 _10057_ (.A(_04355_),
    .B(_04356_),
    .Y(_04357_));
 sky130_fd_sc_hd__inv_2 _10058_ (.A(_04357_),
    .Y(_04358_));
 sky130_fd_sc_hd__nand2_1 _10059_ (.A(_04341_),
    .B(_04358_),
    .Y(_04360_));
 sky130_fd_sc_hd__nand3_1 _10060_ (.A(_04336_),
    .B(_04357_),
    .C(_04340_),
    .Y(_04361_));
 sky130_fd_sc_hd__nand2_1 _10061_ (.A(_04360_),
    .B(_04361_),
    .Y(_04362_));
 sky130_fd_sc_hd__nand2_1 _10062_ (.A(_04100_),
    .B(_04102_),
    .Y(_04363_));
 sky130_fd_sc_hd__nor2_1 _10063_ (.A(_04102_),
    .B(_04100_),
    .Y(_04364_));
 sky130_fd_sc_hd__a21oi_1 _10064_ (.A1(_04363_),
    .A2(_04107_),
    .B1(_04364_),
    .Y(_04365_));
 sky130_fd_sc_hd__inv_2 _10065_ (.A(_04365_),
    .Y(_04366_));
 sky130_fd_sc_hd__nand2_1 _10066_ (.A(_04362_),
    .B(_04366_),
    .Y(_04367_));
 sky130_fd_sc_hd__nand3_1 _10067_ (.A(_04360_),
    .B(_04361_),
    .C(_04365_),
    .Y(_04368_));
 sky130_fd_sc_hd__nand2_1 _10068_ (.A(_04367_),
    .B(_04368_),
    .Y(_04369_));
 sky130_fd_sc_hd__o21ai_1 _10069_ (.A1(_03970_),
    .A2(_03966_),
    .B1(_04000_),
    .Y(_04371_));
 sky130_fd_sc_hd__nand2_1 _10070_ (.A(_04369_),
    .B(_04371_),
    .Y(_04372_));
 sky130_fd_sc_hd__nand3b_1 _10071_ (.A_N(_04371_),
    .B(_04367_),
    .C(_04368_),
    .Y(_04373_));
 sky130_fd_sc_hd__nand2_1 _10072_ (.A(_04372_),
    .B(_04373_),
    .Y(_04374_));
 sky130_fd_sc_hd__inv_2 _10073_ (.A(_04374_),
    .Y(_04375_));
 sky130_fd_sc_hd__nand2_1 _10074_ (.A(_04318_),
    .B(_04375_),
    .Y(_04376_));
 sky130_fd_sc_hd__nand3_1 _10075_ (.A(_04374_),
    .B(_04313_),
    .C(_04317_),
    .Y(_04377_));
 sky130_fd_sc_hd__nand3_1 _10076_ (.A(_04236_),
    .B(_04376_),
    .C(_04377_),
    .Y(_04378_));
 sky130_fd_sc_hd__nand2_1 _10077_ (.A(_04376_),
    .B(_04377_),
    .Y(_04379_));
 sky130_fd_sc_hd__nand2_1 _10078_ (.A(_04120_),
    .B(_04119_),
    .Y(_04380_));
 sky130_fd_sc_hd__nand2_1 _10079_ (.A(_04379_),
    .B(_04380_),
    .Y(_04382_));
 sky130_fd_sc_hd__nand2_1 _10080_ (.A(_04378_),
    .B(_04382_),
    .Y(_04383_));
 sky130_fd_sc_hd__a21oi_1 _10081_ (.A1(_03990_),
    .A2(_03988_),
    .B1(_03989_),
    .Y(_04384_));
 sky130_fd_sc_hd__inv_2 _10082_ (.A(_04384_),
    .Y(_04385_));
 sky130_fd_sc_hd__nand2_1 _10083_ (.A(net51),
    .B(_00656_),
    .Y(_04386_));
 sky130_fd_sc_hd__or4_1 _10084_ (.A(_03042_),
    .B(_02699_),
    .C(_04135_),
    .D(_02451_),
    .X(_04387_));
 sky130_fd_sc_hd__a22o_1 _10085_ (.A1(net49),
    .A2(_05028_),
    .B1(net50),
    .B2(_04928_),
    .X(_04388_));
 sky130_fd_sc_hd__nand2_1 _10086_ (.A(_04387_),
    .B(_04388_),
    .Y(_04389_));
 sky130_fd_sc_hd__xnor2_1 _10087_ (.A(_04386_),
    .B(_04389_),
    .Y(_04390_));
 sky130_fd_sc_hd__or2_1 _10088_ (.A(_04385_),
    .B(_04390_),
    .X(_04391_));
 sky130_fd_sc_hd__nand2_1 _10089_ (.A(_04390_),
    .B(_04385_),
    .Y(_04393_));
 sky130_fd_sc_hd__nand2_1 _10090_ (.A(_04391_),
    .B(_04393_),
    .Y(_04394_));
 sky130_fd_sc_hd__nand2_1 _10091_ (.A(_04140_),
    .B(_04136_),
    .Y(_04395_));
 sky130_fd_sc_hd__nand2_1 _10092_ (.A(_04394_),
    .B(_04395_),
    .Y(_04396_));
 sky130_fd_sc_hd__nand3b_1 _10093_ (.A_N(_04395_),
    .B(_04391_),
    .C(_04393_),
    .Y(_04397_));
 sky130_fd_sc_hd__nand2_1 _10094_ (.A(_04396_),
    .B(_04397_),
    .Y(_04398_));
 sky130_fd_sc_hd__a21oi_1 _10095_ (.A1(_03995_),
    .A2(_03994_),
    .B1(_03984_),
    .Y(_04399_));
 sky130_fd_sc_hd__inv_2 _10096_ (.A(_04399_),
    .Y(_04400_));
 sky130_fd_sc_hd__nand2_1 _10097_ (.A(_04398_),
    .B(_04400_),
    .Y(_04401_));
 sky130_fd_sc_hd__nand3_1 _10098_ (.A(_04399_),
    .B(_04396_),
    .C(_04397_),
    .Y(_04402_));
 sky130_fd_sc_hd__nand2_1 _10099_ (.A(_04401_),
    .B(_04402_),
    .Y(_04404_));
 sky130_fd_sc_hd__nand2_1 _10100_ (.A(_04151_),
    .B(_04149_),
    .Y(_04405_));
 sky130_fd_sc_hd__nand2_1 _10101_ (.A(_04404_),
    .B(_04405_),
    .Y(_04406_));
 sky130_fd_sc_hd__nand3b_1 _10102_ (.A_N(_04405_),
    .B(_04401_),
    .C(_04402_),
    .Y(_04407_));
 sky130_fd_sc_hd__nand2_1 _10103_ (.A(_04406_),
    .B(_04407_),
    .Y(_04408_));
 sky130_fd_sc_hd__a21oi_1 _10104_ (.A1(_04157_),
    .A2(_04156_),
    .B1(_04153_),
    .Y(_04409_));
 sky130_fd_sc_hd__inv_2 _10105_ (.A(_04409_),
    .Y(_04410_));
 sky130_fd_sc_hd__nand2_1 _10106_ (.A(_04408_),
    .B(_04410_),
    .Y(_04411_));
 sky130_fd_sc_hd__nand3_1 _10107_ (.A(_04406_),
    .B(_04407_),
    .C(_04409_),
    .Y(_04412_));
 sky130_fd_sc_hd__nand2_1 _10108_ (.A(_04411_),
    .B(_04412_),
    .Y(_04413_));
 sky130_fd_sc_hd__and3_1 _10109_ (.A(_04177_),
    .B(_04171_),
    .C(_04178_),
    .X(_04415_));
 sky130_fd_sc_hd__nor2_1 _10110_ (.A(_04170_),
    .B(_04184_),
    .Y(_04416_));
 sky130_fd_sc_hd__nand2_1 _10111_ (.A(net56),
    .B(_04991_),
    .Y(_04417_));
 sky130_fd_sc_hd__nand2_1 _10112_ (.A(net54),
    .B(_04828_),
    .Y(_04418_));
 sky130_fd_sc_hd__or4_1 _10113_ (.A(_03624_),
    .B(_00111_),
    .C(_03625_),
    .D(_02464_),
    .X(_04419_));
 sky130_fd_sc_hd__a22o_1 _10114_ (.A1(net52),
    .A2(_00254_),
    .B1(net53),
    .B2(_00522_),
    .X(_04420_));
 sky130_fd_sc_hd__nand2_1 _10115_ (.A(_04419_),
    .B(_04420_),
    .Y(_04421_));
 sky130_fd_sc_hd__xnor2_1 _10116_ (.A(_04418_),
    .B(_04421_),
    .Y(_04422_));
 sky130_fd_sc_hd__nand2_1 _10117_ (.A(_04177_),
    .B(_04174_),
    .Y(_04423_));
 sky130_fd_sc_hd__xnor2_1 _10118_ (.A(_04422_),
    .B(_04423_),
    .Y(_04424_));
 sky130_fd_sc_hd__or2_1 _10119_ (.A(_04417_),
    .B(_04424_),
    .X(_04426_));
 sky130_fd_sc_hd__nand2_1 _10120_ (.A(_04424_),
    .B(_04417_),
    .Y(_04427_));
 sky130_fd_sc_hd__nand2_1 _10121_ (.A(_04426_),
    .B(_04427_),
    .Y(_04428_));
 sky130_fd_sc_hd__o21ai_1 _10122_ (.A1(_04415_),
    .A2(_04416_),
    .B1(_04428_),
    .Y(_04429_));
 sky130_fd_sc_hd__o21a_1 _10123_ (.A1(_04170_),
    .A2(_04181_),
    .B1(_04182_),
    .X(_04430_));
 sky130_fd_sc_hd__nand3_1 _10124_ (.A(_04426_),
    .B(_04430_),
    .C(_04427_),
    .Y(_04431_));
 sky130_fd_sc_hd__nand2_1 _10125_ (.A(_04429_),
    .B(_04431_),
    .Y(_04432_));
 sky130_fd_sc_hd__nand2_1 _10126_ (.A(net57),
    .B(_04992_),
    .Y(_04433_));
 sky130_fd_sc_hd__nand2_1 _10127_ (.A(_04432_),
    .B(_04433_),
    .Y(_04434_));
 sky130_fd_sc_hd__nand3b_1 _10128_ (.A_N(_04433_),
    .B(_04429_),
    .C(_04431_),
    .Y(_04435_));
 sky130_fd_sc_hd__nand3_1 _10129_ (.A(_04413_),
    .B(_04434_),
    .C(_04435_),
    .Y(_04437_));
 sky130_fd_sc_hd__nand2_1 _10130_ (.A(_04434_),
    .B(_04435_),
    .Y(_04438_));
 sky130_fd_sc_hd__nand3_1 _10131_ (.A(_04438_),
    .B(_04411_),
    .C(_04412_),
    .Y(_04439_));
 sky130_fd_sc_hd__nand2_1 _10132_ (.A(_04437_),
    .B(_04439_),
    .Y(_04440_));
 sky130_fd_sc_hd__nand2_1 _10133_ (.A(_04002_),
    .B(_04003_),
    .Y(_04441_));
 sky130_fd_sc_hd__nor2_1 _10134_ (.A(_04003_),
    .B(_04002_),
    .Y(_04442_));
 sky130_fd_sc_hd__a21oi_2 _10135_ (.A1(_04441_),
    .A2(_04012_),
    .B1(_04442_),
    .Y(_04443_));
 sky130_fd_sc_hd__inv_2 _10136_ (.A(_04443_),
    .Y(_04444_));
 sky130_fd_sc_hd__nand2_1 _10137_ (.A(_04440_),
    .B(_04444_),
    .Y(_04445_));
 sky130_fd_sc_hd__nand3_1 _10138_ (.A(_04437_),
    .B(_04439_),
    .C(_04443_),
    .Y(_04446_));
 sky130_fd_sc_hd__nand2_1 _10139_ (.A(_04445_),
    .B(_04446_),
    .Y(_04448_));
 sky130_fd_sc_hd__nor2_1 _10140_ (.A(_04165_),
    .B(_04164_),
    .Y(_04449_));
 sky130_fd_sc_hd__inv_2 _10141_ (.A(_04192_),
    .Y(_04450_));
 sky130_fd_sc_hd__nor2_1 _10142_ (.A(_04449_),
    .B(_04450_),
    .Y(_04451_));
 sky130_fd_sc_hd__inv_2 _10143_ (.A(_04451_),
    .Y(_04452_));
 sky130_fd_sc_hd__nand2_1 _10144_ (.A(_04448_),
    .B(_04452_),
    .Y(_04453_));
 sky130_fd_sc_hd__nand3_1 _10145_ (.A(_04445_),
    .B(_04446_),
    .C(_04451_),
    .Y(_04454_));
 sky130_fd_sc_hd__nand2_1 _10146_ (.A(_04453_),
    .B(_04454_),
    .Y(_04455_));
 sky130_fd_sc_hd__inv_2 _10147_ (.A(_04455_),
    .Y(_04456_));
 sky130_fd_sc_hd__nand2_1 _10148_ (.A(_04383_),
    .B(_04456_),
    .Y(_04457_));
 sky130_fd_sc_hd__nand3_1 _10149_ (.A(_04378_),
    .B(_04455_),
    .C(_04382_),
    .Y(_04459_));
 sky130_fd_sc_hd__nand2_1 _10150_ (.A(_04457_),
    .B(_04459_),
    .Y(_04460_));
 sky130_fd_sc_hd__a21boi_1 _10151_ (.A1(_04126_),
    .A2(_04211_),
    .B1_N(_04127_),
    .Y(_04461_));
 sky130_fd_sc_hd__inv_2 _10152_ (.A(_04461_),
    .Y(_04462_));
 sky130_fd_sc_hd__nand2_1 _10153_ (.A(_04460_),
    .B(_04462_),
    .Y(_04463_));
 sky130_fd_sc_hd__nand3_1 _10154_ (.A(_04461_),
    .B(_04457_),
    .C(_04459_),
    .Y(_04464_));
 sky130_fd_sc_hd__nand2_1 _10155_ (.A(_04463_),
    .B(_04464_),
    .Y(_04465_));
 sky130_fd_sc_hd__nor2_1 _10156_ (.A(_04199_),
    .B(_04195_),
    .Y(_04466_));
 sky130_fd_sc_hd__inv_2 _10157_ (.A(_04207_),
    .Y(_04467_));
 sky130_fd_sc_hd__nor2_1 _10158_ (.A(_04466_),
    .B(_04467_),
    .Y(_04468_));
 sky130_fd_sc_hd__inv_2 _10159_ (.A(_04468_),
    .Y(_04470_));
 sky130_fd_sc_hd__nand2_1 _10160_ (.A(_04465_),
    .B(_04470_),
    .Y(_04471_));
 sky130_fd_sc_hd__nand3_1 _10161_ (.A(_04463_),
    .B(_04464_),
    .C(_04468_),
    .Y(_04472_));
 sky130_fd_sc_hd__nand2_1 _10162_ (.A(_04471_),
    .B(_04472_),
    .Y(_04473_));
 sky130_fd_sc_hd__a21oi_1 _10163_ (.A1(_04217_),
    .A2(_04223_),
    .B1(_04214_),
    .Y(_04474_));
 sky130_fd_sc_hd__inv_2 _10164_ (.A(_04474_),
    .Y(_04475_));
 sky130_fd_sc_hd__nand2_1 _10165_ (.A(_04473_),
    .B(_04475_),
    .Y(_04476_));
 sky130_fd_sc_hd__nand3_1 _10166_ (.A(_04471_),
    .B(_04474_),
    .C(_04472_),
    .Y(_04477_));
 sky130_fd_sc_hd__nand2_1 _10167_ (.A(_04476_),
    .B(_04477_),
    .Y(_04478_));
 sky130_fd_sc_hd__nand2_1 _10168_ (.A(_04478_),
    .B(_04189_),
    .Y(_04479_));
 sky130_fd_sc_hd__nand3b_1 _10169_ (.A_N(_04189_),
    .B(_04476_),
    .C(_04477_),
    .Y(_04481_));
 sky130_fd_sc_hd__nand2_1 _10170_ (.A(_04479_),
    .B(_04481_),
    .Y(_04482_));
 sky130_fd_sc_hd__nand2_1 _10171_ (.A(_04482_),
    .B(_04225_),
    .Y(_04483_));
 sky130_fd_sc_hd__nand3b_1 _10172_ (.A_N(_04225_),
    .B(_04479_),
    .C(_04481_),
    .Y(_04484_));
 sky130_fd_sc_hd__nand2_2 _10173_ (.A(_04483_),
    .B(_04484_),
    .Y(_04485_));
 sky130_fd_sc_hd__nand2_1 _10174_ (.A(_04235_),
    .B(_04485_),
    .Y(_04486_));
 sky130_fd_sc_hd__inv_2 _10175_ (.A(_04485_),
    .Y(_04487_));
 sky130_fd_sc_hd__nand3_1 _10176_ (.A(_04234_),
    .B(_04487_),
    .C(_04231_),
    .Y(_04488_));
 sky130_fd_sc_hd__nand2_1 _10177_ (.A(_04486_),
    .B(_04488_),
    .Y(\ab[21] ));
 sky130_fd_sc_hd__nand2_1 _10178_ (.A(net66),
    .B(net144),
    .Y(_04489_));
 sky130_fd_sc_hd__inv_2 _10179_ (.A(net77),
    .Y(_04491_));
 sky130_fd_sc_hd__inv_2 _10180_ (.A(net153),
    .Y(_04492_));
 sky130_fd_sc_hd__nand2_1 _10181_ (.A(_04491_),
    .B(_04492_),
    .Y(_04493_));
 sky130_fd_sc_hd__nand2_1 _10182_ (.A(net186),
    .B(net153),
    .Y(_04494_));
 sky130_fd_sc_hd__nand2_1 _10183_ (.A(net154),
    .B(_04494_),
    .Y(_04495_));
 sky130_fd_sc_hd__or2_1 _10184_ (.A(_04489_),
    .B(net155),
    .X(_04496_));
 sky130_fd_sc_hd__nand2_1 _10185_ (.A(net155),
    .B(_04489_),
    .Y(_04497_));
 sky130_fd_sc_hd__and2_1 _10186_ (.A(_04496_),
    .B(net156),
    .X(_04498_));
 sky130_fd_sc_hd__clkbuf_1 _10187_ (.A(net157),
    .X(\absum[1] ));
 sky130_fd_sc_hd__or2_1 _10188_ (.A(net88),
    .B(net118),
    .X(_04499_));
 sky130_fd_sc_hd__nand2_1 _10189_ (.A(net88),
    .B(net118),
    .Y(_04501_));
 sky130_fd_sc_hd__and2_1 _10190_ (.A(_04499_),
    .B(net119),
    .X(_04502_));
 sky130_fd_sc_hd__nand2_1 _10191_ (.A(_04496_),
    .B(_04494_),
    .Y(_04503_));
 sky130_fd_sc_hd__or2_1 _10192_ (.A(_04502_),
    .B(_04503_),
    .X(_04504_));
 sky130_fd_sc_hd__nand2_1 _10193_ (.A(net187),
    .B(_04502_),
    .Y(_04505_));
 sky130_fd_sc_hd__and2_1 _10194_ (.A(net188),
    .B(_04505_),
    .X(_04506_));
 sky130_fd_sc_hd__clkbuf_1 _10195_ (.A(net189),
    .X(\absum[2] ));
 sky130_fd_sc_hd__nor2_1 _10196_ (.A(net91),
    .B(net195),
    .Y(_04507_));
 sky130_fd_sc_hd__nand2_1 _10197_ (.A(net91),
    .B(net195),
    .Y(_04508_));
 sky130_fd_sc_hd__and2b_1 _10198_ (.A_N(_04507_),
    .B(_04508_),
    .X(_04509_));
 sky130_fd_sc_hd__nand2_1 _10199_ (.A(_04505_),
    .B(net119),
    .Y(_04511_));
 sky130_fd_sc_hd__xor2_1 _10200_ (.A(_04509_),
    .B(net120),
    .X(\absum[3] ));
 sky130_fd_sc_hd__or2_1 _10201_ (.A(net92),
    .B(net176),
    .X(_04512_));
 sky130_fd_sc_hd__nand2_1 _10202_ (.A(net92),
    .B(net176),
    .Y(_04513_));
 sky130_fd_sc_hd__and2_1 _10203_ (.A(_04512_),
    .B(net177),
    .X(_04514_));
 sky130_fd_sc_hd__o21ai_1 _10204_ (.A1(net119),
    .A2(_04507_),
    .B1(net196),
    .Y(_04515_));
 sky130_fd_sc_hd__a31o_1 _10205_ (.A1(_04503_),
    .A2(_04502_),
    .A3(_04509_),
    .B1(net197),
    .X(_04516_));
 sky130_fd_sc_hd__or2_1 _10206_ (.A(_04514_),
    .B(_04516_),
    .X(_04517_));
 sky130_fd_sc_hd__nand2_1 _10207_ (.A(_04516_),
    .B(_04514_),
    .Y(_04518_));
 sky130_fd_sc_hd__and2_1 _10208_ (.A(net198),
    .B(_04518_),
    .X(_04519_));
 sky130_fd_sc_hd__clkbuf_1 _10209_ (.A(net199),
    .X(\absum[4] ));
 sky130_fd_sc_hd__or2_1 _10210_ (.A(net93),
    .B(net171),
    .X(_04521_));
 sky130_fd_sc_hd__nand2_1 _10211_ (.A(net93),
    .B(net171),
    .Y(_04522_));
 sky130_fd_sc_hd__and2_1 _10212_ (.A(_04521_),
    .B(net172),
    .X(_04523_));
 sky130_fd_sc_hd__nand2_1 _10213_ (.A(_04518_),
    .B(net177),
    .Y(_04524_));
 sky130_fd_sc_hd__or2_1 _10214_ (.A(_04523_),
    .B(net178),
    .X(_04525_));
 sky130_fd_sc_hd__nand2_1 _10215_ (.A(net178),
    .B(_04523_),
    .Y(_04526_));
 sky130_fd_sc_hd__and2_1 _10216_ (.A(net179),
    .B(_04526_),
    .X(_04527_));
 sky130_fd_sc_hd__clkbuf_1 _10217_ (.A(net180),
    .X(\absum[5] ));
 sky130_fd_sc_hd__or2_1 _10218_ (.A(net94),
    .B(net136),
    .X(_04528_));
 sky130_fd_sc_hd__nand2_1 _10219_ (.A(net94),
    .B(net136),
    .Y(_04530_));
 sky130_fd_sc_hd__and2_1 _10220_ (.A(_04528_),
    .B(net137),
    .X(_04531_));
 sky130_fd_sc_hd__nand2_1 _10221_ (.A(_04526_),
    .B(net172),
    .Y(_04532_));
 sky130_fd_sc_hd__or2_1 _10222_ (.A(_04531_),
    .B(net173),
    .X(_04533_));
 sky130_fd_sc_hd__nand2_1 _10223_ (.A(net173),
    .B(_04531_),
    .Y(_04534_));
 sky130_fd_sc_hd__and2_1 _10224_ (.A(net174),
    .B(_04534_),
    .X(_04535_));
 sky130_fd_sc_hd__clkbuf_1 _10225_ (.A(net175),
    .X(\absum[6] ));
 sky130_fd_sc_hd__nor2_1 _10226_ (.A(net95),
    .B(net190),
    .Y(_04536_));
 sky130_fd_sc_hd__nand2_1 _10227_ (.A(net95),
    .B(net190),
    .Y(_04537_));
 sky130_fd_sc_hd__and2b_1 _10228_ (.A_N(_04536_),
    .B(_04537_),
    .X(_04538_));
 sky130_fd_sc_hd__nand2_1 _10229_ (.A(_04534_),
    .B(net137),
    .Y(_04540_));
 sky130_fd_sc_hd__xor2_1 _10230_ (.A(_04538_),
    .B(net138),
    .X(\absum[7] ));
 sky130_fd_sc_hd__nor2_1 _10231_ (.A(net96),
    .B(net140),
    .Y(_04541_));
 sky130_fd_sc_hd__nand2_1 _10232_ (.A(net96),
    .B(net140),
    .Y(_04542_));
 sky130_fd_sc_hd__inv_2 _10233_ (.A(net141),
    .Y(_04543_));
 sky130_fd_sc_hd__nor2_1 _10234_ (.A(_04541_),
    .B(_04543_),
    .Y(_04544_));
 sky130_fd_sc_hd__inv_2 _10235_ (.A(net138),
    .Y(_04545_));
 sky130_fd_sc_hd__o21ai_2 _10236_ (.A1(_04536_),
    .A2(_04545_),
    .B1(net191),
    .Y(_04546_));
 sky130_fd_sc_hd__or2_1 _10237_ (.A(_04544_),
    .B(net192),
    .X(_04547_));
 sky130_fd_sc_hd__nand2_1 _10238_ (.A(net192),
    .B(_04544_),
    .Y(_04548_));
 sky130_fd_sc_hd__and2_1 _10239_ (.A(net193),
    .B(_04548_),
    .X(_04550_));
 sky130_fd_sc_hd__clkbuf_1 _10240_ (.A(net194),
    .X(\absum[8] ));
 sky130_fd_sc_hd__nor2_1 _10241_ (.A(net97),
    .B(\abprod[9] ),
    .Y(_04551_));
 sky130_fd_sc_hd__nand2_1 _10242_ (.A(net97),
    .B(\abprod[9] ),
    .Y(_04552_));
 sky130_fd_sc_hd__and2b_1 _10243_ (.A_N(_04551_),
    .B(_04552_),
    .X(_04553_));
 sky130_fd_sc_hd__nand2_1 _10244_ (.A(_04548_),
    .B(net141),
    .Y(_04554_));
 sky130_fd_sc_hd__xor2_1 _10245_ (.A(_04553_),
    .B(net142),
    .X(\absum[9] ));
 sky130_fd_sc_hd__nor2_1 _10246_ (.A(net200),
    .B(net124),
    .Y(_04555_));
 sky130_fd_sc_hd__nand2_1 _10247_ (.A(net67),
    .B(net124),
    .Y(_04556_));
 sky130_fd_sc_hd__inv_2 _10248_ (.A(net125),
    .Y(_04557_));
 sky130_fd_sc_hd__nor2_1 _10249_ (.A(_04555_),
    .B(_04557_),
    .Y(_04559_));
 sky130_fd_sc_hd__and2_1 _10250_ (.A(_04553_),
    .B(_04544_),
    .X(_04560_));
 sky130_fd_sc_hd__o21ai_1 _10251_ (.A1(_04542_),
    .A2(_04551_),
    .B1(_04552_),
    .Y(_04561_));
 sky130_fd_sc_hd__a21o_1 _10252_ (.A1(_04546_),
    .A2(_04560_),
    .B1(_04561_),
    .X(_04562_));
 sky130_fd_sc_hd__or2_1 _10253_ (.A(_04559_),
    .B(_04562_),
    .X(_04563_));
 sky130_fd_sc_hd__nand2_1 _10254_ (.A(_04562_),
    .B(_04559_),
    .Y(_04564_));
 sky130_fd_sc_hd__and2_1 _10255_ (.A(_04563_),
    .B(net201),
    .X(_04565_));
 sky130_fd_sc_hd__clkbuf_1 _10256_ (.A(net202),
    .X(\absum[10] ));
 sky130_fd_sc_hd__nor2_1 _10257_ (.A(net68),
    .B(net203),
    .Y(_04566_));
 sky130_fd_sc_hd__nand2_1 _10258_ (.A(net68),
    .B(net203),
    .Y(_04567_));
 sky130_fd_sc_hd__inv_2 _10259_ (.A(net204),
    .Y(_04569_));
 sky130_fd_sc_hd__nor2_1 _10260_ (.A(_04566_),
    .B(_04569_),
    .Y(_04570_));
 sky130_fd_sc_hd__nand2_1 _10261_ (.A(_04564_),
    .B(net125),
    .Y(_04571_));
 sky130_fd_sc_hd__xor2_1 _10262_ (.A(_04570_),
    .B(net126),
    .X(\absum[11] ));
 sky130_fd_sc_hd__nor2_1 _10263_ (.A(net69),
    .B(net132),
    .Y(_04572_));
 sky130_fd_sc_hd__nand2_1 _10264_ (.A(net69),
    .B(net132),
    .Y(_04573_));
 sky130_fd_sc_hd__and2b_1 _10265_ (.A_N(_04572_),
    .B(net133),
    .X(_04574_));
 sky130_fd_sc_hd__and2_1 _10266_ (.A(_04559_),
    .B(_04570_),
    .X(_04575_));
 sky130_fd_sc_hd__nand2_1 _10267_ (.A(_04560_),
    .B(_04575_),
    .Y(_04576_));
 sky130_fd_sc_hd__inv_2 _10268_ (.A(_04546_),
    .Y(_04577_));
 sky130_fd_sc_hd__a221oi_2 _10269_ (.A1(_04557_),
    .A2(_04570_),
    .B1(_04575_),
    .B2(_04561_),
    .C1(_04569_),
    .Y(_04579_));
 sky130_fd_sc_hd__o21ai_1 _10270_ (.A1(_04576_),
    .A2(_04577_),
    .B1(net205),
    .Y(_04580_));
 sky130_fd_sc_hd__or2_1 _10271_ (.A(_04574_),
    .B(_04580_),
    .X(_04581_));
 sky130_fd_sc_hd__nand2_1 _10272_ (.A(_04580_),
    .B(_04574_),
    .Y(_04582_));
 sky130_fd_sc_hd__and2_1 _10273_ (.A(net206),
    .B(_04582_),
    .X(_04583_));
 sky130_fd_sc_hd__clkbuf_1 _10274_ (.A(net207),
    .X(\absum[12] ));
 sky130_fd_sc_hd__nor2_1 _10275_ (.A(net70),
    .B(net181),
    .Y(_04584_));
 sky130_fd_sc_hd__nand2_1 _10276_ (.A(net70),
    .B(net181),
    .Y(_04585_));
 sky130_fd_sc_hd__and2b_1 _10277_ (.A_N(_04584_),
    .B(_04585_),
    .X(_04586_));
 sky130_fd_sc_hd__nand2_1 _10278_ (.A(_04582_),
    .B(net133),
    .Y(_04587_));
 sky130_fd_sc_hd__xor2_1 _10279_ (.A(_04586_),
    .B(net134),
    .X(\absum[13] ));
 sky130_fd_sc_hd__nor2_1 _10280_ (.A(net71),
    .B(net128),
    .Y(_04589_));
 sky130_fd_sc_hd__nand2_1 _10281_ (.A(net71),
    .B(net128),
    .Y(_04590_));
 sky130_fd_sc_hd__inv_2 _10282_ (.A(net129),
    .Y(_04591_));
 sky130_fd_sc_hd__nor2_1 _10283_ (.A(_04589_),
    .B(_04591_),
    .Y(_04592_));
 sky130_fd_sc_hd__inv_2 _10284_ (.A(_04592_),
    .Y(_04593_));
 sky130_fd_sc_hd__a31o_1 _10285_ (.A1(_04582_),
    .A2(net133),
    .A3(_04585_),
    .B1(net182),
    .X(_04594_));
 sky130_fd_sc_hd__or2_1 _10286_ (.A(_04593_),
    .B(net183),
    .X(_04595_));
 sky130_fd_sc_hd__nand2_1 _10287_ (.A(net183),
    .B(_04593_),
    .Y(_04596_));
 sky130_fd_sc_hd__and2_1 _10288_ (.A(_04595_),
    .B(net184),
    .X(_04597_));
 sky130_fd_sc_hd__clkbuf_1 _10289_ (.A(net185),
    .X(\absum[14] ));
 sky130_fd_sc_hd__nor2_1 _10290_ (.A(net72),
    .B(net214),
    .Y(_04599_));
 sky130_fd_sc_hd__nand2_1 _10291_ (.A(net72),
    .B(net214),
    .Y(_04600_));
 sky130_fd_sc_hd__and2b_1 _10292_ (.A_N(_04599_),
    .B(_04600_),
    .X(_04601_));
 sky130_fd_sc_hd__nand2_1 _10293_ (.A(_04595_),
    .B(net129),
    .Y(_04602_));
 sky130_fd_sc_hd__xor2_1 _10294_ (.A(_04601_),
    .B(net130),
    .X(\absum[15] ));
 sky130_fd_sc_hd__nor2_1 _10295_ (.A(net73),
    .B(net110),
    .Y(_04603_));
 sky130_fd_sc_hd__nand2_1 _10296_ (.A(net73),
    .B(net110),
    .Y(_04604_));
 sky130_fd_sc_hd__and2b_1 _10297_ (.A_N(_04603_),
    .B(net111),
    .X(_04605_));
 sky130_fd_sc_hd__nand2_1 _10298_ (.A(_04601_),
    .B(_04592_),
    .Y(_04606_));
 sky130_fd_sc_hd__nand3b_1 _10299_ (.A_N(_04606_),
    .B(_04574_),
    .C(_04586_),
    .Y(_04608_));
 sky130_fd_sc_hd__o21a_1 _10300_ (.A1(_04573_),
    .A2(_04584_),
    .B1(_04585_),
    .X(_04609_));
 sky130_fd_sc_hd__o21a_1 _10301_ (.A1(_04590_),
    .A2(_04599_),
    .B1(net215),
    .X(_04610_));
 sky130_fd_sc_hd__o221a_1 _10302_ (.A1(_04609_),
    .A2(_04606_),
    .B1(_04608_),
    .B2(_04579_),
    .C1(_04610_),
    .X(_04611_));
 sky130_fd_sc_hd__o31ai_2 _10303_ (.A1(_04576_),
    .A2(_04608_),
    .A3(_04577_),
    .B1(_04611_),
    .Y(_04612_));
 sky130_fd_sc_hd__or2_1 _10304_ (.A(_04605_),
    .B(_04612_),
    .X(_04613_));
 sky130_fd_sc_hd__nand2_1 _10305_ (.A(_04612_),
    .B(_04605_),
    .Y(_04614_));
 sky130_fd_sc_hd__and2_1 _10306_ (.A(net216),
    .B(_04614_),
    .X(_04615_));
 sky130_fd_sc_hd__clkbuf_1 _10307_ (.A(net217),
    .X(\absum[16] ));
 sky130_fd_sc_hd__nor2_1 _10308_ (.A(net74),
    .B(net218),
    .Y(_04616_));
 sky130_fd_sc_hd__nand2_1 _10309_ (.A(net74),
    .B(net218),
    .Y(_04618_));
 sky130_fd_sc_hd__and2b_1 _10310_ (.A_N(_04616_),
    .B(_04618_),
    .X(_04619_));
 sky130_fd_sc_hd__nand2_1 _10311_ (.A(_04614_),
    .B(net111),
    .Y(_04620_));
 sky130_fd_sc_hd__xor2_1 _10312_ (.A(_04619_),
    .B(net112),
    .X(\absum[17] ));
 sky130_fd_sc_hd__nor2_1 _10313_ (.A(net75),
    .B(net114),
    .Y(_04621_));
 sky130_fd_sc_hd__nand2_1 _10314_ (.A(net75),
    .B(net114),
    .Y(_04622_));
 sky130_fd_sc_hd__and2b_1 _10315_ (.A_N(_04621_),
    .B(net115),
    .X(_04623_));
 sky130_fd_sc_hd__o21ai_1 _10316_ (.A1(net111),
    .A2(_04616_),
    .B1(net219),
    .Y(_04624_));
 sky130_fd_sc_hd__a31o_1 _10317_ (.A1(_04612_),
    .A2(_04605_),
    .A3(_04619_),
    .B1(net220),
    .X(_04625_));
 sky130_fd_sc_hd__or2_1 _10318_ (.A(_04623_),
    .B(_04625_),
    .X(_04626_));
 sky130_fd_sc_hd__nand2_1 _10319_ (.A(_04625_),
    .B(_04623_),
    .Y(_04628_));
 sky130_fd_sc_hd__and2_1 _10320_ (.A(net221),
    .B(_04628_),
    .X(_04629_));
 sky130_fd_sc_hd__clkbuf_1 _10321_ (.A(net222),
    .X(\absum[18] ));
 sky130_fd_sc_hd__nor2_1 _10322_ (.A(net76),
    .B(net208),
    .Y(_04630_));
 sky130_fd_sc_hd__nand2_1 _10323_ (.A(net76),
    .B(net208),
    .Y(_04631_));
 sky130_fd_sc_hd__and2b_1 _10324_ (.A_N(_04630_),
    .B(_04631_),
    .X(_04632_));
 sky130_fd_sc_hd__nand2_1 _10325_ (.A(_04628_),
    .B(net115),
    .Y(_04633_));
 sky130_fd_sc_hd__xor2_1 _10326_ (.A(_04632_),
    .B(net116),
    .X(\absum[19] ));
 sky130_fd_sc_hd__or2_1 _10327_ (.A(net78),
    .B(net106),
    .X(_04634_));
 sky130_fd_sc_hd__nand2_1 _10328_ (.A(net78),
    .B(net106),
    .Y(_04635_));
 sky130_fd_sc_hd__and2_1 _10329_ (.A(_04634_),
    .B(net107),
    .X(_04637_));
 sky130_fd_sc_hd__o21ai_1 _10330_ (.A1(net115),
    .A2(_04630_),
    .B1(net209),
    .Y(_04638_));
 sky130_fd_sc_hd__a31o_1 _10331_ (.A1(_04625_),
    .A2(_04623_),
    .A3(_04632_),
    .B1(net210),
    .X(_04639_));
 sky130_fd_sc_hd__or2_1 _10332_ (.A(_04637_),
    .B(net211),
    .X(_04640_));
 sky130_fd_sc_hd__nand2_1 _10333_ (.A(_04639_),
    .B(_04637_),
    .Y(_04641_));
 sky130_fd_sc_hd__and2_1 _10334_ (.A(net212),
    .B(_04641_),
    .X(_04642_));
 sky130_fd_sc_hd__clkbuf_1 _10335_ (.A(net213),
    .X(\absum[20] ));
 sky130_fd_sc_hd__nor2_1 _10336_ (.A(net79),
    .B(\abprod[21] ),
    .Y(_04643_));
 sky130_fd_sc_hd__nand2_1 _10337_ (.A(net79),
    .B(\abprod[21] ),
    .Y(_04644_));
 sky130_fd_sc_hd__and2b_1 _10338_ (.A_N(_04643_),
    .B(_04644_),
    .X(_04645_));
 sky130_fd_sc_hd__nand2_1 _10339_ (.A(_04641_),
    .B(net107),
    .Y(_04647_));
 sky130_fd_sc_hd__xor2_1 _10340_ (.A(_04645_),
    .B(net108),
    .X(\absum[21] ));
 sky130_fd_sc_hd__o21ai_1 _10341_ (.A1(net107),
    .A2(_04643_),
    .B1(_04644_),
    .Y(_04648_));
 sky130_fd_sc_hd__a31o_1 _10342_ (.A1(_04639_),
    .A2(_04637_),
    .A3(_04645_),
    .B1(_04648_),
    .X(_04649_));
 sky130_fd_sc_hd__or2_1 _10343_ (.A(net167),
    .B(_04649_),
    .X(_04650_));
 sky130_fd_sc_hd__nand2_1 _10344_ (.A(_04649_),
    .B(net167),
    .Y(_04651_));
 sky130_fd_sc_hd__and2_1 _10345_ (.A(net168),
    .B(_04651_),
    .X(_04652_));
 sky130_fd_sc_hd__clkbuf_1 _10346_ (.A(net169),
    .X(\absum[22] ));
 sky130_fd_sc_hd__inv_2 _10347_ (.A(net147),
    .Y(_04653_));
 sky130_fd_sc_hd__nor2_2 _10348_ (.A(_04653_),
    .B(_04651_),
    .Y(_04654_));
 sky130_fd_sc_hd__and2_1 _10349_ (.A(_04651_),
    .B(_04653_),
    .X(_04656_));
 sky130_fd_sc_hd__nor2_1 _10350_ (.A(_04654_),
    .B(net148),
    .Y(\absum[23] ));
 sky130_fd_sc_hd__or2_1 _10351_ (.A(net164),
    .B(_04654_),
    .X(_04657_));
 sky130_fd_sc_hd__nand2_1 _10352_ (.A(_04654_),
    .B(net164),
    .Y(_04658_));
 sky130_fd_sc_hd__and2_1 _10353_ (.A(net165),
    .B(_04658_),
    .X(_04659_));
 sky130_fd_sc_hd__clkbuf_1 _10354_ (.A(net166),
    .X(\absum[24] ));
 sky130_fd_sc_hd__inv_2 _10355_ (.A(net150),
    .Y(_04660_));
 sky130_fd_sc_hd__nor2_1 _10356_ (.A(_04660_),
    .B(_04658_),
    .Y(_04661_));
 sky130_fd_sc_hd__and2_1 _10357_ (.A(_04658_),
    .B(_04660_),
    .X(_04662_));
 sky130_fd_sc_hd__nor2_1 _10358_ (.A(_04661_),
    .B(net151),
    .Y(\absum[25] ));
 sky130_fd_sc_hd__or2_1 _10359_ (.A(net161),
    .B(_04661_),
    .X(_04664_));
 sky130_fd_sc_hd__nand2_1 _10360_ (.A(_04661_),
    .B(net161),
    .Y(_04665_));
 sky130_fd_sc_hd__and2_1 _10361_ (.A(net162),
    .B(_04665_),
    .X(_04666_));
 sky130_fd_sc_hd__clkbuf_1 _10362_ (.A(net163),
    .X(\absum[26] ));
 sky130_fd_sc_hd__inv_2 _10363_ (.A(net158),
    .Y(_04667_));
 sky130_fd_sc_hd__nor2_1 _10364_ (.A(_04667_),
    .B(_04665_),
    .Y(_04668_));
 sky130_fd_sc_hd__nand2_1 _10365_ (.A(_04665_),
    .B(_04667_),
    .Y(_04669_));
 sky130_fd_sc_hd__and2b_1 _10366_ (.A_N(_04668_),
    .B(net159),
    .X(_04670_));
 sky130_fd_sc_hd__clkbuf_1 _10367_ (.A(net160),
    .X(\absum[27] ));
 sky130_fd_sc_hd__nor2_1 _10368_ (.A(net170),
    .B(_04668_),
    .Y(_04671_));
 sky130_fd_sc_hd__and4_1 _10369_ (.A(net164),
    .B(net150),
    .C(net161),
    .D(net158),
    .X(_04673_));
 sky130_fd_sc_hd__nand3_1 _10370_ (.A(_04654_),
    .B(net170),
    .C(_04673_),
    .Y(_04674_));
 sky130_fd_sc_hd__and2b_1 _10371_ (.A_N(_04671_),
    .B(_04674_),
    .X(_04675_));
 sky130_fd_sc_hd__clkbuf_1 _10372_ (.A(_04675_),
    .X(\absum[28] ));
 sky130_fd_sc_hd__xnor2_1 _10373_ (.A(net102),
    .B(_04674_),
    .Y(\absum[29] ));
 sky130_fd_sc_hd__inv_2 _10374_ (.A(net122),
    .Y(_04676_));
 sky130_fd_sc_hd__nand2_1 _10375_ (.A(net86),
    .B(net102),
    .Y(_04677_));
 sky130_fd_sc_hd__nand3b_1 _10376_ (.A_N(_04677_),
    .B(_04654_),
    .C(_04673_),
    .Y(_04678_));
 sky130_fd_sc_hd__xor2_1 _10377_ (.A(_04676_),
    .B(_04678_),
    .X(\absum[30] ));
 sky130_fd_sc_hd__nor2_1 _10378_ (.A(_04676_),
    .B(_04678_),
    .Y(_04679_));
 sky130_fd_sc_hd__xor2_1 _10379_ (.A(net104),
    .B(_04679_),
    .X(\absum[31] ));
 sky130_fd_sc_hd__or2_1 _10380_ (.A(net66),
    .B(net144),
    .X(_04681_));
 sky130_fd_sc_hd__and2_1 _10381_ (.A(net145),
    .B(_04489_),
    .X(_04682_));
 sky130_fd_sc_hd__clkbuf_1 _10382_ (.A(net146),
    .X(\absum[0] ));
 sky130_fd_sc_hd__and3_1 _10383_ (.A(_02299_),
    .B(_02268_),
    .C(_02267_),
    .X(_04683_));
 sky130_fd_sc_hd__nand3b_1 _10384_ (.A_N(_02272_),
    .B(_02304_),
    .C(_04683_),
    .Y(_04684_));
 sky130_fd_sc_hd__or3_1 _10385_ (.A(_02308_),
    .B(_02241_),
    .C(_04684_),
    .X(_04685_));
 sky130_fd_sc_hd__or2_1 _10386_ (.A(_02282_),
    .B(_04685_),
    .X(_04686_));
 sky130_fd_sc_hd__nand2_1 _10387_ (.A(_04685_),
    .B(_02282_),
    .Y(_04687_));
 sky130_fd_sc_hd__and2_1 _10388_ (.A(_04686_),
    .B(_04687_),
    .X(_04688_));
 sky130_fd_sc_hd__clkbuf_1 _10389_ (.A(_04688_),
    .X(\ab[0] ));
 sky130_fd_sc_hd__nand2_1 _10390_ (.A(_04686_),
    .B(_02281_),
    .Y(_04690_));
 sky130_fd_sc_hd__xnor2_1 _10391_ (.A(_02289_),
    .B(_04690_),
    .Y(\ab[1] ));
 sky130_fd_sc_hd__o21ai_1 _10392_ (.A1(_02289_),
    .A2(_04686_),
    .B1(_02314_),
    .Y(_04691_));
 sky130_fd_sc_hd__or2_1 _10393_ (.A(_02185_),
    .B(_04691_),
    .X(_04692_));
 sky130_fd_sc_hd__nand2_1 _10394_ (.A(_04691_),
    .B(_02185_),
    .Y(_04693_));
 sky130_fd_sc_hd__and2_1 _10395_ (.A(_04692_),
    .B(_04693_),
    .X(_04694_));
 sky130_fd_sc_hd__clkbuf_1 _10396_ (.A(_04694_),
    .X(\ab[2] ));
 sky130_fd_sc_hd__nand2_1 _10397_ (.A(_04693_),
    .B(_02182_),
    .Y(_04695_));
 sky130_fd_sc_hd__xor2_1 _10398_ (.A(_02187_),
    .B(_04695_),
    .X(\ab[3] ));
 sky130_fd_sc_hd__a21o_1 _10399_ (.A1(_02311_),
    .A2(_02314_),
    .B1(_02188_),
    .X(_04697_));
 sky130_fd_sc_hd__nand2_1 _10400_ (.A(_04697_),
    .B(_02172_),
    .Y(_04698_));
 sky130_fd_sc_hd__or2_1 _10401_ (.A(_02176_),
    .B(_04698_),
    .X(_04699_));
 sky130_fd_sc_hd__nand2_1 _10402_ (.A(_04698_),
    .B(_02176_),
    .Y(_04700_));
 sky130_fd_sc_hd__and2_1 _10403_ (.A(_04699_),
    .B(_04700_),
    .X(_04701_));
 sky130_fd_sc_hd__clkbuf_1 _10404_ (.A(_04701_),
    .X(\ab[4] ));
 sky130_fd_sc_hd__nand2_1 _10405_ (.A(_04700_),
    .B(_01998_),
    .Y(_04702_));
 sky130_fd_sc_hd__xnor2_1 _10406_ (.A(_02006_),
    .B(_04702_),
    .Y(\ab[5] ));
 sky130_fd_sc_hd__xor2_1 _10407_ (.A(_02323_),
    .B(_02317_),
    .X(\ab[6] ));
 sky130_fd_sc_hd__a21bo_1 _10408_ (.A1(_02317_),
    .A2(_02321_),
    .B1_N(_01712_),
    .X(_04703_));
 sky130_fd_sc_hd__xor2_1 _10409_ (.A(_02319_),
    .B(_04703_),
    .X(\ab[7] ));
 sky130_fd_sc_hd__inv_2 _10410_ (.A(_01766_),
    .Y(_04705_));
 sky130_fd_sc_hd__a31o_1 _10411_ (.A1(_02317_),
    .A2(_02319_),
    .A3(_02323_),
    .B1(_01740_),
    .X(_04706_));
 sky130_fd_sc_hd__or2_1 _10412_ (.A(_04705_),
    .B(_04706_),
    .X(_04707_));
 sky130_fd_sc_hd__nand2_1 _10413_ (.A(_04706_),
    .B(_04705_),
    .Y(_04708_));
 sky130_fd_sc_hd__and2_1 _10414_ (.A(_04707_),
    .B(_04708_),
    .X(_04709_));
 sky130_fd_sc_hd__clkbuf_1 _10415_ (.A(_04709_),
    .X(\ab[8] ));
 sky130_fd_sc_hd__nand2_1 _10416_ (.A(_04708_),
    .B(_01765_),
    .Y(_04710_));
 sky130_fd_sc_hd__xnor2_1 _10417_ (.A(_01758_),
    .B(_04710_),
    .Y(\ab[9] ));
 sky130_fd_sc_hd__inv_2 _10418_ (.A(_01773_),
    .Y(_04711_));
 sky130_fd_sc_hd__a21bo_1 _10419_ (.A1(_02317_),
    .A2(_02325_),
    .B1_N(_01770_),
    .X(_04713_));
 sky130_fd_sc_hd__or2_1 _10420_ (.A(_04711_),
    .B(_04713_),
    .X(_04714_));
 sky130_fd_sc_hd__nand2_1 _10421_ (.A(_04713_),
    .B(_04711_),
    .Y(_04715_));
 sky130_fd_sc_hd__and2_1 _10422_ (.A(_04714_),
    .B(_04715_),
    .X(_04716_));
 sky130_fd_sc_hd__clkbuf_1 _10423_ (.A(_04716_),
    .X(\ab[10] ));
 sky130_fd_sc_hd__nand2_1 _10424_ (.A(_04715_),
    .B(_01162_),
    .Y(_04717_));
 sky130_fd_sc_hd__xnor2_1 _10425_ (.A(_01777_),
    .B(_04717_),
    .Y(\ab[11] ));
 sky130_fd_sc_hd__inv_2 _10426_ (.A(_00798_),
    .Y(_04718_));
 sky130_fd_sc_hd__nand2_1 _10427_ (.A(_04713_),
    .B(_01778_),
    .Y(_04719_));
 sky130_fd_sc_hd__or2_1 _10428_ (.A(_01162_),
    .B(_01777_),
    .X(_04720_));
 sky130_fd_sc_hd__nand3_1 _10429_ (.A(_04719_),
    .B(_01167_),
    .C(_04720_),
    .Y(_04722_));
 sky130_fd_sc_hd__or2_1 _10430_ (.A(_04718_),
    .B(_04722_),
    .X(_04723_));
 sky130_fd_sc_hd__nand2_1 _10431_ (.A(_04722_),
    .B(_04718_),
    .Y(_04724_));
 sky130_fd_sc_hd__and2_1 _10432_ (.A(_04723_),
    .B(_04724_),
    .X(_04725_));
 sky130_fd_sc_hd__clkbuf_1 _10433_ (.A(_04725_),
    .X(\ab[12] ));
 sky130_fd_sc_hd__nand2_1 _10434_ (.A(_04724_),
    .B(_00797_),
    .Y(_04726_));
 sky130_fd_sc_hd__xnor2_1 _10435_ (.A(_00611_),
    .B(_04726_),
    .Y(\ab[13] ));
 sky130_fd_sc_hd__or2_1 _10436_ (.A(_02832_),
    .B(_02327_),
    .X(_04727_));
 sky130_fd_sc_hd__nand2_1 _10437_ (.A(_02327_),
    .B(_02832_),
    .Y(_04728_));
 sky130_fd_sc_hd__and2_1 _10438_ (.A(_04727_),
    .B(_04728_),
    .X(_04729_));
 sky130_fd_sc_hd__clkbuf_1 _10439_ (.A(_04729_),
    .X(\ab[14] ));
 sky130_fd_sc_hd__nand2_1 _10440_ (.A(_04728_),
    .B(_02829_),
    .Y(_04731_));
 sky130_fd_sc_hd__xor2_1 _10441_ (.A(_02823_),
    .B(_04731_),
    .X(\ab[15] ));
 sky130_fd_sc_hd__inv_2 _10442_ (.A(_02833_),
    .Y(_04732_));
 sky130_fd_sc_hd__a21o_1 _10443_ (.A1(_02327_),
    .A2(_04732_),
    .B1(_03404_),
    .X(_04733_));
 sky130_fd_sc_hd__or2_1 _10444_ (.A(_03397_),
    .B(_04733_),
    .X(_04734_));
 sky130_fd_sc_hd__nand2_1 _10445_ (.A(_04733_),
    .B(_03397_),
    .Y(_04735_));
 sky130_fd_sc_hd__and2_1 _10446_ (.A(_04734_),
    .B(_04735_),
    .X(_04736_));
 sky130_fd_sc_hd__clkbuf_1 _10447_ (.A(_04736_),
    .X(\ab[16] ));
 sky130_fd_sc_hd__nand2_1 _10448_ (.A(_04735_),
    .B(_03395_),
    .Y(_04737_));
 sky130_fd_sc_hd__xor2_1 _10449_ (.A(_03389_),
    .B(_04737_),
    .X(\ab[17] ));
 sky130_fd_sc_hd__inv_2 _10450_ (.A(_03670_),
    .Y(_04739_));
 sky130_fd_sc_hd__or2_1 _10451_ (.A(_04739_),
    .B(_03410_),
    .X(_04740_));
 sky130_fd_sc_hd__nand2_1 _10452_ (.A(_03410_),
    .B(_04739_),
    .Y(_04741_));
 sky130_fd_sc_hd__and2_1 _10453_ (.A(_04740_),
    .B(_04741_),
    .X(_04742_));
 sky130_fd_sc_hd__buf_1 _10454_ (.A(_04742_),
    .X(\ab[18] ));
 sky130_fd_sc_hd__nand2_1 _10455_ (.A(_04741_),
    .B(_03669_),
    .Y(_04743_));
 sky130_fd_sc_hd__xnor2_1 _10456_ (.A(_03938_),
    .B(_04743_),
    .Y(\ab[19] ));
 sky130_fd_sc_hd__xor2_1 _10457_ (.A(_04233_),
    .B(_03944_),
    .X(\ab[20] ));
 sky130_fd_sc_hd__dfrtp_1 _10458_ (.CLK(clknet_2_0__leaf_clk),
    .D(\ab[0] ),
    .RESET_B(net98),
    .Q(\abprod[0] ));
 sky130_fd_sc_hd__dfrtp_1 _10459_ (.CLK(clknet_2_1__leaf_clk),
    .D(\ab[1] ),
    .RESET_B(net98),
    .Q(\abprod[1] ));
 sky130_fd_sc_hd__dfrtp_1 _10460_ (.CLK(clknet_2_0__leaf_clk),
    .D(\ab[2] ),
    .RESET_B(net98),
    .Q(\abprod[2] ));
 sky130_fd_sc_hd__dfrtp_1 _10461_ (.CLK(clknet_2_1__leaf_clk),
    .D(\ab[3] ),
    .RESET_B(net98),
    .Q(\abprod[3] ));
 sky130_fd_sc_hd__dfrtp_1 _10462_ (.CLK(clknet_2_0__leaf_clk),
    .D(\ab[4] ),
    .RESET_B(net98),
    .Q(\abprod[4] ));
 sky130_fd_sc_hd__dfrtp_1 _10463_ (.CLK(clknet_2_1__leaf_clk),
    .D(\ab[5] ),
    .RESET_B(net98),
    .Q(\abprod[5] ));
 sky130_fd_sc_hd__dfrtp_1 _10464_ (.CLK(clknet_2_0__leaf_clk),
    .D(\ab[6] ),
    .RESET_B(net98),
    .Q(\abprod[6] ));
 sky130_fd_sc_hd__dfrtp_1 _10465_ (.CLK(clknet_2_1__leaf_clk),
    .D(\ab[7] ),
    .RESET_B(net98),
    .Q(\abprod[7] ));
 sky130_fd_sc_hd__dfrtp_1 _10466_ (.CLK(clknet_2_0__leaf_clk),
    .D(\ab[8] ),
    .RESET_B(net98),
    .Q(\abprod[8] ));
 sky130_fd_sc_hd__dfrtp_1 _10467_ (.CLK(clknet_2_1__leaf_clk),
    .D(\ab[9] ),
    .RESET_B(net99),
    .Q(\abprod[9] ));
 sky130_fd_sc_hd__dfrtp_1 _10468_ (.CLK(clknet_2_0__leaf_clk),
    .D(\ab[10] ),
    .RESET_B(net99),
    .Q(\abprod[10] ));
 sky130_fd_sc_hd__dfrtp_1 _10469_ (.CLK(clknet_2_1__leaf_clk),
    .D(\ab[11] ),
    .RESET_B(net99),
    .Q(\abprod[11] ));
 sky130_fd_sc_hd__dfrtp_1 _10470_ (.CLK(clknet_2_0__leaf_clk),
    .D(\ab[12] ),
    .RESET_B(net99),
    .Q(\abprod[12] ));
 sky130_fd_sc_hd__dfrtp_1 _10471_ (.CLK(clknet_2_1__leaf_clk),
    .D(\ab[13] ),
    .RESET_B(net99),
    .Q(\abprod[13] ));
 sky130_fd_sc_hd__dfrtp_1 _10472_ (.CLK(clknet_2_0__leaf_clk),
    .D(\ab[14] ),
    .RESET_B(net99),
    .Q(\abprod[14] ));
 sky130_fd_sc_hd__dfrtp_1 _10473_ (.CLK(clknet_2_3__leaf_clk),
    .D(\ab[15] ),
    .RESET_B(net100),
    .Q(\abprod[15] ));
 sky130_fd_sc_hd__dfrtp_1 _10474_ (.CLK(clknet_2_2__leaf_clk),
    .D(\ab[16] ),
    .RESET_B(net100),
    .Q(\abprod[16] ));
 sky130_fd_sc_hd__dfrtp_1 _10475_ (.CLK(clknet_2_3__leaf_clk),
    .D(\ab[17] ),
    .RESET_B(net100),
    .Q(\abprod[17] ));
 sky130_fd_sc_hd__dfrtp_1 _10476_ (.CLK(clknet_2_2__leaf_clk),
    .D(\ab[18] ),
    .RESET_B(net100),
    .Q(\abprod[18] ));
 sky130_fd_sc_hd__dfrtp_1 _10477_ (.CLK(clknet_2_3__leaf_clk),
    .D(\ab[19] ),
    .RESET_B(net100),
    .Q(\abprod[19] ));
 sky130_fd_sc_hd__dfrtp_1 _10478_ (.CLK(clknet_2_2__leaf_clk),
    .D(\ab[20] ),
    .RESET_B(net100),
    .Q(\abprod[20] ));
 sky130_fd_sc_hd__dfrtp_1 _10479_ (.CLK(clknet_2_3__leaf_clk),
    .D(\ab[21] ),
    .RESET_B(net100),
    .Q(\abprod[21] ));
 sky130_fd_sc_hd__dfrtp_1 _10480_ (.CLK(clknet_2_0__leaf_clk),
    .D(\absum[0] ),
    .RESET_B(net98),
    .Q(net66));
 sky130_fd_sc_hd__dfrtp_2 _10481_ (.CLK(clknet_2_0__leaf_clk),
    .D(\absum[1] ),
    .RESET_B(net98),
    .Q(net77));
 sky130_fd_sc_hd__dfrtp_1 _10482_ (.CLK(clknet_2_0__leaf_clk),
    .D(\absum[2] ),
    .RESET_B(net98),
    .Q(net88));
 sky130_fd_sc_hd__dfrtp_2 _10483_ (.CLK(clknet_2_1__leaf_clk),
    .D(net121),
    .RESET_B(net98),
    .Q(net91));
 sky130_fd_sc_hd__dfrtp_1 _10484_ (.CLK(clknet_2_0__leaf_clk),
    .D(\absum[4] ),
    .RESET_B(net98),
    .Q(net92));
 sky130_fd_sc_hd__dfrtp_2 _10485_ (.CLK(clknet_2_1__leaf_clk),
    .D(\absum[5] ),
    .RESET_B(net98),
    .Q(net93));
 sky130_fd_sc_hd__dfrtp_1 _10486_ (.CLK(clknet_2_0__leaf_clk),
    .D(\absum[6] ),
    .RESET_B(net98),
    .Q(net94));
 sky130_fd_sc_hd__dfrtp_2 _10487_ (.CLK(clknet_2_1__leaf_clk),
    .D(net139),
    .RESET_B(net99),
    .Q(net95));
 sky130_fd_sc_hd__dfrtp_2 _10488_ (.CLK(clknet_2_0__leaf_clk),
    .D(\absum[8] ),
    .RESET_B(net99),
    .Q(net96));
 sky130_fd_sc_hd__dfrtp_2 _10489_ (.CLK(clknet_2_1__leaf_clk),
    .D(net143),
    .RESET_B(net99),
    .Q(net97));
 sky130_fd_sc_hd__dfrtp_1 _10490_ (.CLK(clknet_2_0__leaf_clk),
    .D(\absum[10] ),
    .RESET_B(net99),
    .Q(net67));
 sky130_fd_sc_hd__dfrtp_2 _10491_ (.CLK(clknet_2_0__leaf_clk),
    .D(net127),
    .RESET_B(net99),
    .Q(net68));
 sky130_fd_sc_hd__dfrtp_2 _10492_ (.CLK(clknet_2_0__leaf_clk),
    .D(\absum[12] ),
    .RESET_B(net99),
    .Q(net69));
 sky130_fd_sc_hd__dfrtp_2 _10493_ (.CLK(clknet_2_1__leaf_clk),
    .D(net135),
    .RESET_B(net99),
    .Q(net70));
 sky130_fd_sc_hd__dfrtp_2 _10494_ (.CLK(clknet_2_0__leaf_clk),
    .D(\absum[14] ),
    .RESET_B(net99),
    .Q(net71));
 sky130_fd_sc_hd__dfrtp_1 _10495_ (.CLK(clknet_2_1__leaf_clk),
    .D(net131),
    .RESET_B(net99),
    .Q(net72));
 sky130_fd_sc_hd__dfrtp_2 _10496_ (.CLK(clknet_2_2__leaf_clk),
    .D(\absum[16] ),
    .RESET_B(net100),
    .Q(net73));
 sky130_fd_sc_hd__dfrtp_2 _10497_ (.CLK(clknet_2_3__leaf_clk),
    .D(net113),
    .RESET_B(net100),
    .Q(net74));
 sky130_fd_sc_hd__dfrtp_2 _10498_ (.CLK(clknet_2_2__leaf_clk),
    .D(\absum[18] ),
    .RESET_B(net100),
    .Q(net75));
 sky130_fd_sc_hd__dfrtp_2 _10499_ (.CLK(clknet_2_3__leaf_clk),
    .D(net117),
    .RESET_B(net100),
    .Q(net76));
 sky130_fd_sc_hd__dfrtp_2 _10500_ (.CLK(clknet_2_2__leaf_clk),
    .D(\absum[20] ),
    .RESET_B(net100),
    .Q(net78));
 sky130_fd_sc_hd__dfrtp_2 _10501_ (.CLK(clknet_2_3__leaf_clk),
    .D(net109),
    .RESET_B(net100),
    .Q(net79));
 sky130_fd_sc_hd__dfrtp_1 _10502_ (.CLK(clknet_2_2__leaf_clk),
    .D(\absum[22] ),
    .RESET_B(net100),
    .Q(net80));
 sky130_fd_sc_hd__dfrtp_1 _10503_ (.CLK(clknet_2_3__leaf_clk),
    .D(net149),
    .RESET_B(net100),
    .Q(net81));
 sky130_fd_sc_hd__dfrtp_1 _10504_ (.CLK(clknet_2_2__leaf_clk),
    .D(\absum[24] ),
    .RESET_B(net100),
    .Q(net82));
 sky130_fd_sc_hd__dfrtp_1 _10505_ (.CLK(clknet_2_2__leaf_clk),
    .D(net152),
    .RESET_B(net101),
    .Q(net83));
 sky130_fd_sc_hd__dfrtp_1 _10506_ (.CLK(clknet_2_3__leaf_clk),
    .D(\absum[26] ),
    .RESET_B(net101),
    .Q(net84));
 sky130_fd_sc_hd__dfrtp_1 _10507_ (.CLK(clknet_2_3__leaf_clk),
    .D(\absum[27] ),
    .RESET_B(net101),
    .Q(net85));
 sky130_fd_sc_hd__dfrtp_1 _10508_ (.CLK(clknet_2_3__leaf_clk),
    .D(\absum[28] ),
    .RESET_B(net101),
    .Q(net86));
 sky130_fd_sc_hd__dfrtp_1 _10509_ (.CLK(clknet_2_3__leaf_clk),
    .D(net103),
    .RESET_B(net101),
    .Q(net87));
 sky130_fd_sc_hd__dfrtp_1 _10510_ (.CLK(clknet_2_2__leaf_clk),
    .D(net123),
    .RESET_B(net101),
    .Q(net89));
 sky130_fd_sc_hd__dfrtp_1 _10511_ (.CLK(clknet_2_2__leaf_clk),
    .D(net105),
    .RESET_B(net101),
    .Q(net90));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_0__f_clk (.A(clknet_0_clk),
    .X(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_1__f_clk (.A(clknet_0_clk),
    .X(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_2__f_clk (.A(clknet_0_clk),
    .X(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_3__f_clk (.A(clknet_0_clk),
    .X(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__clkbuf_8 fanout100 (.A(net101),
    .X(net100));
 sky130_fd_sc_hd__buf_4 fanout101 (.A(net65),
    .X(net101));
 sky130_fd_sc_hd__clkbuf_8 fanout98 (.A(net99),
    .X(net98));
 sky130_fd_sc_hd__clkbuf_8 fanout99 (.A(net101),
    .X(net99));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1 (.A(net87),
    .X(net102));
 sky130_fd_sc_hd__dlygate4sd3_1 hold10 (.A(_04604_),
    .X(net111));
 sky130_fd_sc_hd__dlygate4sd3_1 hold100 (.A(_04564_),
    .X(net201));
 sky130_fd_sc_hd__dlygate4sd3_1 hold101 (.A(_04565_),
    .X(net202));
 sky130_fd_sc_hd__dlygate4sd3_1 hold102 (.A(\abprod[11] ),
    .X(net203));
 sky130_fd_sc_hd__dlygate4sd3_1 hold103 (.A(_04567_),
    .X(net204));
 sky130_fd_sc_hd__dlygate4sd3_1 hold104 (.A(_04579_),
    .X(net205));
 sky130_fd_sc_hd__dlygate4sd3_1 hold105 (.A(_04581_),
    .X(net206));
 sky130_fd_sc_hd__dlygate4sd3_1 hold106 (.A(_04583_),
    .X(net207));
 sky130_fd_sc_hd__dlygate4sd3_1 hold107 (.A(\abprod[19] ),
    .X(net208));
 sky130_fd_sc_hd__dlygate4sd3_1 hold108 (.A(_04631_),
    .X(net209));
 sky130_fd_sc_hd__dlygate4sd3_1 hold109 (.A(_04638_),
    .X(net210));
 sky130_fd_sc_hd__dlygate4sd3_1 hold11 (.A(_04620_),
    .X(net112));
 sky130_fd_sc_hd__dlygate4sd3_1 hold110 (.A(_04639_),
    .X(net211));
 sky130_fd_sc_hd__dlygate4sd3_1 hold111 (.A(_04640_),
    .X(net212));
 sky130_fd_sc_hd__dlygate4sd3_1 hold112 (.A(_04642_),
    .X(net213));
 sky130_fd_sc_hd__dlygate4sd3_1 hold113 (.A(\abprod[15] ),
    .X(net214));
 sky130_fd_sc_hd__dlygate4sd3_1 hold114 (.A(_04600_),
    .X(net215));
 sky130_fd_sc_hd__dlygate4sd3_1 hold115 (.A(_04613_),
    .X(net216));
 sky130_fd_sc_hd__dlygate4sd3_1 hold116 (.A(_04615_),
    .X(net217));
 sky130_fd_sc_hd__dlygate4sd3_1 hold117 (.A(\abprod[17] ),
    .X(net218));
 sky130_fd_sc_hd__dlygate4sd3_1 hold118 (.A(_04618_),
    .X(net219));
 sky130_fd_sc_hd__dlygate4sd3_1 hold119 (.A(_04624_),
    .X(net220));
 sky130_fd_sc_hd__dlygate4sd3_1 hold12 (.A(\absum[17] ),
    .X(net113));
 sky130_fd_sc_hd__dlygate4sd3_1 hold120 (.A(_04626_),
    .X(net221));
 sky130_fd_sc_hd__dlygate4sd3_1 hold121 (.A(_04629_),
    .X(net222));
 sky130_fd_sc_hd__dlygate4sd3_1 hold13 (.A(\abprod[18] ),
    .X(net114));
 sky130_fd_sc_hd__dlygate4sd3_1 hold14 (.A(_04622_),
    .X(net115));
 sky130_fd_sc_hd__dlygate4sd3_1 hold15 (.A(_04633_),
    .X(net116));
 sky130_fd_sc_hd__dlygate4sd3_1 hold16 (.A(\absum[19] ),
    .X(net117));
 sky130_fd_sc_hd__dlygate4sd3_1 hold17 (.A(\abprod[2] ),
    .X(net118));
 sky130_fd_sc_hd__dlygate4sd3_1 hold18 (.A(_04501_),
    .X(net119));
 sky130_fd_sc_hd__dlygate4sd3_1 hold19 (.A(_04511_),
    .X(net120));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(\absum[29] ),
    .X(net103));
 sky130_fd_sc_hd__dlygate4sd3_1 hold20 (.A(\absum[3] ),
    .X(net121));
 sky130_fd_sc_hd__dlygate4sd3_1 hold21 (.A(net89),
    .X(net122));
 sky130_fd_sc_hd__dlygate4sd3_1 hold22 (.A(\absum[30] ),
    .X(net123));
 sky130_fd_sc_hd__dlygate4sd3_1 hold23 (.A(\abprod[10] ),
    .X(net124));
 sky130_fd_sc_hd__dlygate4sd3_1 hold24 (.A(_04556_),
    .X(net125));
 sky130_fd_sc_hd__dlygate4sd3_1 hold25 (.A(_04571_),
    .X(net126));
 sky130_fd_sc_hd__dlygate4sd3_1 hold26 (.A(\absum[11] ),
    .X(net127));
 sky130_fd_sc_hd__dlygate4sd3_1 hold27 (.A(\abprod[14] ),
    .X(net128));
 sky130_fd_sc_hd__dlygate4sd3_1 hold28 (.A(_04590_),
    .X(net129));
 sky130_fd_sc_hd__dlygate4sd3_1 hold29 (.A(_04602_),
    .X(net130));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3 (.A(net90),
    .X(net104));
 sky130_fd_sc_hd__dlygate4sd3_1 hold30 (.A(\absum[15] ),
    .X(net131));
 sky130_fd_sc_hd__dlygate4sd3_1 hold31 (.A(\abprod[12] ),
    .X(net132));
 sky130_fd_sc_hd__dlygate4sd3_1 hold32 (.A(_04573_),
    .X(net133));
 sky130_fd_sc_hd__dlygate4sd3_1 hold33 (.A(_04587_),
    .X(net134));
 sky130_fd_sc_hd__dlygate4sd3_1 hold34 (.A(\absum[13] ),
    .X(net135));
 sky130_fd_sc_hd__dlygate4sd3_1 hold35 (.A(\abprod[6] ),
    .X(net136));
 sky130_fd_sc_hd__dlygate4sd3_1 hold36 (.A(_04530_),
    .X(net137));
 sky130_fd_sc_hd__buf_1 hold37 (.A(_04540_),
    .X(net138));
 sky130_fd_sc_hd__dlygate4sd3_1 hold38 (.A(\absum[7] ),
    .X(net139));
 sky130_fd_sc_hd__dlygate4sd3_1 hold39 (.A(\abprod[8] ),
    .X(net140));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4 (.A(\absum[31] ),
    .X(net105));
 sky130_fd_sc_hd__dlygate4sd3_1 hold40 (.A(_04542_),
    .X(net141));
 sky130_fd_sc_hd__dlygate4sd3_1 hold41 (.A(_04554_),
    .X(net142));
 sky130_fd_sc_hd__dlygate4sd3_1 hold42 (.A(\absum[9] ),
    .X(net143));
 sky130_fd_sc_hd__dlygate4sd3_1 hold43 (.A(\abprod[0] ),
    .X(net144));
 sky130_fd_sc_hd__dlygate4sd3_1 hold44 (.A(_04681_),
    .X(net145));
 sky130_fd_sc_hd__dlygate4sd3_1 hold45 (.A(_04682_),
    .X(net146));
 sky130_fd_sc_hd__dlygate4sd3_1 hold46 (.A(net81),
    .X(net147));
 sky130_fd_sc_hd__dlygate4sd3_1 hold47 (.A(_04656_),
    .X(net148));
 sky130_fd_sc_hd__dlygate4sd3_1 hold48 (.A(\absum[23] ),
    .X(net149));
 sky130_fd_sc_hd__dlygate4sd3_1 hold49 (.A(net83),
    .X(net150));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5 (.A(\abprod[20] ),
    .X(net106));
 sky130_fd_sc_hd__dlygate4sd3_1 hold50 (.A(_04662_),
    .X(net151));
 sky130_fd_sc_hd__dlygate4sd3_1 hold51 (.A(\absum[25] ),
    .X(net152));
 sky130_fd_sc_hd__dlygate4sd3_1 hold52 (.A(\abprod[1] ),
    .X(net153));
 sky130_fd_sc_hd__dlygate4sd3_1 hold53 (.A(_04493_),
    .X(net154));
 sky130_fd_sc_hd__dlygate4sd3_1 hold54 (.A(_04495_),
    .X(net155));
 sky130_fd_sc_hd__dlygate4sd3_1 hold55 (.A(_04497_),
    .X(net156));
 sky130_fd_sc_hd__dlygate4sd3_1 hold56 (.A(_04498_),
    .X(net157));
 sky130_fd_sc_hd__dlygate4sd3_1 hold57 (.A(net85),
    .X(net158));
 sky130_fd_sc_hd__dlygate4sd3_1 hold58 (.A(_04669_),
    .X(net159));
 sky130_fd_sc_hd__dlygate4sd3_1 hold59 (.A(_04670_),
    .X(net160));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6 (.A(_04635_),
    .X(net107));
 sky130_fd_sc_hd__dlygate4sd3_1 hold60 (.A(net84),
    .X(net161));
 sky130_fd_sc_hd__dlygate4sd3_1 hold61 (.A(_04664_),
    .X(net162));
 sky130_fd_sc_hd__dlygate4sd3_1 hold62 (.A(_04666_),
    .X(net163));
 sky130_fd_sc_hd__dlygate4sd3_1 hold63 (.A(net82),
    .X(net164));
 sky130_fd_sc_hd__dlygate4sd3_1 hold64 (.A(_04657_),
    .X(net165));
 sky130_fd_sc_hd__dlygate4sd3_1 hold65 (.A(_04659_),
    .X(net166));
 sky130_fd_sc_hd__dlygate4sd3_1 hold66 (.A(net80),
    .X(net167));
 sky130_fd_sc_hd__dlygate4sd3_1 hold67 (.A(_04650_),
    .X(net168));
 sky130_fd_sc_hd__dlygate4sd3_1 hold68 (.A(_04652_),
    .X(net169));
 sky130_fd_sc_hd__dlygate4sd3_1 hold69 (.A(net86),
    .X(net170));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7 (.A(_04647_),
    .X(net108));
 sky130_fd_sc_hd__dlygate4sd3_1 hold70 (.A(\abprod[5] ),
    .X(net171));
 sky130_fd_sc_hd__dlygate4sd3_1 hold71 (.A(_04522_),
    .X(net172));
 sky130_fd_sc_hd__dlygate4sd3_1 hold72 (.A(_04532_),
    .X(net173));
 sky130_fd_sc_hd__dlygate4sd3_1 hold73 (.A(_04533_),
    .X(net174));
 sky130_fd_sc_hd__dlygate4sd3_1 hold74 (.A(_04535_),
    .X(net175));
 sky130_fd_sc_hd__dlygate4sd3_1 hold75 (.A(\abprod[4] ),
    .X(net176));
 sky130_fd_sc_hd__dlygate4sd3_1 hold76 (.A(_04513_),
    .X(net177));
 sky130_fd_sc_hd__dlygate4sd3_1 hold77 (.A(_04524_),
    .X(net178));
 sky130_fd_sc_hd__dlygate4sd3_1 hold78 (.A(_04525_),
    .X(net179));
 sky130_fd_sc_hd__dlygate4sd3_1 hold79 (.A(_04527_),
    .X(net180));
 sky130_fd_sc_hd__dlygate4sd3_1 hold8 (.A(\absum[21] ),
    .X(net109));
 sky130_fd_sc_hd__dlygate4sd3_1 hold80 (.A(\abprod[13] ),
    .X(net181));
 sky130_fd_sc_hd__dlygate4sd3_1 hold81 (.A(_04584_),
    .X(net182));
 sky130_fd_sc_hd__dlygate4sd3_1 hold82 (.A(_04594_),
    .X(net183));
 sky130_fd_sc_hd__dlygate4sd3_1 hold83 (.A(_04596_),
    .X(net184));
 sky130_fd_sc_hd__dlygate4sd3_1 hold84 (.A(_04597_),
    .X(net185));
 sky130_fd_sc_hd__dlygate4sd3_1 hold85 (.A(net77),
    .X(net186));
 sky130_fd_sc_hd__dlygate4sd3_1 hold86 (.A(_04503_),
    .X(net187));
 sky130_fd_sc_hd__dlygate4sd3_1 hold87 (.A(_04504_),
    .X(net188));
 sky130_fd_sc_hd__dlygate4sd3_1 hold88 (.A(_04506_),
    .X(net189));
 sky130_fd_sc_hd__dlygate4sd3_1 hold89 (.A(\abprod[7] ),
    .X(net190));
 sky130_fd_sc_hd__dlygate4sd3_1 hold9 (.A(\abprod[16] ),
    .X(net110));
 sky130_fd_sc_hd__dlygate4sd3_1 hold90 (.A(_04537_),
    .X(net191));
 sky130_fd_sc_hd__dlygate4sd3_1 hold91 (.A(_04546_),
    .X(net192));
 sky130_fd_sc_hd__dlygate4sd3_1 hold92 (.A(_04547_),
    .X(net193));
 sky130_fd_sc_hd__dlygate4sd3_1 hold93 (.A(_04550_),
    .X(net194));
 sky130_fd_sc_hd__dlygate4sd3_1 hold94 (.A(\abprod[3] ),
    .X(net195));
 sky130_fd_sc_hd__dlygate4sd3_1 hold95 (.A(_04508_),
    .X(net196));
 sky130_fd_sc_hd__dlygate4sd3_1 hold96 (.A(_04515_),
    .X(net197));
 sky130_fd_sc_hd__dlygate4sd3_1 hold97 (.A(_04517_),
    .X(net198));
 sky130_fd_sc_hd__dlygate4sd3_1 hold98 (.A(_04519_),
    .X(net199));
 sky130_fd_sc_hd__dlygate4sd3_1 hold99 (.A(net67),
    .X(net200));
 sky130_fd_sc_hd__clkbuf_4 input1 (.A(a_i[0]),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_1 input10 (.A(a_i[18]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_1 input11 (.A(a_i[19]),
    .X(net11));
 sky130_fd_sc_hd__buf_2 input12 (.A(a_i[1]),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_1 input13 (.A(a_i[20]),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_1 input14 (.A(a_i[21]),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_1 input15 (.A(a_i[22]),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_1 input16 (.A(a_i[23]),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_4 input17 (.A(a_i[24]),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_4 input18 (.A(a_i[25]),
    .X(net18));
 sky130_fd_sc_hd__buf_2 input19 (.A(a_i[26]),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(a_i[10]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_2 input20 (.A(a_i[27]),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_2 input21 (.A(a_i[28]),
    .X(net21));
 sky130_fd_sc_hd__buf_1 input22 (.A(a_i[29]),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_2 input23 (.A(a_i[2]),
    .X(net23));
 sky130_fd_sc_hd__buf_1 input24 (.A(a_i[30]),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_1 input25 (.A(a_i[31]),
    .X(net25));
 sky130_fd_sc_hd__buf_1 input26 (.A(a_i[3]),
    .X(net26));
 sky130_fd_sc_hd__buf_1 input27 (.A(a_i[4]),
    .X(net27));
 sky130_fd_sc_hd__buf_1 input28 (.A(a_i[5]),
    .X(net28));
 sky130_fd_sc_hd__buf_1 input29 (.A(a_i[6]),
    .X(net29));
 sky130_fd_sc_hd__clkbuf_4 input3 (.A(a_i[11]),
    .X(net3));
 sky130_fd_sc_hd__buf_1 input30 (.A(a_i[7]),
    .X(net30));
 sky130_fd_sc_hd__buf_1 input31 (.A(a_i[8]),
    .X(net31));
 sky130_fd_sc_hd__clkbuf_1 input32 (.A(a_i[9]),
    .X(net32));
 sky130_fd_sc_hd__clkbuf_2 input33 (.A(b_i[0]),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_1 input34 (.A(b_i[10]),
    .X(net34));
 sky130_fd_sc_hd__clkbuf_4 input35 (.A(b_i[11]),
    .X(net35));
 sky130_fd_sc_hd__clkbuf_4 input36 (.A(b_i[12]),
    .X(net36));
 sky130_fd_sc_hd__clkbuf_4 input37 (.A(b_i[13]),
    .X(net37));
 sky130_fd_sc_hd__buf_2 input38 (.A(b_i[14]),
    .X(net38));
 sky130_fd_sc_hd__clkbuf_2 input39 (.A(b_i[15]),
    .X(net39));
 sky130_fd_sc_hd__buf_2 input4 (.A(a_i[12]),
    .X(net4));
 sky130_fd_sc_hd__buf_2 input40 (.A(b_i[16]),
    .X(net40));
 sky130_fd_sc_hd__clkbuf_1 input41 (.A(b_i[17]),
    .X(net41));
 sky130_fd_sc_hd__buf_1 input42 (.A(b_i[18]),
    .X(net42));
 sky130_fd_sc_hd__clkbuf_2 input43 (.A(b_i[19]),
    .X(net43));
 sky130_fd_sc_hd__buf_4 input44 (.A(b_i[1]),
    .X(net44));
 sky130_fd_sc_hd__buf_1 input45 (.A(b_i[20]),
    .X(net45));
 sky130_fd_sc_hd__buf_4 input46 (.A(b_i[21]),
    .X(net46));
 sky130_fd_sc_hd__buf_1 input47 (.A(b_i[22]),
    .X(net47));
 sky130_fd_sc_hd__buf_1 input48 (.A(b_i[23]),
    .X(net48));
 sky130_fd_sc_hd__buf_4 input49 (.A(b_i[24]),
    .X(net49));
 sky130_fd_sc_hd__buf_4 input5 (.A(a_i[13]),
    .X(net5));
 sky130_fd_sc_hd__buf_4 input50 (.A(b_i[25]),
    .X(net50));
 sky130_fd_sc_hd__clkbuf_4 input51 (.A(b_i[26]),
    .X(net51));
 sky130_fd_sc_hd__clkbuf_4 input52 (.A(b_i[27]),
    .X(net52));
 sky130_fd_sc_hd__clkbuf_4 input53 (.A(b_i[28]),
    .X(net53));
 sky130_fd_sc_hd__buf_2 input54 (.A(b_i[29]),
    .X(net54));
 sky130_fd_sc_hd__clkbuf_4 input55 (.A(b_i[2]),
    .X(net55));
 sky130_fd_sc_hd__clkbuf_2 input56 (.A(b_i[30]),
    .X(net56));
 sky130_fd_sc_hd__dlymetal6s2s_1 input57 (.A(b_i[31]),
    .X(net57));
 sky130_fd_sc_hd__buf_1 input58 (.A(b_i[3]),
    .X(net58));
 sky130_fd_sc_hd__buf_1 input59 (.A(b_i[4]),
    .X(net59));
 sky130_fd_sc_hd__clkbuf_4 input6 (.A(a_i[14]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_1 input60 (.A(b_i[5]),
    .X(net60));
 sky130_fd_sc_hd__clkbuf_1 input61 (.A(b_i[6]),
    .X(net61));
 sky130_fd_sc_hd__clkbuf_1 input62 (.A(b_i[7]),
    .X(net62));
 sky130_fd_sc_hd__buf_1 input63 (.A(b_i[8]),
    .X(net63));
 sky130_fd_sc_hd__buf_1 input64 (.A(b_i[9]),
    .X(net64));
 sky130_fd_sc_hd__clkbuf_2 input65 (.A(nrst),
    .X(net65));
 sky130_fd_sc_hd__clkbuf_2 input7 (.A(a_i[15]),
    .X(net7));
 sky130_fd_sc_hd__buf_2 input8 (.A(a_i[16]),
    .X(net8));
 sky130_fd_sc_hd__dlymetal6s2s_1 input9 (.A(a_i[17]),
    .X(net9));
 sky130_fd_sc_hd__buf_12 output66 (.A(net66),
    .X(y_o[0]));
 sky130_fd_sc_hd__buf_12 output67 (.A(net67),
    .X(y_o[10]));
 sky130_fd_sc_hd__buf_12 output68 (.A(net68),
    .X(y_o[11]));
 sky130_fd_sc_hd__buf_12 output69 (.A(net69),
    .X(y_o[12]));
 sky130_fd_sc_hd__buf_12 output70 (.A(net70),
    .X(y_o[13]));
 sky130_fd_sc_hd__buf_12 output71 (.A(net71),
    .X(y_o[14]));
 sky130_fd_sc_hd__buf_12 output72 (.A(net72),
    .X(y_o[15]));
 sky130_fd_sc_hd__buf_12 output73 (.A(net73),
    .X(y_o[16]));
 sky130_fd_sc_hd__buf_12 output74 (.A(net74),
    .X(y_o[17]));
 sky130_fd_sc_hd__buf_12 output75 (.A(net75),
    .X(y_o[18]));
 sky130_fd_sc_hd__buf_12 output76 (.A(net76),
    .X(y_o[19]));
 sky130_fd_sc_hd__buf_12 output77 (.A(net77),
    .X(y_o[1]));
 sky130_fd_sc_hd__buf_12 output78 (.A(net78),
    .X(y_o[20]));
 sky130_fd_sc_hd__buf_12 output79 (.A(net79),
    .X(y_o[21]));
 sky130_fd_sc_hd__buf_12 output80 (.A(net80),
    .X(y_o[22]));
 sky130_fd_sc_hd__buf_12 output81 (.A(net81),
    .X(y_o[23]));
 sky130_fd_sc_hd__buf_12 output82 (.A(net82),
    .X(y_o[24]));
 sky130_fd_sc_hd__buf_12 output83 (.A(net83),
    .X(y_o[25]));
 sky130_fd_sc_hd__buf_12 output84 (.A(net84),
    .X(y_o[26]));
 sky130_fd_sc_hd__buf_12 output85 (.A(net85),
    .X(y_o[27]));
 sky130_fd_sc_hd__buf_12 output86 (.A(net86),
    .X(y_o[28]));
 sky130_fd_sc_hd__buf_12 output87 (.A(net87),
    .X(y_o[29]));
 sky130_fd_sc_hd__buf_12 output88 (.A(net88),
    .X(y_o[2]));
 sky130_fd_sc_hd__buf_12 output89 (.A(net89),
    .X(y_o[30]));
 sky130_fd_sc_hd__buf_12 output90 (.A(net90),
    .X(y_o[31]));
 sky130_fd_sc_hd__buf_12 output91 (.A(net91),
    .X(y_o[3]));
 sky130_fd_sc_hd__buf_12 output92 (.A(net92),
    .X(y_o[4]));
 sky130_fd_sc_hd__buf_12 output93 (.A(net93),
    .X(y_o[5]));
 sky130_fd_sc_hd__buf_12 output94 (.A(net94),
    .X(y_o[6]));
 sky130_fd_sc_hd__buf_12 output95 (.A(net95),
    .X(y_o[7]));
 sky130_fd_sc_hd__buf_12 output96 (.A(net96),
    .X(y_o[8]));
 sky130_fd_sc_hd__buf_12 output97 (.A(net97),
    .X(y_o[9]));
endmodule

