magic
tech sky130A
magscale 1 2
timestamp 1763328624
<< obsli1 >>
rect 1104 2159 48852 47345
<< obsm1 >>
rect 934 1708 49022 47376
<< metal2 >>
rect 12438 0 12494 800
rect 37370 0 37426 800
<< obsm2 >>
rect 938 856 49018 47365
rect 938 800 12382 856
rect 12550 800 37314 856
rect 37482 800 49018 856
<< metal3 >>
rect 0 45976 800 46096
rect 0 44616 800 44736
rect 0 43256 800 43376
rect 0 41896 800 42016
rect 49200 41896 50000 42016
rect 49200 41352 50000 41472
rect 49200 40808 50000 40928
rect 0 40536 800 40656
rect 49200 40264 50000 40384
rect 49200 39720 50000 39840
rect 0 39176 800 39296
rect 49200 39176 50000 39296
rect 49200 38632 50000 38752
rect 49200 38088 50000 38208
rect 0 37816 800 37936
rect 49200 37544 50000 37664
rect 49200 37000 50000 37120
rect 0 36456 800 36576
rect 49200 36456 50000 36576
rect 49200 35912 50000 36032
rect 49200 35368 50000 35488
rect 0 35096 800 35216
rect 49200 34824 50000 34944
rect 49200 34280 50000 34400
rect 0 33736 800 33856
rect 49200 33736 50000 33856
rect 49200 33192 50000 33312
rect 49200 32648 50000 32768
rect 0 32376 800 32496
rect 49200 32104 50000 32224
rect 49200 31560 50000 31680
rect 0 31016 800 31136
rect 49200 31016 50000 31136
rect 49200 30472 50000 30592
rect 49200 29928 50000 30048
rect 0 29656 800 29776
rect 49200 29384 50000 29504
rect 49200 28840 50000 28960
rect 0 28296 800 28416
rect 49200 28296 50000 28416
rect 49200 27752 50000 27872
rect 49200 27208 50000 27328
rect 0 26936 800 27056
rect 49200 26664 50000 26784
rect 49200 26120 50000 26240
rect 0 25576 800 25696
rect 49200 25576 50000 25696
rect 49200 25032 50000 25152
rect 49200 24488 50000 24608
rect 0 24216 800 24336
rect 49200 23944 50000 24064
rect 49200 23400 50000 23520
rect 0 22856 800 22976
rect 49200 22856 50000 22976
rect 49200 22312 50000 22432
rect 49200 21768 50000 21888
rect 0 21496 800 21616
rect 49200 21224 50000 21344
rect 49200 20680 50000 20800
rect 0 20136 800 20256
rect 49200 20136 50000 20256
rect 49200 19592 50000 19712
rect 49200 19048 50000 19168
rect 0 18776 800 18896
rect 49200 18504 50000 18624
rect 49200 17960 50000 18080
rect 0 17416 800 17536
rect 49200 17416 50000 17536
rect 49200 16872 50000 16992
rect 49200 16328 50000 16448
rect 0 16056 800 16176
rect 49200 15784 50000 15904
rect 49200 15240 50000 15360
rect 0 14696 800 14816
rect 49200 14696 50000 14816
rect 49200 14152 50000 14272
rect 49200 13608 50000 13728
rect 0 13336 800 13456
rect 49200 13064 50000 13184
rect 49200 12520 50000 12640
rect 0 11976 800 12096
rect 49200 11976 50000 12096
rect 49200 11432 50000 11552
rect 49200 10888 50000 11008
rect 0 10616 800 10736
rect 49200 10344 50000 10464
rect 49200 9800 50000 9920
rect 0 9256 800 9376
rect 49200 9256 50000 9376
rect 49200 8712 50000 8832
rect 49200 8168 50000 8288
rect 0 7896 800 8016
rect 49200 7624 50000 7744
rect 0 6536 800 6656
rect 0 5176 800 5296
rect 0 3816 800 3936
<< obsm3 >>
rect 798 46176 49200 47361
rect 880 45896 49200 46176
rect 798 44816 49200 45896
rect 880 44536 49200 44816
rect 798 43456 49200 44536
rect 880 43176 49200 43456
rect 798 42096 49200 43176
rect 880 41816 49120 42096
rect 798 41552 49200 41816
rect 798 41272 49120 41552
rect 798 41008 49200 41272
rect 798 40736 49120 41008
rect 880 40728 49120 40736
rect 880 40464 49200 40728
rect 880 40456 49120 40464
rect 798 40184 49120 40456
rect 798 39920 49200 40184
rect 798 39640 49120 39920
rect 798 39376 49200 39640
rect 880 39096 49120 39376
rect 798 38832 49200 39096
rect 798 38552 49120 38832
rect 798 38288 49200 38552
rect 798 38016 49120 38288
rect 880 38008 49120 38016
rect 880 37744 49200 38008
rect 880 37736 49120 37744
rect 798 37464 49120 37736
rect 798 37200 49200 37464
rect 798 36920 49120 37200
rect 798 36656 49200 36920
rect 880 36376 49120 36656
rect 798 36112 49200 36376
rect 798 35832 49120 36112
rect 798 35568 49200 35832
rect 798 35296 49120 35568
rect 880 35288 49120 35296
rect 880 35024 49200 35288
rect 880 35016 49120 35024
rect 798 34744 49120 35016
rect 798 34480 49200 34744
rect 798 34200 49120 34480
rect 798 33936 49200 34200
rect 880 33656 49120 33936
rect 798 33392 49200 33656
rect 798 33112 49120 33392
rect 798 32848 49200 33112
rect 798 32576 49120 32848
rect 880 32568 49120 32576
rect 880 32304 49200 32568
rect 880 32296 49120 32304
rect 798 32024 49120 32296
rect 798 31760 49200 32024
rect 798 31480 49120 31760
rect 798 31216 49200 31480
rect 880 30936 49120 31216
rect 798 30672 49200 30936
rect 798 30392 49120 30672
rect 798 30128 49200 30392
rect 798 29856 49120 30128
rect 880 29848 49120 29856
rect 880 29584 49200 29848
rect 880 29576 49120 29584
rect 798 29304 49120 29576
rect 798 29040 49200 29304
rect 798 28760 49120 29040
rect 798 28496 49200 28760
rect 880 28216 49120 28496
rect 798 27952 49200 28216
rect 798 27672 49120 27952
rect 798 27408 49200 27672
rect 798 27136 49120 27408
rect 880 27128 49120 27136
rect 880 26864 49200 27128
rect 880 26856 49120 26864
rect 798 26584 49120 26856
rect 798 26320 49200 26584
rect 798 26040 49120 26320
rect 798 25776 49200 26040
rect 880 25496 49120 25776
rect 798 25232 49200 25496
rect 798 24952 49120 25232
rect 798 24688 49200 24952
rect 798 24416 49120 24688
rect 880 24408 49120 24416
rect 880 24144 49200 24408
rect 880 24136 49120 24144
rect 798 23864 49120 24136
rect 798 23600 49200 23864
rect 798 23320 49120 23600
rect 798 23056 49200 23320
rect 880 22776 49120 23056
rect 798 22512 49200 22776
rect 798 22232 49120 22512
rect 798 21968 49200 22232
rect 798 21696 49120 21968
rect 880 21688 49120 21696
rect 880 21424 49200 21688
rect 880 21416 49120 21424
rect 798 21144 49120 21416
rect 798 20880 49200 21144
rect 798 20600 49120 20880
rect 798 20336 49200 20600
rect 880 20056 49120 20336
rect 798 19792 49200 20056
rect 798 19512 49120 19792
rect 798 19248 49200 19512
rect 798 18976 49120 19248
rect 880 18968 49120 18976
rect 880 18704 49200 18968
rect 880 18696 49120 18704
rect 798 18424 49120 18696
rect 798 18160 49200 18424
rect 798 17880 49120 18160
rect 798 17616 49200 17880
rect 880 17336 49120 17616
rect 798 17072 49200 17336
rect 798 16792 49120 17072
rect 798 16528 49200 16792
rect 798 16256 49120 16528
rect 880 16248 49120 16256
rect 880 15984 49200 16248
rect 880 15976 49120 15984
rect 798 15704 49120 15976
rect 798 15440 49200 15704
rect 798 15160 49120 15440
rect 798 14896 49200 15160
rect 880 14616 49120 14896
rect 798 14352 49200 14616
rect 798 14072 49120 14352
rect 798 13808 49200 14072
rect 798 13536 49120 13808
rect 880 13528 49120 13536
rect 880 13264 49200 13528
rect 880 13256 49120 13264
rect 798 12984 49120 13256
rect 798 12720 49200 12984
rect 798 12440 49120 12720
rect 798 12176 49200 12440
rect 880 11896 49120 12176
rect 798 11632 49200 11896
rect 798 11352 49120 11632
rect 798 11088 49200 11352
rect 798 10816 49120 11088
rect 880 10808 49120 10816
rect 880 10544 49200 10808
rect 880 10536 49120 10544
rect 798 10264 49120 10536
rect 798 10000 49200 10264
rect 798 9720 49120 10000
rect 798 9456 49200 9720
rect 880 9176 49120 9456
rect 798 8912 49200 9176
rect 798 8632 49120 8912
rect 798 8368 49200 8632
rect 798 8096 49120 8368
rect 880 8088 49120 8096
rect 880 7824 49200 8088
rect 880 7816 49120 7824
rect 798 7544 49120 7816
rect 798 6736 49200 7544
rect 880 6456 49200 6736
rect 798 5376 49200 6456
rect 880 5096 49200 5376
rect 798 4016 49200 5096
rect 880 3736 49200 4016
rect 798 2143 49200 3736
<< metal4 >>
rect 4208 2128 4528 47376
rect 19568 2128 19888 47376
rect 34928 2128 35248 47376
<< obsm4 >>
rect 3923 3843 4128 45661
rect 4608 3843 19488 45661
rect 19968 3843 34848 45661
rect 35328 3843 48149 45661
<< labels >>
rlabel metal3 s 49200 7624 50000 7744 6 a_i[0]
port 1 nsew signal input
rlabel metal3 s 49200 13064 50000 13184 6 a_i[10]
port 2 nsew signal input
rlabel metal3 s 49200 13608 50000 13728 6 a_i[11]
port 3 nsew signal input
rlabel metal3 s 49200 14152 50000 14272 6 a_i[12]
port 4 nsew signal input
rlabel metal3 s 49200 14696 50000 14816 6 a_i[13]
port 5 nsew signal input
rlabel metal3 s 49200 15240 50000 15360 6 a_i[14]
port 6 nsew signal input
rlabel metal3 s 49200 15784 50000 15904 6 a_i[15]
port 7 nsew signal input
rlabel metal3 s 49200 16328 50000 16448 6 a_i[16]
port 8 nsew signal input
rlabel metal3 s 49200 16872 50000 16992 6 a_i[17]
port 9 nsew signal input
rlabel metal3 s 49200 17416 50000 17536 6 a_i[18]
port 10 nsew signal input
rlabel metal3 s 49200 17960 50000 18080 6 a_i[19]
port 11 nsew signal input
rlabel metal3 s 49200 8168 50000 8288 6 a_i[1]
port 12 nsew signal input
rlabel metal3 s 49200 18504 50000 18624 6 a_i[20]
port 13 nsew signal input
rlabel metal3 s 49200 19048 50000 19168 6 a_i[21]
port 14 nsew signal input
rlabel metal3 s 49200 19592 50000 19712 6 a_i[22]
port 15 nsew signal input
rlabel metal3 s 49200 20136 50000 20256 6 a_i[23]
port 16 nsew signal input
rlabel metal3 s 49200 20680 50000 20800 6 a_i[24]
port 17 nsew signal input
rlabel metal3 s 49200 21224 50000 21344 6 a_i[25]
port 18 nsew signal input
rlabel metal3 s 49200 21768 50000 21888 6 a_i[26]
port 19 nsew signal input
rlabel metal3 s 49200 22312 50000 22432 6 a_i[27]
port 20 nsew signal input
rlabel metal3 s 49200 22856 50000 22976 6 a_i[28]
port 21 nsew signal input
rlabel metal3 s 49200 23400 50000 23520 6 a_i[29]
port 22 nsew signal input
rlabel metal3 s 49200 8712 50000 8832 6 a_i[2]
port 23 nsew signal input
rlabel metal3 s 49200 23944 50000 24064 6 a_i[30]
port 24 nsew signal input
rlabel metal3 s 49200 24488 50000 24608 6 a_i[31]
port 25 nsew signal input
rlabel metal3 s 49200 9256 50000 9376 6 a_i[3]
port 26 nsew signal input
rlabel metal3 s 49200 9800 50000 9920 6 a_i[4]
port 27 nsew signal input
rlabel metal3 s 49200 10344 50000 10464 6 a_i[5]
port 28 nsew signal input
rlabel metal3 s 49200 10888 50000 11008 6 a_i[6]
port 29 nsew signal input
rlabel metal3 s 49200 11432 50000 11552 6 a_i[7]
port 30 nsew signal input
rlabel metal3 s 49200 11976 50000 12096 6 a_i[8]
port 31 nsew signal input
rlabel metal3 s 49200 12520 50000 12640 6 a_i[9]
port 32 nsew signal input
rlabel metal3 s 49200 25032 50000 25152 6 b_i[0]
port 33 nsew signal input
rlabel metal3 s 49200 30472 50000 30592 6 b_i[10]
port 34 nsew signal input
rlabel metal3 s 49200 31016 50000 31136 6 b_i[11]
port 35 nsew signal input
rlabel metal3 s 49200 31560 50000 31680 6 b_i[12]
port 36 nsew signal input
rlabel metal3 s 49200 32104 50000 32224 6 b_i[13]
port 37 nsew signal input
rlabel metal3 s 49200 32648 50000 32768 6 b_i[14]
port 38 nsew signal input
rlabel metal3 s 49200 33192 50000 33312 6 b_i[15]
port 39 nsew signal input
rlabel metal3 s 49200 33736 50000 33856 6 b_i[16]
port 40 nsew signal input
rlabel metal3 s 49200 34280 50000 34400 6 b_i[17]
port 41 nsew signal input
rlabel metal3 s 49200 34824 50000 34944 6 b_i[18]
port 42 nsew signal input
rlabel metal3 s 49200 35368 50000 35488 6 b_i[19]
port 43 nsew signal input
rlabel metal3 s 49200 25576 50000 25696 6 b_i[1]
port 44 nsew signal input
rlabel metal3 s 49200 35912 50000 36032 6 b_i[20]
port 45 nsew signal input
rlabel metal3 s 49200 36456 50000 36576 6 b_i[21]
port 46 nsew signal input
rlabel metal3 s 49200 37000 50000 37120 6 b_i[22]
port 47 nsew signal input
rlabel metal3 s 49200 37544 50000 37664 6 b_i[23]
port 48 nsew signal input
rlabel metal3 s 49200 38088 50000 38208 6 b_i[24]
port 49 nsew signal input
rlabel metal3 s 49200 38632 50000 38752 6 b_i[25]
port 50 nsew signal input
rlabel metal3 s 49200 39176 50000 39296 6 b_i[26]
port 51 nsew signal input
rlabel metal3 s 49200 39720 50000 39840 6 b_i[27]
port 52 nsew signal input
rlabel metal3 s 49200 40264 50000 40384 6 b_i[28]
port 53 nsew signal input
rlabel metal3 s 49200 40808 50000 40928 6 b_i[29]
port 54 nsew signal input
rlabel metal3 s 49200 26120 50000 26240 6 b_i[2]
port 55 nsew signal input
rlabel metal3 s 49200 41352 50000 41472 6 b_i[30]
port 56 nsew signal input
rlabel metal3 s 49200 41896 50000 42016 6 b_i[31]
port 57 nsew signal input
rlabel metal3 s 49200 26664 50000 26784 6 b_i[3]
port 58 nsew signal input
rlabel metal3 s 49200 27208 50000 27328 6 b_i[4]
port 59 nsew signal input
rlabel metal3 s 49200 27752 50000 27872 6 b_i[5]
port 60 nsew signal input
rlabel metal3 s 49200 28296 50000 28416 6 b_i[6]
port 61 nsew signal input
rlabel metal3 s 49200 28840 50000 28960 6 b_i[7]
port 62 nsew signal input
rlabel metal3 s 49200 29384 50000 29504 6 b_i[8]
port 63 nsew signal input
rlabel metal3 s 49200 29928 50000 30048 6 b_i[9]
port 64 nsew signal input
rlabel metal2 s 12438 0 12494 800 6 clk
port 65 nsew signal input
rlabel metal2 s 37370 0 37426 800 6 nrst
port 66 nsew signal input
rlabel metal4 s 4208 2128 4528 47376 6 vccd1
port 67 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 47376 6 vccd1
port 67 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 47376 6 vssd1
port 68 nsew ground bidirectional
rlabel metal3 s 0 3816 800 3936 6 y_o[0]
port 69 nsew signal output
rlabel metal3 s 0 17416 800 17536 6 y_o[10]
port 70 nsew signal output
rlabel metal3 s 0 18776 800 18896 6 y_o[11]
port 71 nsew signal output
rlabel metal3 s 0 20136 800 20256 6 y_o[12]
port 72 nsew signal output
rlabel metal3 s 0 21496 800 21616 6 y_o[13]
port 73 nsew signal output
rlabel metal3 s 0 22856 800 22976 6 y_o[14]
port 74 nsew signal output
rlabel metal3 s 0 24216 800 24336 6 y_o[15]
port 75 nsew signal output
rlabel metal3 s 0 25576 800 25696 6 y_o[16]
port 76 nsew signal output
rlabel metal3 s 0 26936 800 27056 6 y_o[17]
port 77 nsew signal output
rlabel metal3 s 0 28296 800 28416 6 y_o[18]
port 78 nsew signal output
rlabel metal3 s 0 29656 800 29776 6 y_o[19]
port 79 nsew signal output
rlabel metal3 s 0 5176 800 5296 6 y_o[1]
port 80 nsew signal output
rlabel metal3 s 0 31016 800 31136 6 y_o[20]
port 81 nsew signal output
rlabel metal3 s 0 32376 800 32496 6 y_o[21]
port 82 nsew signal output
rlabel metal3 s 0 33736 800 33856 6 y_o[22]
port 83 nsew signal output
rlabel metal3 s 0 35096 800 35216 6 y_o[23]
port 84 nsew signal output
rlabel metal3 s 0 36456 800 36576 6 y_o[24]
port 85 nsew signal output
rlabel metal3 s 0 37816 800 37936 6 y_o[25]
port 86 nsew signal output
rlabel metal3 s 0 39176 800 39296 6 y_o[26]
port 87 nsew signal output
rlabel metal3 s 0 40536 800 40656 6 y_o[27]
port 88 nsew signal output
rlabel metal3 s 0 41896 800 42016 6 y_o[28]
port 89 nsew signal output
rlabel metal3 s 0 43256 800 43376 6 y_o[29]
port 90 nsew signal output
rlabel metal3 s 0 6536 800 6656 6 y_o[2]
port 91 nsew signal output
rlabel metal3 s 0 44616 800 44736 6 y_o[30]
port 92 nsew signal output
rlabel metal3 s 0 45976 800 46096 6 y_o[31]
port 93 nsew signal output
rlabel metal3 s 0 7896 800 8016 6 y_o[3]
port 94 nsew signal output
rlabel metal3 s 0 9256 800 9376 6 y_o[4]
port 95 nsew signal output
rlabel metal3 s 0 10616 800 10736 6 y_o[5]
port 96 nsew signal output
rlabel metal3 s 0 11976 800 12096 6 y_o[6]
port 97 nsew signal output
rlabel metal3 s 0 13336 800 13456 6 y_o[7]
port 98 nsew signal output
rlabel metal3 s 0 14696 800 14816 6 y_o[8]
port 99 nsew signal output
rlabel metal3 s 0 16056 800 16176 6 y_o[9]
port 100 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 50000 50000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 11131228
string GDS_FILE /home/sforde22/Caravel/sdmay26-24/openlane/mac/runs/25_11_16_15_25/results/signoff/mac.magic.gds
string GDS_START 431116
<< end >>

