VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO mac_piped
  CLASS BLOCK ;
  FOREIGN mac_piped ;
  ORIGIN 0.000 0.000 ;
  SIZE 300.000 BY 300.000 ;
  PIN a_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 296.000 20.440 300.000 21.040 ;
    END
  END a_i[0]
  PIN a_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 61.240 300.000 61.840 ;
    END
  END a_i[10]
  PIN a_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 296.000 65.320 300.000 65.920 ;
    END
  END a_i[11]
  PIN a_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 296.000 69.400 300.000 70.000 ;
    END
  END a_i[12]
  PIN a_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 73.480 300.000 74.080 ;
    END
  END a_i[13]
  PIN a_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 296.000 77.560 300.000 78.160 ;
    END
  END a_i[14]
  PIN a_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 296.000 81.640 300.000 82.240 ;
    END
  END a_i[15]
  PIN a_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 296.000 85.720 300.000 86.320 ;
    END
  END a_i[16]
  PIN a_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 296.000 89.800 300.000 90.400 ;
    END
  END a_i[17]
  PIN a_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 93.880 300.000 94.480 ;
    END
  END a_i[18]
  PIN a_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 97.960 300.000 98.560 ;
    END
  END a_i[19]
  PIN a_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 296.000 24.520 300.000 25.120 ;
    END
  END a_i[1]
  PIN a_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 102.040 300.000 102.640 ;
    END
  END a_i[20]
  PIN a_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 106.120 300.000 106.720 ;
    END
  END a_i[21]
  PIN a_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 110.200 300.000 110.800 ;
    END
  END a_i[22]
  PIN a_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 114.280 300.000 114.880 ;
    END
  END a_i[23]
  PIN a_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 296.000 118.360 300.000 118.960 ;
    END
  END a_i[24]
  PIN a_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 296.000 122.440 300.000 123.040 ;
    END
  END a_i[25]
  PIN a_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 296.000 126.520 300.000 127.120 ;
    END
  END a_i[26]
  PIN a_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 296.000 130.600 300.000 131.200 ;
    END
  END a_i[27]
  PIN a_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 296.000 134.680 300.000 135.280 ;
    END
  END a_i[28]
  PIN a_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 138.760 300.000 139.360 ;
    END
  END a_i[29]
  PIN a_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 296.000 28.600 300.000 29.200 ;
    END
  END a_i[2]
  PIN a_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 142.840 300.000 143.440 ;
    END
  END a_i[30]
  PIN a_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 146.920 300.000 147.520 ;
    END
  END a_i[31]
  PIN a_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 32.680 300.000 33.280 ;
    END
  END a_i[3]
  PIN a_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 36.760 300.000 37.360 ;
    END
  END a_i[4]
  PIN a_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 40.840 300.000 41.440 ;
    END
  END a_i[5]
  PIN a_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 44.920 300.000 45.520 ;
    END
  END a_i[6]
  PIN a_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 49.000 300.000 49.600 ;
    END
  END a_i[7]
  PIN a_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 53.080 300.000 53.680 ;
    END
  END a_i[8]
  PIN a_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 57.160 300.000 57.760 ;
    END
  END a_i[9]
  PIN b_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 296.000 151.000 300.000 151.600 ;
    END
  END b_i[0]
  PIN b_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 191.800 300.000 192.400 ;
    END
  END b_i[10]
  PIN b_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 296.000 195.880 300.000 196.480 ;
    END
  END b_i[11]
  PIN b_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 296.000 199.960 300.000 200.560 ;
    END
  END b_i[12]
  PIN b_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 296.000 204.040 300.000 204.640 ;
    END
  END b_i[13]
  PIN b_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 296.000 208.120 300.000 208.720 ;
    END
  END b_i[14]
  PIN b_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 296.000 212.200 300.000 212.800 ;
    END
  END b_i[15]
  PIN b_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 296.000 216.280 300.000 216.880 ;
    END
  END b_i[16]
  PIN b_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 220.360 300.000 220.960 ;
    END
  END b_i[17]
  PIN b_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 224.440 300.000 225.040 ;
    END
  END b_i[18]
  PIN b_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 296.000 228.520 300.000 229.120 ;
    END
  END b_i[19]
  PIN b_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 155.080 300.000 155.680 ;
    END
  END b_i[1]
  PIN b_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 232.600 300.000 233.200 ;
    END
  END b_i[20]
  PIN b_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 236.680 300.000 237.280 ;
    END
  END b_i[21]
  PIN b_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 240.760 300.000 241.360 ;
    END
  END b_i[22]
  PIN b_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 244.840 300.000 245.440 ;
    END
  END b_i[23]
  PIN b_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 248.920 300.000 249.520 ;
    END
  END b_i[24]
  PIN b_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 253.000 300.000 253.600 ;
    END
  END b_i[25]
  PIN b_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 296.000 257.080 300.000 257.680 ;
    END
  END b_i[26]
  PIN b_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 296.000 261.160 300.000 261.760 ;
    END
  END b_i[27]
  PIN b_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 296.000 265.240 300.000 265.840 ;
    END
  END b_i[28]
  PIN b_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 296.000 269.320 300.000 269.920 ;
    END
  END b_i[29]
  PIN b_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 296.000 159.160 300.000 159.760 ;
    END
  END b_i[2]
  PIN b_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 296.000 273.400 300.000 274.000 ;
    END
  END b_i[30]
  PIN b_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 296.000 277.480 300.000 278.080 ;
    END
  END b_i[31]
  PIN b_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 163.240 300.000 163.840 ;
    END
  END b_i[3]
  PIN b_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 167.320 300.000 167.920 ;
    END
  END b_i[4]
  PIN b_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 171.400 300.000 172.000 ;
    END
  END b_i[5]
  PIN b_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 175.480 300.000 176.080 ;
    END
  END b_i[6]
  PIN b_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 179.560 300.000 180.160 ;
    END
  END b_i[7]
  PIN b_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 183.640 300.000 184.240 ;
    END
  END b_i[8]
  PIN b_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 187.720 300.000 188.320 ;
    END
  END b_i[9]
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met2 ;
        RECT 74.610 0.000 74.890 4.000 ;
    END
  END clk
  PIN nrst
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 224.570 0.000 224.850 4.000 ;
    END
  END nrst
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 288.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 288.560 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 288.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 288.560 ;
    END
  END vssd1
  PIN y_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 23.160 4.000 23.760 ;
    END
  END y_o[0]
  PIN y_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 104.760 4.000 105.360 ;
    END
  END y_o[10]
  PIN y_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 112.920 4.000 113.520 ;
    END
  END y_o[11]
  PIN y_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 121.080 4.000 121.680 ;
    END
  END y_o[12]
  PIN y_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 129.240 4.000 129.840 ;
    END
  END y_o[13]
  PIN y_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 137.400 4.000 138.000 ;
    END
  END y_o[14]
  PIN y_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 145.560 4.000 146.160 ;
    END
  END y_o[15]
  PIN y_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 153.720 4.000 154.320 ;
    END
  END y_o[16]
  PIN y_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 161.880 4.000 162.480 ;
    END
  END y_o[17]
  PIN y_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 170.040 4.000 170.640 ;
    END
  END y_o[18]
  PIN y_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 178.200 4.000 178.800 ;
    END
  END y_o[19]
  PIN y_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 31.320 4.000 31.920 ;
    END
  END y_o[1]
  PIN y_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 186.360 4.000 186.960 ;
    END
  END y_o[20]
  PIN y_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 194.520 4.000 195.120 ;
    END
  END y_o[21]
  PIN y_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 202.680 4.000 203.280 ;
    END
  END y_o[22]
  PIN y_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 210.840 4.000 211.440 ;
    END
  END y_o[23]
  PIN y_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 219.000 4.000 219.600 ;
    END
  END y_o[24]
  PIN y_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 227.160 4.000 227.760 ;
    END
  END y_o[25]
  PIN y_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 235.320 4.000 235.920 ;
    END
  END y_o[26]
  PIN y_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 243.480 4.000 244.080 ;
    END
  END y_o[27]
  PIN y_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 251.640 4.000 252.240 ;
    END
  END y_o[28]
  PIN y_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 259.800 4.000 260.400 ;
    END
  END y_o[29]
  PIN y_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 39.480 4.000 40.080 ;
    END
  END y_o[2]
  PIN y_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 267.960 4.000 268.560 ;
    END
  END y_o[30]
  PIN y_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 276.120 4.000 276.720 ;
    END
  END y_o[31]
  PIN y_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 47.640 4.000 48.240 ;
    END
  END y_o[3]
  PIN y_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 55.800 4.000 56.400 ;
    END
  END y_o[4]
  PIN y_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 63.960 4.000 64.560 ;
    END
  END y_o[5]
  PIN y_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 72.120 4.000 72.720 ;
    END
  END y_o[6]
  PIN y_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 80.280 4.000 80.880 ;
    END
  END y_o[7]
  PIN y_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 88.440 4.000 89.040 ;
    END
  END y_o[8]
  PIN y_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 96.600 4.000 97.200 ;
    END
  END y_o[9]
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 294.400 288.405 ;
      LAYER met1 ;
        RECT 4.670 10.640 298.930 288.560 ;
      LAYER met2 ;
        RECT 4.690 4.280 298.900 288.505 ;
        RECT 4.690 4.000 74.330 4.280 ;
        RECT 75.170 4.000 224.290 4.280 ;
        RECT 225.130 4.000 298.900 4.280 ;
      LAYER met3 ;
        RECT 3.990 278.480 296.000 288.485 ;
        RECT 3.990 277.120 295.600 278.480 ;
        RECT 4.400 277.080 295.600 277.120 ;
        RECT 4.400 275.720 296.000 277.080 ;
        RECT 3.990 274.400 296.000 275.720 ;
        RECT 3.990 273.000 295.600 274.400 ;
        RECT 3.990 270.320 296.000 273.000 ;
        RECT 3.990 268.960 295.600 270.320 ;
        RECT 4.400 268.920 295.600 268.960 ;
        RECT 4.400 267.560 296.000 268.920 ;
        RECT 3.990 266.240 296.000 267.560 ;
        RECT 3.990 264.840 295.600 266.240 ;
        RECT 3.990 262.160 296.000 264.840 ;
        RECT 3.990 260.800 295.600 262.160 ;
        RECT 4.400 260.760 295.600 260.800 ;
        RECT 4.400 259.400 296.000 260.760 ;
        RECT 3.990 258.080 296.000 259.400 ;
        RECT 3.990 256.680 295.600 258.080 ;
        RECT 3.990 254.000 296.000 256.680 ;
        RECT 3.990 252.640 295.600 254.000 ;
        RECT 4.400 252.600 295.600 252.640 ;
        RECT 4.400 251.240 296.000 252.600 ;
        RECT 3.990 249.920 296.000 251.240 ;
        RECT 3.990 248.520 295.600 249.920 ;
        RECT 3.990 245.840 296.000 248.520 ;
        RECT 3.990 244.480 295.600 245.840 ;
        RECT 4.400 244.440 295.600 244.480 ;
        RECT 4.400 243.080 296.000 244.440 ;
        RECT 3.990 241.760 296.000 243.080 ;
        RECT 3.990 240.360 295.600 241.760 ;
        RECT 3.990 237.680 296.000 240.360 ;
        RECT 3.990 236.320 295.600 237.680 ;
        RECT 4.400 236.280 295.600 236.320 ;
        RECT 4.400 234.920 296.000 236.280 ;
        RECT 3.990 233.600 296.000 234.920 ;
        RECT 3.990 232.200 295.600 233.600 ;
        RECT 3.990 229.520 296.000 232.200 ;
        RECT 3.990 228.160 295.600 229.520 ;
        RECT 4.400 228.120 295.600 228.160 ;
        RECT 4.400 226.760 296.000 228.120 ;
        RECT 3.990 225.440 296.000 226.760 ;
        RECT 3.990 224.040 295.600 225.440 ;
        RECT 3.990 221.360 296.000 224.040 ;
        RECT 3.990 220.000 295.600 221.360 ;
        RECT 4.400 219.960 295.600 220.000 ;
        RECT 4.400 218.600 296.000 219.960 ;
        RECT 3.990 217.280 296.000 218.600 ;
        RECT 3.990 215.880 295.600 217.280 ;
        RECT 3.990 213.200 296.000 215.880 ;
        RECT 3.990 211.840 295.600 213.200 ;
        RECT 4.400 211.800 295.600 211.840 ;
        RECT 4.400 210.440 296.000 211.800 ;
        RECT 3.990 209.120 296.000 210.440 ;
        RECT 3.990 207.720 295.600 209.120 ;
        RECT 3.990 205.040 296.000 207.720 ;
        RECT 3.990 203.680 295.600 205.040 ;
        RECT 4.400 203.640 295.600 203.680 ;
        RECT 4.400 202.280 296.000 203.640 ;
        RECT 3.990 200.960 296.000 202.280 ;
        RECT 3.990 199.560 295.600 200.960 ;
        RECT 3.990 196.880 296.000 199.560 ;
        RECT 3.990 195.520 295.600 196.880 ;
        RECT 4.400 195.480 295.600 195.520 ;
        RECT 4.400 194.120 296.000 195.480 ;
        RECT 3.990 192.800 296.000 194.120 ;
        RECT 3.990 191.400 295.600 192.800 ;
        RECT 3.990 188.720 296.000 191.400 ;
        RECT 3.990 187.360 295.600 188.720 ;
        RECT 4.400 187.320 295.600 187.360 ;
        RECT 4.400 185.960 296.000 187.320 ;
        RECT 3.990 184.640 296.000 185.960 ;
        RECT 3.990 183.240 295.600 184.640 ;
        RECT 3.990 180.560 296.000 183.240 ;
        RECT 3.990 179.200 295.600 180.560 ;
        RECT 4.400 179.160 295.600 179.200 ;
        RECT 4.400 177.800 296.000 179.160 ;
        RECT 3.990 176.480 296.000 177.800 ;
        RECT 3.990 175.080 295.600 176.480 ;
        RECT 3.990 172.400 296.000 175.080 ;
        RECT 3.990 171.040 295.600 172.400 ;
        RECT 4.400 171.000 295.600 171.040 ;
        RECT 4.400 169.640 296.000 171.000 ;
        RECT 3.990 168.320 296.000 169.640 ;
        RECT 3.990 166.920 295.600 168.320 ;
        RECT 3.990 164.240 296.000 166.920 ;
        RECT 3.990 162.880 295.600 164.240 ;
        RECT 4.400 162.840 295.600 162.880 ;
        RECT 4.400 161.480 296.000 162.840 ;
        RECT 3.990 160.160 296.000 161.480 ;
        RECT 3.990 158.760 295.600 160.160 ;
        RECT 3.990 156.080 296.000 158.760 ;
        RECT 3.990 154.720 295.600 156.080 ;
        RECT 4.400 154.680 295.600 154.720 ;
        RECT 4.400 153.320 296.000 154.680 ;
        RECT 3.990 152.000 296.000 153.320 ;
        RECT 3.990 150.600 295.600 152.000 ;
        RECT 3.990 147.920 296.000 150.600 ;
        RECT 3.990 146.560 295.600 147.920 ;
        RECT 4.400 146.520 295.600 146.560 ;
        RECT 4.400 145.160 296.000 146.520 ;
        RECT 3.990 143.840 296.000 145.160 ;
        RECT 3.990 142.440 295.600 143.840 ;
        RECT 3.990 139.760 296.000 142.440 ;
        RECT 3.990 138.400 295.600 139.760 ;
        RECT 4.400 138.360 295.600 138.400 ;
        RECT 4.400 137.000 296.000 138.360 ;
        RECT 3.990 135.680 296.000 137.000 ;
        RECT 3.990 134.280 295.600 135.680 ;
        RECT 3.990 131.600 296.000 134.280 ;
        RECT 3.990 130.240 295.600 131.600 ;
        RECT 4.400 130.200 295.600 130.240 ;
        RECT 4.400 128.840 296.000 130.200 ;
        RECT 3.990 127.520 296.000 128.840 ;
        RECT 3.990 126.120 295.600 127.520 ;
        RECT 3.990 123.440 296.000 126.120 ;
        RECT 3.990 122.080 295.600 123.440 ;
        RECT 4.400 122.040 295.600 122.080 ;
        RECT 4.400 120.680 296.000 122.040 ;
        RECT 3.990 119.360 296.000 120.680 ;
        RECT 3.990 117.960 295.600 119.360 ;
        RECT 3.990 115.280 296.000 117.960 ;
        RECT 3.990 113.920 295.600 115.280 ;
        RECT 4.400 113.880 295.600 113.920 ;
        RECT 4.400 112.520 296.000 113.880 ;
        RECT 3.990 111.200 296.000 112.520 ;
        RECT 3.990 109.800 295.600 111.200 ;
        RECT 3.990 107.120 296.000 109.800 ;
        RECT 3.990 105.760 295.600 107.120 ;
        RECT 4.400 105.720 295.600 105.760 ;
        RECT 4.400 104.360 296.000 105.720 ;
        RECT 3.990 103.040 296.000 104.360 ;
        RECT 3.990 101.640 295.600 103.040 ;
        RECT 3.990 98.960 296.000 101.640 ;
        RECT 3.990 97.600 295.600 98.960 ;
        RECT 4.400 97.560 295.600 97.600 ;
        RECT 4.400 96.200 296.000 97.560 ;
        RECT 3.990 94.880 296.000 96.200 ;
        RECT 3.990 93.480 295.600 94.880 ;
        RECT 3.990 90.800 296.000 93.480 ;
        RECT 3.990 89.440 295.600 90.800 ;
        RECT 4.400 89.400 295.600 89.440 ;
        RECT 4.400 88.040 296.000 89.400 ;
        RECT 3.990 86.720 296.000 88.040 ;
        RECT 3.990 85.320 295.600 86.720 ;
        RECT 3.990 82.640 296.000 85.320 ;
        RECT 3.990 81.280 295.600 82.640 ;
        RECT 4.400 81.240 295.600 81.280 ;
        RECT 4.400 79.880 296.000 81.240 ;
        RECT 3.990 78.560 296.000 79.880 ;
        RECT 3.990 77.160 295.600 78.560 ;
        RECT 3.990 74.480 296.000 77.160 ;
        RECT 3.990 73.120 295.600 74.480 ;
        RECT 4.400 73.080 295.600 73.120 ;
        RECT 4.400 71.720 296.000 73.080 ;
        RECT 3.990 70.400 296.000 71.720 ;
        RECT 3.990 69.000 295.600 70.400 ;
        RECT 3.990 66.320 296.000 69.000 ;
        RECT 3.990 64.960 295.600 66.320 ;
        RECT 4.400 64.920 295.600 64.960 ;
        RECT 4.400 63.560 296.000 64.920 ;
        RECT 3.990 62.240 296.000 63.560 ;
        RECT 3.990 60.840 295.600 62.240 ;
        RECT 3.990 58.160 296.000 60.840 ;
        RECT 3.990 56.800 295.600 58.160 ;
        RECT 4.400 56.760 295.600 56.800 ;
        RECT 4.400 55.400 296.000 56.760 ;
        RECT 3.990 54.080 296.000 55.400 ;
        RECT 3.990 52.680 295.600 54.080 ;
        RECT 3.990 50.000 296.000 52.680 ;
        RECT 3.990 48.640 295.600 50.000 ;
        RECT 4.400 48.600 295.600 48.640 ;
        RECT 4.400 47.240 296.000 48.600 ;
        RECT 3.990 45.920 296.000 47.240 ;
        RECT 3.990 44.520 295.600 45.920 ;
        RECT 3.990 41.840 296.000 44.520 ;
        RECT 3.990 40.480 295.600 41.840 ;
        RECT 4.400 40.440 295.600 40.480 ;
        RECT 4.400 39.080 296.000 40.440 ;
        RECT 3.990 37.760 296.000 39.080 ;
        RECT 3.990 36.360 295.600 37.760 ;
        RECT 3.990 33.680 296.000 36.360 ;
        RECT 3.990 32.320 295.600 33.680 ;
        RECT 4.400 32.280 295.600 32.320 ;
        RECT 4.400 30.920 296.000 32.280 ;
        RECT 3.990 29.600 296.000 30.920 ;
        RECT 3.990 28.200 295.600 29.600 ;
        RECT 3.990 25.520 296.000 28.200 ;
        RECT 3.990 24.160 295.600 25.520 ;
        RECT 4.400 24.120 295.600 24.160 ;
        RECT 4.400 22.760 296.000 24.120 ;
        RECT 3.990 21.440 296.000 22.760 ;
        RECT 3.990 20.040 295.600 21.440 ;
        RECT 3.990 10.715 296.000 20.040 ;
      LAYER met4 ;
        RECT 30.655 32.135 97.440 240.545 ;
        RECT 99.840 32.135 174.240 240.545 ;
        RECT 176.640 32.135 251.040 240.545 ;
        RECT 253.440 32.135 289.505 240.545 ;
  END
END mac_piped
END LIBRARY

