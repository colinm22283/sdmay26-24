magic
tech sky130A
magscale 1 2
timestamp 1761579139
<< viali >>
rect 28549 27489 28583 27523
rect 27169 26945 27203 26979
rect 28365 26877 28399 26911
rect 26709 26741 26743 26775
rect 27169 26333 27203 26367
rect 26985 26265 27019 26299
rect 28365 26265 28399 26299
rect 27169 25245 27203 25279
rect 28365 25177 28399 25211
rect 26985 25109 27019 25143
rect 27169 24769 27203 24803
rect 28365 24701 28399 24735
rect 26709 24565 26743 24599
rect 1409 23681 1443 23715
rect 27169 23681 27203 23715
rect 28365 23613 28399 23647
rect 1593 23477 1627 23511
rect 26709 23477 26743 23511
rect 1593 23205 1627 23239
rect 1409 23069 1443 23103
rect 1685 23069 1719 23103
rect 27169 23069 27203 23103
rect 28365 23001 28399 23035
rect 1869 22933 1903 22967
rect 26985 22933 27019 22967
rect 1409 22593 1443 22627
rect 1685 22593 1719 22627
rect 1593 22389 1627 22423
rect 1869 22389 1903 22423
rect 28365 22049 28399 22083
rect 1409 21981 1443 22015
rect 1685 21981 1719 22015
rect 27169 21981 27203 22015
rect 1593 21845 1627 21879
rect 1869 21845 1903 21879
rect 26985 21845 27019 21879
rect 1409 21505 1443 21539
rect 1685 21505 1719 21539
rect 26709 21505 26743 21539
rect 27169 21505 27203 21539
rect 28365 21437 28399 21471
rect 1593 21369 1627 21403
rect 1869 21301 1903 21335
rect 1593 21029 1627 21063
rect 1409 20893 1443 20927
rect 1685 20893 1719 20927
rect 1869 20757 1903 20791
rect 1409 20417 1443 20451
rect 1685 20417 1719 20451
rect 27169 20417 27203 20451
rect 28365 20349 28399 20383
rect 1593 20213 1627 20247
rect 1869 20213 1903 20247
rect 26709 20213 26743 20247
rect 1593 19941 1627 19975
rect 1409 19805 1443 19839
rect 1685 19805 1719 19839
rect 27169 19805 27203 19839
rect 28365 19737 28399 19771
rect 1869 19669 1903 19703
rect 26985 19669 27019 19703
rect 1593 19465 1627 19499
rect 1869 19465 1903 19499
rect 1409 19329 1443 19363
rect 1685 19329 1719 19363
rect 12817 18921 12851 18955
rect 1593 18853 1627 18887
rect 28365 18785 28399 18819
rect 1409 18717 1443 18751
rect 1685 18717 1719 18751
rect 27169 18717 27203 18751
rect 1869 18581 1903 18615
rect 26985 18581 27019 18615
rect 12265 18377 12299 18411
rect 26709 18309 26743 18343
rect 1409 18241 1443 18275
rect 1685 18241 1719 18275
rect 9229 18241 9263 18275
rect 9413 18241 9447 18275
rect 9689 18241 9723 18275
rect 9873 18241 9907 18275
rect 12173 18241 12207 18275
rect 27169 18241 27203 18275
rect 11989 18173 12023 18207
rect 13277 18173 13311 18207
rect 28365 18173 28399 18207
rect 9597 18105 9631 18139
rect 12633 18105 12667 18139
rect 1593 18037 1627 18071
rect 1869 18037 1903 18071
rect 10057 18037 10091 18071
rect 12725 18037 12759 18071
rect 10609 17833 10643 17867
rect 1593 17765 1627 17799
rect 9229 17765 9263 17799
rect 10241 17697 10275 17731
rect 11437 17697 11471 17731
rect 13461 17697 13495 17731
rect 1409 17629 1443 17663
rect 1685 17629 1719 17663
rect 9873 17629 9907 17663
rect 10425 17629 10459 17663
rect 10701 17629 10735 17663
rect 11345 17561 11379 17595
rect 11713 17561 11747 17595
rect 1869 17493 1903 17527
rect 8493 17493 8527 17527
rect 9321 17493 9355 17527
rect 1593 17289 1627 17323
rect 9321 17289 9355 17323
rect 10057 17289 10091 17323
rect 10517 17289 10551 17323
rect 10885 17289 10919 17323
rect 9689 17221 9723 17255
rect 10149 17221 10183 17255
rect 11989 17221 12023 17255
rect 14657 17221 14691 17255
rect 1409 17153 1443 17187
rect 1685 17153 1719 17187
rect 7573 17153 7607 17187
rect 8125 17153 8159 17187
rect 8309 17153 8343 17187
rect 8493 17153 8527 17187
rect 8861 17153 8895 17187
rect 8953 17153 8987 17187
rect 10977 17153 11011 17187
rect 13737 17153 13771 17187
rect 14749 17153 14783 17187
rect 15025 17153 15059 17187
rect 27169 17153 27203 17187
rect 7205 17085 7239 17119
rect 7757 17085 7791 17119
rect 8769 17085 8803 17119
rect 9965 17085 9999 17119
rect 10701 17085 10735 17119
rect 11713 17085 11747 17119
rect 14381 17085 14415 17119
rect 28365 17085 28399 17119
rect 1869 16949 1903 16983
rect 6653 16949 6687 16983
rect 7389 16949 7423 16983
rect 11345 16949 11379 16983
rect 13829 16949 13863 16983
rect 8769 16745 8803 16779
rect 11253 16745 11287 16779
rect 6377 16609 6411 16643
rect 8125 16609 8159 16643
rect 8401 16609 8435 16643
rect 9229 16609 9263 16643
rect 11989 16609 12023 16643
rect 1409 16541 1443 16575
rect 1869 16541 1903 16575
rect 6101 16541 6135 16575
rect 8585 16541 8619 16575
rect 8953 16541 8987 16575
rect 10977 16541 11011 16575
rect 11437 16541 11471 16575
rect 11713 16541 11747 16575
rect 13737 16541 13771 16575
rect 27169 16541 27203 16575
rect 28365 16473 28399 16507
rect 1593 16405 1627 16439
rect 1685 16405 1719 16439
rect 11529 16405 11563 16439
rect 6653 16201 6687 16235
rect 6837 16201 6871 16235
rect 7297 16201 7331 16235
rect 13737 16201 13771 16235
rect 11253 16133 11287 16167
rect 13553 16133 13587 16167
rect 1409 16065 1443 16099
rect 1685 16065 1719 16099
rect 6561 16065 6595 16099
rect 7205 16065 7239 16099
rect 8033 16065 8067 16099
rect 8309 16065 8343 16099
rect 11345 16065 11379 16099
rect 11529 16065 11563 16099
rect 13829 16065 13863 16099
rect 7389 15997 7423 16031
rect 7849 15997 7883 16031
rect 8585 15997 8619 16031
rect 10333 15997 10367 16031
rect 10977 15997 11011 16031
rect 11805 15997 11839 16031
rect 10425 15929 10459 15963
rect 1593 15861 1627 15895
rect 1869 15861 1903 15895
rect 8217 15861 8251 15895
rect 9873 15657 9907 15691
rect 11989 15657 12023 15691
rect 13553 15657 13587 15691
rect 14289 15657 14323 15691
rect 1685 15589 1719 15623
rect 9689 15589 9723 15623
rect 11897 15589 11931 15623
rect 7757 15521 7791 15555
rect 9045 15521 9079 15555
rect 9229 15521 9263 15555
rect 11253 15521 11287 15555
rect 12541 15521 12575 15555
rect 1409 15453 1443 15487
rect 1869 15453 1903 15487
rect 9781 15453 9815 15487
rect 11437 15453 11471 15487
rect 13277 15453 13311 15487
rect 13645 15453 13679 15487
rect 27169 15453 27203 15487
rect 11069 15385 11103 15419
rect 11529 15385 11563 15419
rect 28365 15385 28399 15419
rect 1593 15317 1627 15351
rect 8769 15317 8803 15351
rect 9321 15317 9355 15351
rect 10333 15317 10367 15351
rect 12725 15317 12759 15351
rect 26985 15317 27019 15351
rect 1593 15113 1627 15147
rect 12909 15113 12943 15147
rect 13369 15113 13403 15147
rect 14657 15113 14691 15147
rect 12449 15045 12483 15079
rect 1409 14977 1443 15011
rect 7297 14977 7331 15011
rect 7757 14977 7791 15011
rect 12081 14977 12115 15011
rect 12541 14977 12575 15011
rect 14289 14977 14323 15011
rect 27169 14977 27203 15011
rect 6929 14909 6963 14943
rect 7481 14909 7515 14943
rect 12265 14909 12299 14943
rect 13093 14909 13127 14943
rect 13277 14909 13311 14943
rect 28365 14909 28399 14943
rect 6377 14773 6411 14807
rect 7113 14773 7147 14807
rect 7665 14773 7699 14807
rect 13737 14773 13771 14807
rect 14197 14773 14231 14807
rect 26709 14773 26743 14807
rect 1593 14569 1627 14603
rect 11437 14569 11471 14603
rect 12160 14569 12194 14603
rect 6193 14433 6227 14467
rect 11069 14433 11103 14467
rect 14657 14433 14691 14467
rect 15485 14433 15519 14467
rect 15577 14433 15611 14467
rect 1409 14365 1443 14399
rect 1685 14365 1719 14399
rect 5917 14365 5951 14399
rect 9597 14365 9631 14399
rect 10425 14365 10459 14399
rect 10609 14365 10643 14399
rect 10793 14365 10827 14399
rect 10977 14365 11011 14399
rect 11253 14365 11287 14399
rect 11897 14365 11931 14399
rect 15025 14365 15059 14399
rect 15761 14365 15795 14399
rect 7941 14297 7975 14331
rect 13921 14297 13955 14331
rect 1869 14229 1903 14263
rect 9873 14229 9907 14263
rect 14105 14229 14139 14263
rect 14933 14229 14967 14263
rect 15945 14229 15979 14263
rect 1593 14025 1627 14059
rect 1869 14025 1903 14059
rect 6561 14025 6595 14059
rect 7021 14025 7055 14059
rect 9045 14025 9079 14059
rect 9965 14025 9999 14059
rect 11161 14025 11195 14059
rect 26709 14025 26743 14059
rect 7665 13957 7699 13991
rect 10333 13957 10367 13991
rect 11713 13957 11747 13991
rect 12357 13957 12391 13991
rect 14749 13957 14783 13991
rect 15577 13957 15611 13991
rect 1409 13889 1443 13923
rect 1685 13889 1719 13923
rect 6929 13889 6963 13923
rect 9689 13889 9723 13923
rect 10793 13889 10827 13923
rect 10977 13889 11011 13923
rect 15393 13889 15427 13923
rect 15945 13889 15979 13923
rect 16405 13889 16439 13923
rect 27169 13889 27203 13923
rect 7205 13821 7239 13855
rect 9137 13821 9171 13855
rect 9321 13821 9355 13855
rect 10425 13821 10459 13855
rect 10609 13821 10643 13855
rect 12081 13821 12115 13855
rect 14105 13821 14139 13855
rect 15025 13821 15059 13855
rect 15209 13821 15243 13855
rect 15761 13821 15795 13855
rect 16129 13821 16163 13855
rect 28365 13821 28399 13855
rect 8585 13753 8619 13787
rect 8125 13685 8159 13719
rect 8677 13685 8711 13719
rect 9597 13685 9631 13719
rect 9321 13481 9355 13515
rect 26985 13481 27019 13515
rect 1869 13413 1903 13447
rect 5273 13345 5307 13379
rect 7757 13345 7791 13379
rect 8677 13345 8711 13379
rect 9413 13345 9447 13379
rect 9689 13345 9723 13379
rect 11437 13345 11471 13379
rect 16037 13345 16071 13379
rect 16681 13345 16715 13379
rect 1409 13277 1443 13311
rect 1685 13277 1719 13311
rect 5457 13277 5491 13311
rect 5733 13277 5767 13311
rect 8953 13277 8987 13311
rect 9137 13277 9171 13311
rect 11897 13277 11931 13311
rect 15577 13277 15611 13311
rect 15669 13277 15703 13311
rect 16221 13277 16255 13311
rect 27169 13277 27203 13311
rect 6009 13209 6043 13243
rect 12173 13209 12207 13243
rect 13921 13209 13955 13243
rect 15393 13209 15427 13243
rect 28365 13209 28399 13243
rect 1593 13141 1627 13175
rect 5641 13141 5675 13175
rect 8125 13141 8159 13175
rect 15853 13141 15887 13175
rect 16405 13141 16439 13175
rect 1593 12937 1627 12971
rect 5549 12937 5583 12971
rect 6745 12937 6779 12971
rect 6837 12937 6871 12971
rect 7573 12937 7607 12971
rect 10425 12937 10459 12971
rect 10977 12937 11011 12971
rect 13093 12937 13127 12971
rect 13921 12937 13955 12971
rect 14381 12937 14415 12971
rect 8125 12869 8159 12903
rect 8585 12869 8619 12903
rect 14933 12869 14967 12903
rect 1409 12801 1443 12835
rect 1685 12801 1719 12835
rect 5457 12801 5491 12835
rect 8209 12801 8243 12835
rect 8309 12801 8343 12835
rect 10609 12801 10643 12835
rect 10701 12801 10735 12835
rect 11069 12801 11103 12835
rect 12173 12801 12207 12835
rect 12633 12801 12667 12835
rect 14013 12801 14047 12835
rect 15117 12801 15151 12835
rect 15301 12801 15335 12835
rect 16129 12801 16163 12835
rect 6193 12733 6227 12767
rect 7021 12733 7055 12767
rect 7297 12733 7331 12767
rect 7481 12733 7515 12767
rect 10333 12733 10367 12767
rect 12449 12733 12483 12767
rect 12541 12733 12575 12767
rect 13645 12733 13679 12767
rect 15853 12733 15887 12767
rect 15945 12733 15979 12767
rect 1869 12665 1903 12699
rect 6377 12665 6411 12699
rect 7941 12665 7975 12699
rect 13001 12665 13035 12699
rect 15485 12597 15519 12631
rect 16313 12597 16347 12631
rect 15209 12393 15243 12427
rect 16313 12393 16347 12427
rect 1593 12325 1627 12359
rect 5733 12325 5767 12359
rect 10149 12325 10183 12359
rect 11437 12325 11471 12359
rect 13001 12325 13035 12359
rect 7389 12257 7423 12291
rect 9505 12257 9539 12291
rect 10793 12257 10827 12291
rect 11897 12257 11931 12291
rect 11989 12257 12023 12291
rect 12449 12257 12483 12291
rect 13645 12257 13679 12291
rect 15393 12257 15427 12291
rect 16497 12257 16531 12291
rect 1409 12189 1443 12223
rect 1685 12189 1719 12223
rect 8125 12189 8159 12223
rect 8953 12189 8987 12223
rect 9873 12189 9907 12223
rect 9965 12189 9999 12223
rect 10517 12189 10551 12223
rect 11345 12189 11379 12223
rect 12541 12189 12575 12223
rect 14105 12189 14139 12223
rect 15577 12189 15611 12223
rect 16681 12189 16715 12223
rect 27169 12189 27203 12223
rect 7021 12121 7055 12155
rect 11805 12121 11839 12155
rect 12633 12121 12667 12155
rect 15761 12121 15795 12155
rect 28365 12121 28399 12155
rect 1869 12053 1903 12087
rect 5181 12053 5215 12087
rect 7573 12053 7607 12087
rect 7665 12053 7699 12087
rect 8033 12053 8067 12087
rect 8769 12053 8803 12087
rect 10425 12053 10459 12087
rect 13093 12053 13127 12087
rect 14197 12053 14231 12087
rect 16865 12053 16899 12087
rect 6009 11849 6043 11883
rect 6837 11849 6871 11883
rect 9873 11849 9907 11883
rect 17693 11849 17727 11883
rect 12265 11781 12299 11815
rect 1409 11713 1443 11747
rect 1685 11713 1719 11747
rect 5641 11713 5675 11747
rect 5825 11713 5859 11747
rect 6469 11713 6503 11747
rect 6653 11713 6687 11747
rect 9229 11713 9263 11747
rect 10333 11713 10367 11747
rect 11713 11713 11747 11747
rect 11989 11713 12023 11747
rect 14013 11713 14047 11747
rect 17049 11713 17083 11747
rect 17141 11713 17175 11747
rect 27169 11713 27203 11747
rect 6929 11645 6963 11679
rect 8677 11645 8711 11679
rect 8953 11645 8987 11679
rect 9045 11645 9079 11679
rect 10701 11645 10735 11679
rect 28365 11645 28399 11679
rect 1593 11577 1627 11611
rect 1869 11509 1903 11543
rect 9413 11509 9447 11543
rect 11345 11509 11379 11543
rect 11805 11509 11839 11543
rect 17325 11509 17359 11543
rect 26709 11509 26743 11543
rect 11437 11305 11471 11339
rect 1593 11237 1627 11271
rect 4905 11169 4939 11203
rect 5273 11169 5307 11203
rect 8217 11169 8251 11203
rect 8585 11169 8619 11203
rect 8953 11169 8987 11203
rect 9321 11169 9355 11203
rect 9689 11169 9723 11203
rect 10793 11169 10827 11203
rect 1409 11101 1443 11135
rect 1685 11101 1719 11135
rect 5089 11101 5123 11135
rect 5917 11101 5951 11135
rect 6101 11101 6135 11135
rect 8401 11101 8435 11135
rect 9137 11101 9171 11135
rect 9873 11101 9907 11135
rect 11529 11101 11563 11135
rect 13553 11101 13587 11135
rect 14197 11101 14231 11135
rect 14289 11101 14323 11135
rect 6377 11033 6411 11067
rect 8125 11033 8159 11067
rect 10977 11033 11011 11067
rect 11069 11033 11103 11067
rect 11805 11033 11839 11067
rect 14473 11033 14507 11067
rect 1869 10965 1903 10999
rect 5365 10965 5399 10999
rect 10057 10965 10091 10999
rect 5457 10761 5491 10795
rect 7573 10761 7607 10795
rect 10517 10761 10551 10795
rect 4905 10693 4939 10727
rect 13553 10693 13587 10727
rect 15669 10693 15703 10727
rect 1409 10625 1443 10659
rect 1685 10625 1719 10659
rect 4997 10625 5031 10659
rect 5181 10625 5215 10659
rect 5825 10625 5859 10659
rect 6561 10625 6595 10659
rect 7205 10625 7239 10659
rect 7665 10625 7699 10659
rect 7849 10625 7883 10659
rect 13737 10625 13771 10659
rect 13829 10625 13863 10659
rect 15761 10625 15795 10659
rect 15945 10625 15979 10659
rect 27169 10625 27203 10659
rect 5365 10557 5399 10591
rect 5917 10557 5951 10591
rect 6101 10557 6135 10591
rect 9597 10557 9631 10591
rect 10333 10557 10367 10591
rect 11069 10557 11103 10591
rect 11529 10557 11563 10591
rect 11805 10557 11839 10591
rect 28365 10557 28399 10591
rect 1593 10489 1627 10523
rect 1869 10421 1903 10455
rect 4537 10421 4571 10455
rect 9781 10421 9815 10455
rect 14013 10421 14047 10455
rect 16129 10421 16163 10455
rect 8677 10217 8711 10251
rect 9873 10217 9907 10251
rect 11897 10217 11931 10251
rect 12725 10217 12759 10251
rect 26985 10217 27019 10251
rect 1869 10149 1903 10183
rect 11713 10149 11747 10183
rect 4997 10081 5031 10115
rect 7297 10081 7331 10115
rect 9965 10081 9999 10115
rect 10241 10081 10275 10115
rect 12449 10081 12483 10115
rect 1409 10013 1443 10047
rect 1685 10013 1719 10047
rect 8125 10013 8159 10047
rect 9321 10013 9355 10047
rect 12817 10013 12851 10047
rect 27169 10013 27203 10047
rect 5273 9945 5307 9979
rect 7021 9945 7055 9979
rect 28365 9945 28399 9979
rect 1593 9877 1627 9911
rect 2237 9877 2271 9911
rect 4813 9877 4847 9911
rect 1869 9673 1903 9707
rect 4629 9605 4663 9639
rect 4813 9605 4847 9639
rect 7021 9605 7055 9639
rect 9597 9605 9631 9639
rect 10701 9605 10735 9639
rect 1409 9537 1443 9571
rect 1685 9537 1719 9571
rect 1961 9537 1995 9571
rect 2237 9537 2271 9571
rect 4905 9537 4939 9571
rect 5089 9537 5123 9571
rect 5181 9535 5215 9569
rect 6193 9537 6227 9571
rect 6377 9537 6411 9571
rect 7113 9537 7147 9571
rect 9045 9537 9079 9571
rect 9229 9537 9263 9571
rect 10241 9537 10275 9571
rect 11345 9537 11379 9571
rect 12173 9537 12207 9571
rect 14197 9537 14231 9571
rect 10793 9469 10827 9503
rect 10977 9469 11011 9503
rect 11253 9469 11287 9503
rect 14013 9469 14047 9503
rect 1593 9401 1627 9435
rect 2145 9333 2179 9367
rect 2421 9333 2455 9367
rect 2789 9333 2823 9367
rect 3157 9333 3191 9367
rect 4169 9333 4203 9367
rect 5365 9333 5399 9367
rect 5549 9333 5583 9367
rect 8401 9333 8435 9367
rect 9413 9333 9447 9367
rect 10333 9333 10367 9367
rect 11805 9333 11839 9367
rect 14381 9333 14415 9367
rect 1869 9129 1903 9163
rect 5641 9129 5675 9163
rect 8125 9129 8159 9163
rect 1593 9061 1627 9095
rect 4721 9061 4755 9095
rect 4813 8993 4847 9027
rect 6101 8993 6135 9027
rect 7849 8993 7883 9027
rect 8769 8993 8803 9027
rect 12081 8993 12115 9027
rect 28365 8993 28399 9027
rect 1409 8925 1443 8959
rect 1685 8925 1719 8959
rect 2145 8925 2179 8959
rect 2237 8925 2271 8959
rect 2697 8925 2731 8959
rect 4997 8925 5031 8959
rect 5365 8925 5399 8959
rect 5457 8925 5491 8959
rect 5825 8925 5859 8959
rect 8953 8925 8987 8959
rect 10885 8925 10919 8959
rect 11069 8925 11103 8959
rect 12265 8925 12299 8959
rect 27169 8925 27203 8959
rect 9229 8857 9263 8891
rect 11253 8857 11287 8891
rect 1961 8789 1995 8823
rect 2421 8789 2455 8823
rect 2513 8789 2547 8823
rect 3249 8789 3283 8823
rect 3617 8789 3651 8823
rect 4353 8789 4387 8823
rect 5181 8789 5215 8823
rect 10701 8789 10735 8823
rect 11621 8789 11655 8823
rect 12449 8789 12483 8823
rect 1593 8585 1627 8619
rect 2421 8585 2455 8619
rect 2789 8585 2823 8619
rect 6377 8585 6411 8619
rect 6745 8585 6779 8619
rect 7205 8585 7239 8619
rect 8585 8585 8619 8619
rect 9505 8585 9539 8619
rect 10701 8585 10735 8619
rect 11529 8585 11563 8619
rect 5457 8517 5491 8551
rect 6837 8517 6871 8551
rect 9045 8517 9079 8551
rect 1409 8449 1443 8483
rect 1685 8449 1719 8483
rect 1961 8449 1995 8483
rect 2237 8449 2271 8483
rect 2697 8449 2731 8483
rect 2973 8449 3007 8483
rect 3249 8449 3283 8483
rect 3341 8449 3375 8483
rect 4905 8449 4939 8483
rect 5089 8449 5123 8483
rect 8033 8449 8067 8483
rect 10333 8449 10367 8483
rect 10425 8449 10459 8483
rect 10609 8449 10643 8483
rect 27169 8449 27203 8483
rect 6101 8381 6135 8415
rect 6929 8381 6963 8415
rect 7757 8381 7791 8415
rect 8769 8381 8803 8415
rect 8953 8381 8987 8415
rect 10057 8381 10091 8415
rect 11253 8381 11287 8415
rect 12173 8381 12207 8415
rect 28365 8381 28399 8415
rect 1869 8313 1903 8347
rect 2513 8313 2547 8347
rect 3065 8313 3099 8347
rect 3525 8313 3559 8347
rect 4077 8313 4111 8347
rect 4445 8313 4479 8347
rect 4813 8313 4847 8347
rect 5273 8313 5307 8347
rect 9413 8313 9447 8347
rect 26709 8313 26743 8347
rect 2145 8245 2179 8279
rect 8585 8041 8619 8075
rect 8953 8041 8987 8075
rect 11069 8041 11103 8075
rect 26985 8041 27019 8075
rect 7757 7973 7791 8007
rect 3249 7905 3283 7939
rect 3801 7905 3835 7939
rect 4629 7905 4663 7939
rect 5457 7905 5491 7939
rect 7389 7905 7423 7939
rect 27629 7905 27663 7939
rect 1777 7837 1811 7871
rect 2237 7837 2271 7871
rect 2513 7837 2547 7871
rect 2973 7837 3007 7871
rect 3433 7837 3467 7871
rect 3985 7837 4019 7871
rect 4353 7837 4387 7871
rect 4813 7837 4847 7871
rect 5181 7837 5215 7871
rect 7573 7837 7607 7871
rect 7941 7837 7975 7871
rect 9597 7837 9631 7871
rect 9781 7837 9815 7871
rect 9873 7837 9907 7871
rect 10425 7837 10459 7871
rect 10977 7837 11011 7871
rect 11713 7837 11747 7871
rect 27169 7837 27203 7871
rect 1961 7769 1995 7803
rect 3617 7769 3651 7803
rect 7205 7769 7239 7803
rect 1409 7701 1443 7735
rect 1593 7701 1627 7735
rect 1685 7701 1719 7735
rect 2421 7701 2455 7735
rect 2697 7701 2731 7735
rect 3065 7701 3099 7735
rect 4169 7701 4203 7735
rect 4445 7701 4479 7735
rect 4997 7701 5031 7735
rect 10057 7701 10091 7735
rect 1777 7497 1811 7531
rect 3249 7497 3283 7531
rect 5917 7497 5951 7531
rect 6377 7497 6411 7531
rect 8033 7497 8067 7531
rect 8217 7497 8251 7531
rect 9781 7497 9815 7531
rect 3341 7429 3375 7463
rect 5825 7429 5859 7463
rect 7113 7429 7147 7463
rect 10517 7429 10551 7463
rect 26617 7429 26651 7463
rect 1593 7361 1627 7395
rect 2605 7361 2639 7395
rect 4169 7361 4203 7395
rect 4353 7361 4387 7395
rect 4537 7361 4571 7395
rect 4905 7361 4939 7395
rect 4997 7361 5031 7395
rect 8125 7361 8159 7395
rect 9137 7361 9171 7395
rect 9689 7361 9723 7395
rect 10057 7361 10091 7395
rect 10149 7361 10183 7395
rect 10885 7361 10919 7395
rect 25421 7361 25455 7395
rect 27169 7361 27203 7395
rect 1961 7293 1995 7327
rect 3893 7293 3927 7327
rect 4813 7293 4847 7327
rect 6009 7293 6043 7327
rect 7021 7293 7055 7327
rect 7757 7293 7791 7327
rect 8769 7293 8803 7327
rect 8953 7293 8987 7327
rect 28365 7293 28399 7327
rect 2513 7225 2547 7259
rect 5365 7225 5399 7259
rect 5457 7157 5491 7191
rect 9321 7157 9355 7191
rect 11161 7157 11195 7191
rect 1501 6817 1535 6851
rect 3893 6817 3927 6851
rect 4997 6817 5031 6851
rect 5089 6817 5123 6851
rect 7113 6817 7147 6851
rect 8493 6817 8527 6851
rect 8677 6817 8711 6851
rect 9597 6817 9631 6851
rect 9689 6817 9723 6851
rect 1685 6749 1719 6783
rect 1961 6749 1995 6783
rect 2513 6749 2547 6783
rect 2697 6749 2731 6783
rect 2973 6749 3007 6783
rect 3617 6749 3651 6783
rect 4077 6749 4111 6783
rect 4353 6749 4387 6783
rect 7389 6749 7423 6783
rect 8953 6749 8987 6783
rect 9873 6749 9907 6783
rect 10057 6749 10091 6783
rect 25697 6749 25731 6783
rect 27169 6749 27203 6783
rect 4261 6681 4295 6715
rect 5365 6681 5399 6715
rect 8401 6681 8435 6715
rect 10333 6681 10367 6715
rect 25513 6681 25547 6715
rect 26893 6681 26927 6715
rect 28365 6681 28399 6715
rect 1869 6613 1903 6647
rect 2881 6613 2915 6647
rect 7941 6613 7975 6647
rect 8033 6613 8067 6647
rect 10793 6613 10827 6647
rect 2053 6409 2087 6443
rect 4629 6409 4663 6443
rect 5365 6409 5399 6443
rect 6377 6409 6411 6443
rect 10149 6409 10183 6443
rect 5917 6273 5951 6307
rect 7113 6273 7147 6307
rect 7297 6273 7331 6307
rect 7757 6273 7791 6307
rect 9781 6273 9815 6307
rect 23949 6273 23983 6307
rect 25421 6273 25455 6307
rect 27169 6273 27203 6307
rect 1501 6205 1535 6239
rect 2237 6205 2271 6239
rect 3065 6205 3099 6239
rect 4445 6205 4479 6239
rect 5273 6205 5307 6239
rect 7021 6205 7055 6239
rect 8033 6205 8067 6239
rect 24685 6205 24719 6239
rect 26157 6205 26191 6239
rect 28365 6205 28399 6239
rect 3617 6137 3651 6171
rect 2789 6069 2823 6103
rect 3893 6069 3927 6103
rect 7481 6069 7515 6103
rect 10517 6069 10551 6103
rect 23765 6069 23799 6103
rect 2789 5865 2823 5899
rect 3525 5865 3559 5899
rect 4242 5865 4276 5899
rect 7573 5865 7607 5899
rect 8677 5865 8711 5899
rect 9045 5865 9079 5899
rect 9413 5865 9447 5899
rect 9873 5865 9907 5899
rect 10241 5865 10275 5899
rect 2053 5797 2087 5831
rect 7941 5797 7975 5831
rect 2881 5729 2915 5763
rect 3985 5729 4019 5763
rect 26433 5729 26467 5763
rect 28365 5729 28399 5763
rect 1501 5661 1535 5695
rect 2237 5661 2271 5695
rect 8125 5661 8159 5695
rect 8401 5661 8435 5695
rect 9137 5661 9171 5695
rect 22845 5661 22879 5695
rect 25697 5661 25731 5695
rect 27169 5661 27203 5695
rect 6009 5593 6043 5627
rect 6101 5593 6135 5627
rect 24041 5593 24075 5627
rect 8217 5525 8251 5559
rect 3065 5321 3099 5355
rect 4445 5321 4479 5355
rect 5457 5321 5491 5355
rect 6469 5321 6503 5355
rect 8677 5321 8711 5355
rect 26709 5321 26743 5355
rect 4353 5253 4387 5287
rect 7757 5253 7791 5287
rect 9873 5253 9907 5287
rect 10517 5253 10551 5287
rect 1409 5185 1443 5219
rect 1593 5185 1627 5219
rect 4813 5185 4847 5219
rect 6561 5185 6595 5219
rect 8401 5185 8435 5219
rect 8493 5185 8527 5219
rect 8953 5185 8987 5219
rect 9229 5185 9263 5219
rect 9505 5185 9539 5219
rect 21925 5185 21959 5219
rect 23489 5185 23523 5219
rect 24869 5185 24903 5219
rect 26985 5185 27019 5219
rect 1961 5117 1995 5151
rect 4905 5117 4939 5151
rect 4997 5117 5031 5151
rect 6101 5117 6135 5151
rect 7297 5117 7331 5151
rect 7849 5117 7883 5151
rect 8033 5117 8067 5151
rect 23121 5117 23155 5151
rect 24593 5117 24627 5151
rect 25329 5117 25363 5151
rect 27445 5117 27479 5151
rect 1777 5049 1811 5083
rect 7389 5049 7423 5083
rect 9045 5049 9079 5083
rect 2513 4981 2547 5015
rect 6653 4981 6687 5015
rect 8217 4981 8251 5015
rect 8769 4981 8803 5015
rect 9413 4981 9447 5015
rect 10241 4981 10275 5015
rect 10977 4981 11011 5015
rect 3801 4777 3835 4811
rect 3985 4777 4019 4811
rect 5089 4777 5123 4811
rect 5917 4777 5951 4811
rect 9413 4777 9447 4811
rect 10149 4777 10183 4811
rect 2881 4709 2915 4743
rect 3617 4709 3651 4743
rect 4353 4709 4387 4743
rect 1501 4641 1535 4675
rect 5825 4641 5859 4675
rect 6561 4641 6595 4675
rect 7021 4641 7055 4675
rect 8769 4641 8803 4675
rect 8953 4641 8987 4675
rect 10609 4641 10643 4675
rect 25053 4641 25087 4675
rect 26341 4641 26375 4675
rect 2237 4573 2271 4607
rect 3065 4573 3099 4607
rect 4537 4573 4571 4607
rect 5181 4573 5215 4607
rect 6745 4573 6779 4607
rect 9137 4573 9171 4607
rect 9597 4573 9631 4607
rect 9873 4573 9907 4607
rect 21373 4573 21407 4607
rect 22845 4573 22879 4607
rect 24409 4573 24443 4607
rect 25881 4573 25915 4607
rect 2145 4505 2179 4539
rect 22569 4505 22603 4539
rect 24041 4505 24075 4539
rect 3985 4437 4019 4471
rect 9321 4437 9355 4471
rect 9689 4437 9723 4471
rect 10977 4437 11011 4471
rect 1685 4233 1719 4267
rect 4169 4233 4203 4267
rect 8493 4233 8527 4267
rect 9229 4233 9263 4267
rect 2697 4165 2731 4199
rect 4905 4165 4939 4199
rect 9873 4165 9907 4199
rect 10793 4165 10827 4199
rect 1593 4097 1627 4131
rect 2329 4097 2363 4131
rect 5733 4097 5767 4131
rect 5825 4097 5859 4131
rect 9321 4097 9355 4131
rect 9505 4097 9539 4131
rect 9965 4097 9999 4131
rect 10241 4097 10275 4131
rect 10517 4097 10551 4131
rect 20269 4097 20303 4131
rect 22385 4097 22419 4131
rect 23857 4097 23891 4131
rect 25329 4097 25363 4131
rect 27169 4097 27203 4131
rect 2421 4029 2455 4063
rect 4997 4029 5031 4063
rect 5089 4029 5123 4063
rect 5549 4029 5583 4063
rect 6929 4029 6963 4063
rect 7113 4029 7147 4063
rect 7849 4029 7883 4063
rect 8585 4029 8619 4063
rect 9689 4029 9723 4063
rect 21465 4029 21499 4063
rect 22845 4029 22879 4063
rect 24317 4029 24351 4063
rect 25789 4029 25823 4063
rect 27445 4029 27479 4063
rect 6193 3961 6227 3995
rect 11805 3961 11839 3995
rect 1501 3893 1535 3927
rect 4537 3893 4571 3927
rect 6377 3893 6411 3927
rect 7757 3893 7791 3927
rect 10057 3893 10091 3927
rect 10333 3893 10367 3927
rect 11253 3893 11287 3927
rect 1685 3689 1719 3723
rect 5181 3689 5215 3723
rect 8585 3689 8619 3723
rect 10425 3689 10459 3723
rect 10701 3689 10735 3723
rect 11345 3689 11379 3723
rect 11897 3689 11931 3723
rect 12173 3689 12207 3723
rect 24133 3689 24167 3723
rect 27537 3689 27571 3723
rect 3433 3553 3467 3587
rect 5273 3553 5307 3587
rect 5549 3553 5583 3587
rect 22017 3553 22051 3587
rect 24869 3553 24903 3587
rect 26341 3553 26375 3587
rect 1501 3485 1535 3519
rect 3166 3485 3200 3519
rect 3801 3485 3835 3519
rect 4813 3485 4847 3519
rect 4997 3485 5031 3519
rect 7297 3485 7331 3519
rect 7481 3485 7515 3519
rect 7573 3485 7607 3519
rect 7941 3485 7975 3519
rect 8953 3485 8987 3519
rect 9781 3485 9815 3519
rect 10517 3485 10551 3519
rect 10977 3485 11011 3519
rect 11253 3485 11287 3519
rect 11529 3485 11563 3519
rect 20085 3485 20119 3519
rect 21557 3485 21591 3519
rect 24409 3485 24443 3519
rect 25881 3485 25915 3519
rect 28549 3485 28583 3519
rect 4537 3417 4571 3451
rect 7757 3417 7791 3451
rect 21281 3417 21315 3451
rect 2053 3349 2087 3383
rect 9597 3349 9631 3383
rect 10793 3349 10827 3383
rect 11069 3349 11103 3383
rect 2237 3145 2271 3179
rect 7573 3145 7607 3179
rect 8309 3145 8343 3179
rect 9045 3145 9079 3179
rect 10609 3145 10643 3179
rect 11529 3145 11563 3179
rect 11805 3145 11839 3179
rect 12081 3145 12115 3179
rect 12357 3145 12391 3179
rect 2145 3077 2179 3111
rect 6193 3077 6227 3111
rect 19993 3077 20027 3111
rect 2605 3009 2639 3043
rect 3065 3009 3099 3043
rect 3893 3009 3927 3043
rect 4169 3009 4203 3043
rect 6377 3009 6411 3043
rect 6561 3009 6595 3043
rect 11713 3009 11747 3043
rect 11989 3009 12023 3043
rect 12265 3009 12299 3043
rect 12541 3009 12575 3043
rect 18797 3009 18831 3043
rect 20269 3009 20303 3043
rect 21833 3009 21867 3043
rect 23305 3009 23339 3043
rect 24961 3009 24995 3043
rect 26985 3009 27019 3043
rect 1593 2941 1627 2975
rect 2697 2941 2731 2975
rect 2881 2941 2915 2975
rect 4445 2941 4479 2975
rect 7021 2941 7055 2975
rect 7757 2941 7791 2975
rect 8493 2941 8527 2975
rect 9229 2941 9263 2975
rect 9873 2941 9907 2975
rect 10425 2941 10459 2975
rect 11161 2941 11195 2975
rect 21465 2941 21499 2975
rect 22293 2941 22327 2975
rect 23765 2941 23799 2975
rect 25237 2941 25271 2975
rect 27445 2941 27479 2975
rect 6745 2873 6779 2907
rect 9781 2805 9815 2839
rect 3985 2601 4019 2635
rect 6561 2601 6595 2635
rect 8033 2601 8067 2635
rect 11345 2601 11379 2635
rect 12265 2601 12299 2635
rect 12541 2601 12575 2635
rect 9137 2533 9171 2567
rect 2329 2465 2363 2499
rect 4077 2465 4111 2499
rect 5549 2465 5583 2499
rect 6193 2465 6227 2499
rect 8125 2465 8159 2499
rect 10609 2465 10643 2499
rect 20729 2465 20763 2499
rect 22293 2465 22327 2499
rect 24869 2465 24903 2499
rect 27445 2465 27479 2499
rect 1593 2397 1627 2431
rect 3065 2397 3099 2431
rect 3801 2397 3835 2431
rect 4721 2397 4755 2431
rect 4905 2397 4939 2431
rect 6377 2397 6411 2431
rect 7297 2397 7331 2431
rect 7481 2397 7515 2431
rect 8769 2397 8803 2431
rect 8953 2397 8987 2431
rect 9321 2397 9355 2431
rect 10057 2397 10091 2431
rect 10793 2397 10827 2431
rect 11529 2397 11563 2431
rect 12173 2397 12207 2431
rect 12449 2397 12483 2431
rect 12725 2397 12759 2431
rect 13001 2397 13035 2431
rect 13277 2397 13311 2431
rect 17693 2397 17727 2431
rect 20269 2397 20303 2431
rect 21833 2397 21867 2431
rect 24409 2397 24443 2431
rect 26985 2397 27019 2431
rect 6653 2329 6687 2363
rect 18889 2329 18923 2363
rect 2145 2261 2179 2295
rect 2881 2261 2915 2295
rect 3617 2261 3651 2295
rect 5457 2261 5491 2295
rect 9873 2261 9907 2295
rect 12817 2261 12851 2295
rect 13093 2261 13127 2295
rect 20085 2261 20119 2295
rect 26709 2261 26743 2295
<< metal1 >>
rect 1104 27770 28888 27792
rect 1104 27718 4423 27770
rect 4475 27718 4487 27770
rect 4539 27718 4551 27770
rect 4603 27718 4615 27770
rect 4667 27718 4679 27770
rect 4731 27718 11369 27770
rect 11421 27718 11433 27770
rect 11485 27718 11497 27770
rect 11549 27718 11561 27770
rect 11613 27718 11625 27770
rect 11677 27718 18315 27770
rect 18367 27718 18379 27770
rect 18431 27718 18443 27770
rect 18495 27718 18507 27770
rect 18559 27718 18571 27770
rect 18623 27718 25261 27770
rect 25313 27718 25325 27770
rect 25377 27718 25389 27770
rect 25441 27718 25453 27770
rect 25505 27718 25517 27770
rect 25569 27718 28888 27770
rect 1104 27696 28888 27718
rect 28534 27480 28540 27532
rect 28592 27480 28598 27532
rect 1104 27226 29048 27248
rect 1104 27174 7896 27226
rect 7948 27174 7960 27226
rect 8012 27174 8024 27226
rect 8076 27174 8088 27226
rect 8140 27174 8152 27226
rect 8204 27174 14842 27226
rect 14894 27174 14906 27226
rect 14958 27174 14970 27226
rect 15022 27174 15034 27226
rect 15086 27174 15098 27226
rect 15150 27174 21788 27226
rect 21840 27174 21852 27226
rect 21904 27174 21916 27226
rect 21968 27174 21980 27226
rect 22032 27174 22044 27226
rect 22096 27174 28734 27226
rect 28786 27174 28798 27226
rect 28850 27174 28862 27226
rect 28914 27174 28926 27226
rect 28978 27174 28990 27226
rect 29042 27174 29048 27226
rect 1104 27152 29048 27174
rect 27157 26979 27215 26985
rect 27157 26976 27169 26979
rect 26712 26948 27169 26976
rect 22738 26732 22744 26784
rect 22796 26772 22802 26784
rect 26712 26781 26740 26948
rect 27157 26945 27169 26948
rect 27203 26945 27215 26979
rect 27157 26939 27215 26945
rect 28350 26868 28356 26920
rect 28408 26868 28414 26920
rect 26697 26775 26755 26781
rect 26697 26772 26709 26775
rect 22796 26744 26709 26772
rect 22796 26732 22802 26744
rect 26697 26741 26709 26744
rect 26743 26741 26755 26775
rect 26697 26735 26755 26741
rect 1104 26682 28888 26704
rect 1104 26630 4423 26682
rect 4475 26630 4487 26682
rect 4539 26630 4551 26682
rect 4603 26630 4615 26682
rect 4667 26630 4679 26682
rect 4731 26630 11369 26682
rect 11421 26630 11433 26682
rect 11485 26630 11497 26682
rect 11549 26630 11561 26682
rect 11613 26630 11625 26682
rect 11677 26630 18315 26682
rect 18367 26630 18379 26682
rect 18431 26630 18443 26682
rect 18495 26630 18507 26682
rect 18559 26630 18571 26682
rect 18623 26630 25261 26682
rect 25313 26630 25325 26682
rect 25377 26630 25389 26682
rect 25441 26630 25453 26682
rect 25505 26630 25517 26682
rect 25569 26630 28888 26682
rect 1104 26608 28888 26630
rect 27157 26367 27215 26373
rect 27157 26333 27169 26367
rect 27203 26333 27215 26367
rect 27157 26327 27215 26333
rect 14274 26256 14280 26308
rect 14332 26296 14338 26308
rect 26973 26299 27031 26305
rect 26973 26296 26985 26299
rect 14332 26268 26985 26296
rect 14332 26256 14338 26268
rect 26973 26265 26985 26268
rect 27019 26296 27031 26299
rect 27172 26296 27200 26327
rect 27019 26268 27200 26296
rect 27019 26265 27031 26268
rect 26973 26259 27031 26265
rect 28350 26256 28356 26308
rect 28408 26256 28414 26308
rect 1104 26138 29048 26160
rect 1104 26086 7896 26138
rect 7948 26086 7960 26138
rect 8012 26086 8024 26138
rect 8076 26086 8088 26138
rect 8140 26086 8152 26138
rect 8204 26086 14842 26138
rect 14894 26086 14906 26138
rect 14958 26086 14970 26138
rect 15022 26086 15034 26138
rect 15086 26086 15098 26138
rect 15150 26086 21788 26138
rect 21840 26086 21852 26138
rect 21904 26086 21916 26138
rect 21968 26086 21980 26138
rect 22032 26086 22044 26138
rect 22096 26086 28734 26138
rect 28786 26086 28798 26138
rect 28850 26086 28862 26138
rect 28914 26086 28926 26138
rect 28978 26086 28990 26138
rect 29042 26086 29048 26138
rect 1104 26064 29048 26086
rect 1104 25594 28888 25616
rect 1104 25542 4423 25594
rect 4475 25542 4487 25594
rect 4539 25542 4551 25594
rect 4603 25542 4615 25594
rect 4667 25542 4679 25594
rect 4731 25542 11369 25594
rect 11421 25542 11433 25594
rect 11485 25542 11497 25594
rect 11549 25542 11561 25594
rect 11613 25542 11625 25594
rect 11677 25542 18315 25594
rect 18367 25542 18379 25594
rect 18431 25542 18443 25594
rect 18495 25542 18507 25594
rect 18559 25542 18571 25594
rect 18623 25542 25261 25594
rect 25313 25542 25325 25594
rect 25377 25542 25389 25594
rect 25441 25542 25453 25594
rect 25505 25542 25517 25594
rect 25569 25542 28888 25594
rect 1104 25520 28888 25542
rect 27157 25279 27215 25285
rect 27157 25245 27169 25279
rect 27203 25245 27215 25279
rect 27157 25239 27215 25245
rect 25682 25100 25688 25152
rect 25740 25140 25746 25152
rect 26973 25143 27031 25149
rect 26973 25140 26985 25143
rect 25740 25112 26985 25140
rect 25740 25100 25746 25112
rect 26973 25109 26985 25112
rect 27019 25140 27031 25143
rect 27172 25140 27200 25239
rect 28350 25168 28356 25220
rect 28408 25168 28414 25220
rect 27019 25112 27200 25140
rect 27019 25109 27031 25112
rect 26973 25103 27031 25109
rect 1104 25050 29048 25072
rect 1104 24998 7896 25050
rect 7948 24998 7960 25050
rect 8012 24998 8024 25050
rect 8076 24998 8088 25050
rect 8140 24998 8152 25050
rect 8204 24998 14842 25050
rect 14894 24998 14906 25050
rect 14958 24998 14970 25050
rect 15022 24998 15034 25050
rect 15086 24998 15098 25050
rect 15150 24998 21788 25050
rect 21840 24998 21852 25050
rect 21904 24998 21916 25050
rect 21968 24998 21980 25050
rect 22032 24998 22044 25050
rect 22096 24998 28734 25050
rect 28786 24998 28798 25050
rect 28850 24998 28862 25050
rect 28914 24998 28926 25050
rect 28978 24998 28990 25050
rect 29042 24998 29048 25050
rect 1104 24976 29048 24998
rect 27157 24803 27215 24809
rect 27157 24800 27169 24803
rect 26712 24772 27169 24800
rect 12802 24556 12808 24608
rect 12860 24596 12866 24608
rect 26712 24605 26740 24772
rect 27157 24769 27169 24772
rect 27203 24769 27215 24803
rect 27157 24763 27215 24769
rect 28350 24692 28356 24744
rect 28408 24692 28414 24744
rect 26697 24599 26755 24605
rect 26697 24596 26709 24599
rect 12860 24568 26709 24596
rect 12860 24556 12866 24568
rect 26697 24565 26709 24568
rect 26743 24565 26755 24599
rect 26697 24559 26755 24565
rect 1104 24506 28888 24528
rect 1104 24454 4423 24506
rect 4475 24454 4487 24506
rect 4539 24454 4551 24506
rect 4603 24454 4615 24506
rect 4667 24454 4679 24506
rect 4731 24454 11369 24506
rect 11421 24454 11433 24506
rect 11485 24454 11497 24506
rect 11549 24454 11561 24506
rect 11613 24454 11625 24506
rect 11677 24454 18315 24506
rect 18367 24454 18379 24506
rect 18431 24454 18443 24506
rect 18495 24454 18507 24506
rect 18559 24454 18571 24506
rect 18623 24454 25261 24506
rect 25313 24454 25325 24506
rect 25377 24454 25389 24506
rect 25441 24454 25453 24506
rect 25505 24454 25517 24506
rect 25569 24454 28888 24506
rect 1104 24432 28888 24454
rect 1104 23962 29048 23984
rect 1104 23910 7896 23962
rect 7948 23910 7960 23962
rect 8012 23910 8024 23962
rect 8076 23910 8088 23962
rect 8140 23910 8152 23962
rect 8204 23910 14842 23962
rect 14894 23910 14906 23962
rect 14958 23910 14970 23962
rect 15022 23910 15034 23962
rect 15086 23910 15098 23962
rect 15150 23910 21788 23962
rect 21840 23910 21852 23962
rect 21904 23910 21916 23962
rect 21968 23910 21980 23962
rect 22032 23910 22044 23962
rect 22096 23910 28734 23962
rect 28786 23910 28798 23962
rect 28850 23910 28862 23962
rect 28914 23910 28926 23962
rect 28978 23910 28990 23962
rect 29042 23910 29048 23962
rect 1104 23888 29048 23910
rect 1394 23672 1400 23724
rect 1452 23672 1458 23724
rect 27157 23715 27215 23721
rect 27157 23712 27169 23715
rect 26712 23684 27169 23712
rect 1578 23468 1584 23520
rect 1636 23468 1642 23520
rect 25774 23468 25780 23520
rect 25832 23508 25838 23520
rect 26712 23517 26740 23684
rect 27157 23681 27169 23684
rect 27203 23681 27215 23715
rect 27157 23675 27215 23681
rect 28353 23647 28411 23653
rect 28353 23613 28365 23647
rect 28399 23644 28411 23647
rect 28718 23644 28724 23656
rect 28399 23616 28724 23644
rect 28399 23613 28411 23616
rect 28353 23607 28411 23613
rect 28718 23604 28724 23616
rect 28776 23604 28782 23656
rect 26697 23511 26755 23517
rect 26697 23508 26709 23511
rect 25832 23480 26709 23508
rect 25832 23468 25838 23480
rect 26697 23477 26709 23480
rect 26743 23477 26755 23511
rect 26697 23471 26755 23477
rect 1104 23418 28888 23440
rect 1104 23366 4423 23418
rect 4475 23366 4487 23418
rect 4539 23366 4551 23418
rect 4603 23366 4615 23418
rect 4667 23366 4679 23418
rect 4731 23366 11369 23418
rect 11421 23366 11433 23418
rect 11485 23366 11497 23418
rect 11549 23366 11561 23418
rect 11613 23366 11625 23418
rect 11677 23366 18315 23418
rect 18367 23366 18379 23418
rect 18431 23366 18443 23418
rect 18495 23366 18507 23418
rect 18559 23366 18571 23418
rect 18623 23366 25261 23418
rect 25313 23366 25325 23418
rect 25377 23366 25389 23418
rect 25441 23366 25453 23418
rect 25505 23366 25517 23418
rect 25569 23366 28888 23418
rect 1104 23344 28888 23366
rect 1581 23239 1639 23245
rect 1581 23205 1593 23239
rect 1627 23236 1639 23239
rect 4246 23236 4252 23248
rect 1627 23208 4252 23236
rect 1627 23205 1639 23208
rect 1581 23199 1639 23205
rect 4246 23196 4252 23208
rect 4304 23196 4310 23248
rect 934 23060 940 23112
rect 992 23100 998 23112
rect 1397 23103 1455 23109
rect 1397 23100 1409 23103
rect 992 23072 1409 23100
rect 992 23060 998 23072
rect 1397 23069 1409 23072
rect 1443 23069 1455 23103
rect 1397 23063 1455 23069
rect 1673 23103 1731 23109
rect 1673 23069 1685 23103
rect 1719 23069 1731 23103
rect 1673 23063 1731 23069
rect 27157 23103 27215 23109
rect 27157 23069 27169 23103
rect 27203 23069 27215 23103
rect 27157 23063 27215 23069
rect 1026 22992 1032 23044
rect 1084 23032 1090 23044
rect 1688 23032 1716 23063
rect 1084 23004 1716 23032
rect 1084 22992 1090 23004
rect 1854 22924 1860 22976
rect 1912 22924 1918 22976
rect 16022 22924 16028 22976
rect 16080 22964 16086 22976
rect 26973 22967 27031 22973
rect 26973 22964 26985 22967
rect 16080 22936 26985 22964
rect 16080 22924 16086 22936
rect 26973 22933 26985 22936
rect 27019 22964 27031 22967
rect 27172 22964 27200 23063
rect 28350 22992 28356 23044
rect 28408 22992 28414 23044
rect 27019 22936 27200 22964
rect 27019 22933 27031 22936
rect 26973 22927 27031 22933
rect 1104 22874 29048 22896
rect 1104 22822 7896 22874
rect 7948 22822 7960 22874
rect 8012 22822 8024 22874
rect 8076 22822 8088 22874
rect 8140 22822 8152 22874
rect 8204 22822 14842 22874
rect 14894 22822 14906 22874
rect 14958 22822 14970 22874
rect 15022 22822 15034 22874
rect 15086 22822 15098 22874
rect 15150 22822 21788 22874
rect 21840 22822 21852 22874
rect 21904 22822 21916 22874
rect 21968 22822 21980 22874
rect 22032 22822 22044 22874
rect 22096 22822 28734 22874
rect 28786 22822 28798 22874
rect 28850 22822 28862 22874
rect 28914 22822 28926 22874
rect 28978 22822 28990 22874
rect 29042 22822 29048 22874
rect 1104 22800 29048 22822
rect 1026 22584 1032 22636
rect 1084 22624 1090 22636
rect 1397 22627 1455 22633
rect 1397 22624 1409 22627
rect 1084 22596 1409 22624
rect 1084 22584 1090 22596
rect 1397 22593 1409 22596
rect 1443 22593 1455 22627
rect 1397 22587 1455 22593
rect 1673 22627 1731 22633
rect 1673 22593 1685 22627
rect 1719 22593 1731 22627
rect 1673 22587 1731 22593
rect 934 22516 940 22568
rect 992 22556 998 22568
rect 1688 22556 1716 22587
rect 992 22528 1716 22556
rect 992 22516 998 22528
rect 2038 22488 2044 22500
rect 1596 22460 2044 22488
rect 1596 22429 1624 22460
rect 2038 22448 2044 22460
rect 2096 22448 2102 22500
rect 1581 22423 1639 22429
rect 1581 22389 1593 22423
rect 1627 22389 1639 22423
rect 1581 22383 1639 22389
rect 1857 22423 1915 22429
rect 1857 22389 1869 22423
rect 1903 22420 1915 22423
rect 10226 22420 10232 22432
rect 1903 22392 10232 22420
rect 1903 22389 1915 22392
rect 1857 22383 1915 22389
rect 10226 22380 10232 22392
rect 10284 22380 10290 22432
rect 1104 22330 28888 22352
rect 1104 22278 4423 22330
rect 4475 22278 4487 22330
rect 4539 22278 4551 22330
rect 4603 22278 4615 22330
rect 4667 22278 4679 22330
rect 4731 22278 11369 22330
rect 11421 22278 11433 22330
rect 11485 22278 11497 22330
rect 11549 22278 11561 22330
rect 11613 22278 11625 22330
rect 11677 22278 18315 22330
rect 18367 22278 18379 22330
rect 18431 22278 18443 22330
rect 18495 22278 18507 22330
rect 18559 22278 18571 22330
rect 18623 22278 25261 22330
rect 25313 22278 25325 22330
rect 25377 22278 25389 22330
rect 25441 22278 25453 22330
rect 25505 22278 25517 22330
rect 25569 22278 28888 22330
rect 1104 22256 28888 22278
rect 28353 22083 28411 22089
rect 28353 22049 28365 22083
rect 28399 22080 28411 22083
rect 28810 22080 28816 22092
rect 28399 22052 28816 22080
rect 28399 22049 28411 22052
rect 28353 22043 28411 22049
rect 28810 22040 28816 22052
rect 28868 22040 28874 22092
rect 934 21972 940 22024
rect 992 22012 998 22024
rect 1397 22015 1455 22021
rect 1397 22012 1409 22015
rect 992 21984 1409 22012
rect 992 21972 998 21984
rect 1397 21981 1409 21984
rect 1443 21981 1455 22015
rect 1397 21975 1455 21981
rect 1673 22015 1731 22021
rect 1673 21981 1685 22015
rect 1719 21981 1731 22015
rect 1673 21975 1731 21981
rect 27157 22015 27215 22021
rect 27157 21981 27169 22015
rect 27203 21981 27215 22015
rect 27157 21975 27215 21981
rect 1026 21904 1032 21956
rect 1084 21944 1090 21956
rect 1688 21944 1716 21975
rect 9214 21944 9220 21956
rect 1084 21916 1716 21944
rect 1780 21916 9220 21944
rect 1084 21904 1090 21916
rect 1581 21879 1639 21885
rect 1581 21845 1593 21879
rect 1627 21876 1639 21879
rect 1780 21876 1808 21916
rect 9214 21904 9220 21916
rect 9272 21904 9278 21956
rect 1627 21848 1808 21876
rect 1857 21879 1915 21885
rect 1627 21845 1639 21848
rect 1581 21839 1639 21845
rect 1857 21845 1869 21879
rect 1903 21876 1915 21879
rect 9674 21876 9680 21888
rect 1903 21848 9680 21876
rect 1903 21845 1915 21848
rect 1857 21839 1915 21845
rect 9674 21836 9680 21848
rect 9732 21836 9738 21888
rect 14642 21836 14648 21888
rect 14700 21876 14706 21888
rect 26973 21879 27031 21885
rect 26973 21876 26985 21879
rect 14700 21848 26985 21876
rect 14700 21836 14706 21848
rect 26973 21845 26985 21848
rect 27019 21876 27031 21879
rect 27172 21876 27200 21975
rect 27019 21848 27200 21876
rect 27019 21845 27031 21848
rect 26973 21839 27031 21845
rect 1104 21786 29048 21808
rect 1104 21734 7896 21786
rect 7948 21734 7960 21786
rect 8012 21734 8024 21786
rect 8076 21734 8088 21786
rect 8140 21734 8152 21786
rect 8204 21734 14842 21786
rect 14894 21734 14906 21786
rect 14958 21734 14970 21786
rect 15022 21734 15034 21786
rect 15086 21734 15098 21786
rect 15150 21734 21788 21786
rect 21840 21734 21852 21786
rect 21904 21734 21916 21786
rect 21968 21734 21980 21786
rect 22032 21734 22044 21786
rect 22096 21734 28734 21786
rect 28786 21734 28798 21786
rect 28850 21734 28862 21786
rect 28914 21734 28926 21786
rect 28978 21734 28990 21786
rect 29042 21734 29048 21786
rect 1104 21712 29048 21734
rect 1026 21496 1032 21548
rect 1084 21536 1090 21548
rect 1397 21539 1455 21545
rect 1397 21536 1409 21539
rect 1084 21508 1409 21536
rect 1084 21496 1090 21508
rect 1397 21505 1409 21508
rect 1443 21505 1455 21539
rect 1397 21499 1455 21505
rect 1673 21539 1731 21545
rect 1673 21505 1685 21539
rect 1719 21505 1731 21539
rect 1673 21499 1731 21505
rect 934 21428 940 21480
rect 992 21468 998 21480
rect 1688 21468 1716 21499
rect 15746 21496 15752 21548
rect 15804 21536 15810 21548
rect 26697 21539 26755 21545
rect 26697 21536 26709 21539
rect 15804 21508 26709 21536
rect 15804 21496 15810 21508
rect 26697 21505 26709 21508
rect 26743 21536 26755 21539
rect 27157 21539 27215 21545
rect 27157 21536 27169 21539
rect 26743 21508 27169 21536
rect 26743 21505 26755 21508
rect 26697 21499 26755 21505
rect 27157 21505 27169 21508
rect 27203 21505 27215 21539
rect 27157 21499 27215 21505
rect 992 21440 1716 21468
rect 992 21428 998 21440
rect 28350 21428 28356 21480
rect 28408 21428 28414 21480
rect 1581 21403 1639 21409
rect 1581 21369 1593 21403
rect 1627 21400 1639 21403
rect 7466 21400 7472 21412
rect 1627 21372 7472 21400
rect 1627 21369 1639 21372
rect 1581 21363 1639 21369
rect 7466 21360 7472 21372
rect 7524 21360 7530 21412
rect 1857 21335 1915 21341
rect 1857 21301 1869 21335
rect 1903 21332 1915 21335
rect 8386 21332 8392 21344
rect 1903 21304 8392 21332
rect 1903 21301 1915 21304
rect 1857 21295 1915 21301
rect 8386 21292 8392 21304
rect 8444 21292 8450 21344
rect 1104 21242 28888 21264
rect 1104 21190 4423 21242
rect 4475 21190 4487 21242
rect 4539 21190 4551 21242
rect 4603 21190 4615 21242
rect 4667 21190 4679 21242
rect 4731 21190 11369 21242
rect 11421 21190 11433 21242
rect 11485 21190 11497 21242
rect 11549 21190 11561 21242
rect 11613 21190 11625 21242
rect 11677 21190 18315 21242
rect 18367 21190 18379 21242
rect 18431 21190 18443 21242
rect 18495 21190 18507 21242
rect 18559 21190 18571 21242
rect 18623 21190 25261 21242
rect 25313 21190 25325 21242
rect 25377 21190 25389 21242
rect 25441 21190 25453 21242
rect 25505 21190 25517 21242
rect 25569 21190 28888 21242
rect 1104 21168 28888 21190
rect 1581 21063 1639 21069
rect 1581 21029 1593 21063
rect 1627 21060 1639 21063
rect 4062 21060 4068 21072
rect 1627 21032 4068 21060
rect 1627 21029 1639 21032
rect 1581 21023 1639 21029
rect 4062 21020 4068 21032
rect 4120 21020 4126 21072
rect 1394 20884 1400 20936
rect 1452 20884 1458 20936
rect 1673 20927 1731 20933
rect 1673 20893 1685 20927
rect 1719 20893 1731 20927
rect 1673 20887 1731 20893
rect 934 20816 940 20868
rect 992 20856 998 20868
rect 1688 20856 1716 20887
rect 992 20828 1716 20856
rect 992 20816 998 20828
rect 1857 20791 1915 20797
rect 1857 20757 1869 20791
rect 1903 20788 1915 20791
rect 7650 20788 7656 20800
rect 1903 20760 7656 20788
rect 1903 20757 1915 20760
rect 1857 20751 1915 20757
rect 7650 20748 7656 20760
rect 7708 20748 7714 20800
rect 1104 20698 29048 20720
rect 1104 20646 7896 20698
rect 7948 20646 7960 20698
rect 8012 20646 8024 20698
rect 8076 20646 8088 20698
rect 8140 20646 8152 20698
rect 8204 20646 14842 20698
rect 14894 20646 14906 20698
rect 14958 20646 14970 20698
rect 15022 20646 15034 20698
rect 15086 20646 15098 20698
rect 15150 20646 21788 20698
rect 21840 20646 21852 20698
rect 21904 20646 21916 20698
rect 21968 20646 21980 20698
rect 22032 20646 22044 20698
rect 22096 20646 28734 20698
rect 28786 20646 28798 20698
rect 28850 20646 28862 20698
rect 28914 20646 28926 20698
rect 28978 20646 28990 20698
rect 29042 20646 29048 20698
rect 1104 20624 29048 20646
rect 934 20408 940 20460
rect 992 20448 998 20460
rect 1397 20451 1455 20457
rect 1397 20448 1409 20451
rect 992 20420 1409 20448
rect 992 20408 998 20420
rect 1397 20417 1409 20420
rect 1443 20417 1455 20451
rect 1397 20411 1455 20417
rect 1673 20451 1731 20457
rect 1673 20417 1685 20451
rect 1719 20417 1731 20451
rect 27157 20451 27215 20457
rect 27157 20448 27169 20451
rect 1673 20411 1731 20417
rect 26712 20420 27169 20448
rect 1026 20340 1032 20392
rect 1084 20380 1090 20392
rect 1688 20380 1716 20411
rect 1084 20352 1716 20380
rect 1084 20340 1090 20352
rect 1578 20204 1584 20256
rect 1636 20204 1642 20256
rect 1857 20247 1915 20253
rect 1857 20213 1869 20247
rect 1903 20244 1915 20247
rect 5534 20244 5540 20256
rect 1903 20216 5540 20244
rect 1903 20213 1915 20216
rect 1857 20207 1915 20213
rect 5534 20204 5540 20216
rect 5592 20204 5598 20256
rect 16206 20204 16212 20256
rect 16264 20244 16270 20256
rect 26712 20253 26740 20420
rect 27157 20417 27169 20420
rect 27203 20417 27215 20451
rect 27157 20411 27215 20417
rect 28350 20340 28356 20392
rect 28408 20340 28414 20392
rect 26697 20247 26755 20253
rect 26697 20244 26709 20247
rect 16264 20216 26709 20244
rect 16264 20204 16270 20216
rect 26697 20213 26709 20216
rect 26743 20213 26755 20247
rect 26697 20207 26755 20213
rect 1104 20154 28888 20176
rect 1104 20102 4423 20154
rect 4475 20102 4487 20154
rect 4539 20102 4551 20154
rect 4603 20102 4615 20154
rect 4667 20102 4679 20154
rect 4731 20102 11369 20154
rect 11421 20102 11433 20154
rect 11485 20102 11497 20154
rect 11549 20102 11561 20154
rect 11613 20102 11625 20154
rect 11677 20102 18315 20154
rect 18367 20102 18379 20154
rect 18431 20102 18443 20154
rect 18495 20102 18507 20154
rect 18559 20102 18571 20154
rect 18623 20102 25261 20154
rect 25313 20102 25325 20154
rect 25377 20102 25389 20154
rect 25441 20102 25453 20154
rect 25505 20102 25517 20154
rect 25569 20102 28888 20154
rect 1104 20080 28888 20102
rect 1581 19975 1639 19981
rect 1581 19941 1593 19975
rect 1627 19972 1639 19975
rect 5626 19972 5632 19984
rect 1627 19944 5632 19972
rect 1627 19941 1639 19944
rect 1581 19935 1639 19941
rect 5626 19932 5632 19944
rect 5684 19932 5690 19984
rect 934 19796 940 19848
rect 992 19836 998 19848
rect 1397 19839 1455 19845
rect 1397 19836 1409 19839
rect 992 19808 1409 19836
rect 992 19796 998 19808
rect 1397 19805 1409 19808
rect 1443 19805 1455 19839
rect 1397 19799 1455 19805
rect 1673 19839 1731 19845
rect 1673 19805 1685 19839
rect 1719 19805 1731 19839
rect 1673 19799 1731 19805
rect 27157 19839 27215 19845
rect 27157 19805 27169 19839
rect 27203 19805 27215 19839
rect 27157 19799 27215 19805
rect 1026 19728 1032 19780
rect 1084 19768 1090 19780
rect 1688 19768 1716 19799
rect 1084 19740 1716 19768
rect 1084 19728 1090 19740
rect 1854 19660 1860 19712
rect 1912 19660 1918 19712
rect 10778 19660 10784 19712
rect 10836 19700 10842 19712
rect 26973 19703 27031 19709
rect 26973 19700 26985 19703
rect 10836 19672 26985 19700
rect 10836 19660 10842 19672
rect 26973 19669 26985 19672
rect 27019 19700 27031 19703
rect 27172 19700 27200 19799
rect 28350 19728 28356 19780
rect 28408 19728 28414 19780
rect 27019 19672 27200 19700
rect 27019 19669 27031 19672
rect 26973 19663 27031 19669
rect 1104 19610 29048 19632
rect 1104 19558 7896 19610
rect 7948 19558 7960 19610
rect 8012 19558 8024 19610
rect 8076 19558 8088 19610
rect 8140 19558 8152 19610
rect 8204 19558 14842 19610
rect 14894 19558 14906 19610
rect 14958 19558 14970 19610
rect 15022 19558 15034 19610
rect 15086 19558 15098 19610
rect 15150 19558 21788 19610
rect 21840 19558 21852 19610
rect 21904 19558 21916 19610
rect 21968 19558 21980 19610
rect 22032 19558 22044 19610
rect 22096 19558 28734 19610
rect 28786 19558 28798 19610
rect 28850 19558 28862 19610
rect 28914 19558 28926 19610
rect 28978 19558 28990 19610
rect 29042 19558 29048 19610
rect 1104 19536 29048 19558
rect 1581 19499 1639 19505
rect 1581 19465 1593 19499
rect 1627 19465 1639 19499
rect 1581 19459 1639 19465
rect 1857 19499 1915 19505
rect 1857 19465 1869 19499
rect 1903 19496 1915 19499
rect 3602 19496 3608 19508
rect 1903 19468 3608 19496
rect 1903 19465 1915 19468
rect 1857 19459 1915 19465
rect 1596 19428 1624 19459
rect 3602 19456 3608 19468
rect 3660 19456 3666 19508
rect 3970 19428 3976 19440
rect 1596 19400 3976 19428
rect 3970 19388 3976 19400
rect 4028 19388 4034 19440
rect 1394 19320 1400 19372
rect 1452 19320 1458 19372
rect 1670 19320 1676 19372
rect 1728 19320 1734 19372
rect 1104 19066 28888 19088
rect 1104 19014 4423 19066
rect 4475 19014 4487 19066
rect 4539 19014 4551 19066
rect 4603 19014 4615 19066
rect 4667 19014 4679 19066
rect 4731 19014 11369 19066
rect 11421 19014 11433 19066
rect 11485 19014 11497 19066
rect 11549 19014 11561 19066
rect 11613 19014 11625 19066
rect 11677 19014 18315 19066
rect 18367 19014 18379 19066
rect 18431 19014 18443 19066
rect 18495 19014 18507 19066
rect 18559 19014 18571 19066
rect 18623 19014 25261 19066
rect 25313 19014 25325 19066
rect 25377 19014 25389 19066
rect 25441 19014 25453 19066
rect 25505 19014 25517 19066
rect 25569 19014 28888 19066
rect 1104 18992 28888 19014
rect 12802 18912 12808 18964
rect 12860 18912 12866 18964
rect 1581 18887 1639 18893
rect 1581 18853 1593 18887
rect 1627 18884 1639 18887
rect 3326 18884 3332 18896
rect 1627 18856 3332 18884
rect 1627 18853 1639 18856
rect 1581 18847 1639 18853
rect 3326 18844 3332 18856
rect 3384 18844 3390 18896
rect 28353 18819 28411 18825
rect 28353 18785 28365 18819
rect 28399 18816 28411 18819
rect 28810 18816 28816 18828
rect 28399 18788 28816 18816
rect 28399 18785 28411 18788
rect 28353 18779 28411 18785
rect 28810 18776 28816 18788
rect 28868 18776 28874 18828
rect 934 18708 940 18760
rect 992 18748 998 18760
rect 1397 18751 1455 18757
rect 1397 18748 1409 18751
rect 992 18720 1409 18748
rect 992 18708 998 18720
rect 1397 18717 1409 18720
rect 1443 18717 1455 18751
rect 1397 18711 1455 18717
rect 1673 18751 1731 18757
rect 1673 18717 1685 18751
rect 1719 18717 1731 18751
rect 1673 18711 1731 18717
rect 27157 18751 27215 18757
rect 27157 18717 27169 18751
rect 27203 18717 27215 18751
rect 27157 18711 27215 18717
rect 1026 18640 1032 18692
rect 1084 18680 1090 18692
rect 1688 18680 1716 18711
rect 1084 18652 1716 18680
rect 1084 18640 1090 18652
rect 1857 18615 1915 18621
rect 1857 18581 1869 18615
rect 1903 18612 1915 18615
rect 3786 18612 3792 18624
rect 1903 18584 3792 18612
rect 1903 18581 1915 18584
rect 1857 18575 1915 18581
rect 3786 18572 3792 18584
rect 3844 18572 3850 18624
rect 17770 18572 17776 18624
rect 17828 18612 17834 18624
rect 26973 18615 27031 18621
rect 26973 18612 26985 18615
rect 17828 18584 26985 18612
rect 17828 18572 17834 18584
rect 26973 18581 26985 18584
rect 27019 18612 27031 18615
rect 27172 18612 27200 18711
rect 27019 18584 27200 18612
rect 27019 18581 27031 18584
rect 26973 18575 27031 18581
rect 1104 18522 29048 18544
rect 1104 18470 7896 18522
rect 7948 18470 7960 18522
rect 8012 18470 8024 18522
rect 8076 18470 8088 18522
rect 8140 18470 8152 18522
rect 8204 18470 14842 18522
rect 14894 18470 14906 18522
rect 14958 18470 14970 18522
rect 15022 18470 15034 18522
rect 15086 18470 15098 18522
rect 15150 18470 21788 18522
rect 21840 18470 21852 18522
rect 21904 18470 21916 18522
rect 21968 18470 21980 18522
rect 22032 18470 22044 18522
rect 22096 18470 28734 18522
rect 28786 18470 28798 18522
rect 28850 18470 28862 18522
rect 28914 18470 28926 18522
rect 28978 18470 28990 18522
rect 29042 18470 29048 18522
rect 1104 18448 29048 18470
rect 12253 18411 12311 18417
rect 12253 18377 12265 18411
rect 12299 18408 12311 18411
rect 12802 18408 12808 18420
rect 12299 18380 12808 18408
rect 12299 18377 12311 18380
rect 12253 18371 12311 18377
rect 12802 18368 12808 18380
rect 12860 18408 12866 18420
rect 13722 18408 13728 18420
rect 12860 18380 13728 18408
rect 12860 18368 12866 18380
rect 13722 18368 13728 18380
rect 13780 18368 13786 18420
rect 8294 18300 8300 18352
rect 8352 18340 8358 18352
rect 26697 18343 26755 18349
rect 26697 18340 26709 18343
rect 8352 18312 26709 18340
rect 8352 18300 8358 18312
rect 26697 18309 26709 18312
rect 26743 18309 26755 18343
rect 26697 18303 26755 18309
rect 1394 18232 1400 18284
rect 1452 18232 1458 18284
rect 1673 18275 1731 18281
rect 1673 18241 1685 18275
rect 1719 18241 1731 18275
rect 1673 18235 1731 18241
rect 934 18164 940 18216
rect 992 18204 998 18216
rect 1688 18204 1716 18235
rect 9214 18232 9220 18284
rect 9272 18232 9278 18284
rect 9398 18232 9404 18284
rect 9456 18232 9462 18284
rect 9674 18232 9680 18284
rect 9732 18232 9738 18284
rect 9858 18232 9864 18284
rect 9916 18232 9922 18284
rect 10594 18232 10600 18284
rect 10652 18272 10658 18284
rect 12161 18275 12219 18281
rect 12161 18272 12173 18275
rect 10652 18244 12173 18272
rect 10652 18232 10658 18244
rect 12161 18241 12173 18244
rect 12207 18241 12219 18275
rect 26712 18272 26740 18303
rect 27157 18275 27215 18281
rect 27157 18272 27169 18275
rect 26712 18244 27169 18272
rect 12161 18235 12219 18241
rect 27157 18241 27169 18244
rect 27203 18241 27215 18275
rect 27157 18235 27215 18241
rect 992 18176 1716 18204
rect 992 18164 998 18176
rect 4246 18164 4252 18216
rect 4304 18204 4310 18216
rect 10134 18204 10140 18216
rect 4304 18176 10140 18204
rect 4304 18164 4310 18176
rect 10134 18164 10140 18176
rect 10192 18164 10198 18216
rect 10502 18164 10508 18216
rect 10560 18204 10566 18216
rect 11977 18207 12035 18213
rect 11977 18204 11989 18207
rect 10560 18176 11989 18204
rect 10560 18164 10566 18176
rect 11977 18173 11989 18176
rect 12023 18173 12035 18207
rect 13265 18207 13323 18213
rect 13265 18204 13277 18207
rect 11977 18167 12035 18173
rect 12636 18176 13277 18204
rect 3418 18136 3424 18148
rect 1596 18108 3424 18136
rect 1596 18077 1624 18108
rect 3418 18096 3424 18108
rect 3476 18096 3482 18148
rect 9585 18139 9643 18145
rect 9585 18105 9597 18139
rect 9631 18136 9643 18139
rect 10870 18136 10876 18148
rect 9631 18108 10876 18136
rect 9631 18105 9643 18108
rect 9585 18099 9643 18105
rect 10870 18096 10876 18108
rect 10928 18096 10934 18148
rect 12636 18145 12664 18176
rect 13265 18173 13277 18176
rect 13311 18173 13323 18207
rect 13265 18167 13323 18173
rect 28350 18164 28356 18216
rect 28408 18164 28414 18216
rect 12621 18139 12679 18145
rect 12621 18105 12633 18139
rect 12667 18105 12679 18139
rect 12621 18099 12679 18105
rect 1581 18071 1639 18077
rect 1581 18037 1593 18071
rect 1627 18037 1639 18071
rect 1581 18031 1639 18037
rect 1857 18071 1915 18077
rect 1857 18037 1869 18071
rect 1903 18068 1915 18071
rect 4154 18068 4160 18080
rect 1903 18040 4160 18068
rect 1903 18037 1915 18040
rect 1857 18031 1915 18037
rect 4154 18028 4160 18040
rect 4212 18028 4218 18080
rect 10042 18028 10048 18080
rect 10100 18028 10106 18080
rect 12710 18028 12716 18080
rect 12768 18028 12774 18080
rect 1104 17978 28888 18000
rect 1104 17926 4423 17978
rect 4475 17926 4487 17978
rect 4539 17926 4551 17978
rect 4603 17926 4615 17978
rect 4667 17926 4679 17978
rect 4731 17926 11369 17978
rect 11421 17926 11433 17978
rect 11485 17926 11497 17978
rect 11549 17926 11561 17978
rect 11613 17926 11625 17978
rect 11677 17926 18315 17978
rect 18367 17926 18379 17978
rect 18431 17926 18443 17978
rect 18495 17926 18507 17978
rect 18559 17926 18571 17978
rect 18623 17926 25261 17978
rect 25313 17926 25325 17978
rect 25377 17926 25389 17978
rect 25441 17926 25453 17978
rect 25505 17926 25517 17978
rect 25569 17926 28888 17978
rect 1104 17904 28888 17926
rect 10594 17824 10600 17876
rect 10652 17824 10658 17876
rect 1581 17799 1639 17805
rect 1581 17765 1593 17799
rect 1627 17796 1639 17799
rect 3694 17796 3700 17808
rect 1627 17768 3700 17796
rect 1627 17765 1639 17768
rect 1581 17759 1639 17765
rect 3694 17756 3700 17768
rect 3752 17756 3758 17808
rect 9217 17799 9275 17805
rect 9217 17765 9229 17799
rect 9263 17796 9275 17799
rect 9766 17796 9772 17808
rect 9263 17768 9772 17796
rect 9263 17765 9275 17768
rect 9217 17759 9275 17765
rect 9766 17756 9772 17768
rect 9824 17796 9830 17808
rect 10778 17796 10784 17808
rect 9824 17768 10784 17796
rect 9824 17756 9830 17768
rect 10778 17756 10784 17768
rect 10836 17756 10842 17808
rect 10226 17688 10232 17740
rect 10284 17688 10290 17740
rect 11425 17731 11483 17737
rect 11425 17697 11437 17731
rect 11471 17728 11483 17731
rect 11698 17728 11704 17740
rect 11471 17700 11704 17728
rect 11471 17697 11483 17700
rect 11425 17691 11483 17697
rect 11698 17688 11704 17700
rect 11756 17688 11762 17740
rect 11790 17688 11796 17740
rect 11848 17728 11854 17740
rect 13449 17731 13507 17737
rect 13449 17728 13461 17731
rect 11848 17700 13461 17728
rect 11848 17688 11854 17700
rect 13449 17697 13461 17700
rect 13495 17728 13507 17731
rect 16022 17728 16028 17740
rect 13495 17700 16028 17728
rect 13495 17697 13507 17700
rect 13449 17691 13507 17697
rect 16022 17688 16028 17700
rect 16080 17688 16086 17740
rect 1026 17620 1032 17672
rect 1084 17660 1090 17672
rect 1397 17663 1455 17669
rect 1397 17660 1409 17663
rect 1084 17632 1409 17660
rect 1084 17620 1090 17632
rect 1397 17629 1409 17632
rect 1443 17629 1455 17663
rect 1397 17623 1455 17629
rect 1673 17663 1731 17669
rect 1673 17629 1685 17663
rect 1719 17629 1731 17663
rect 1673 17623 1731 17629
rect 934 17552 940 17604
rect 992 17592 998 17604
rect 1688 17592 1716 17623
rect 9858 17620 9864 17672
rect 9916 17620 9922 17672
rect 10410 17620 10416 17672
rect 10468 17620 10474 17672
rect 10686 17620 10692 17672
rect 10744 17620 10750 17672
rect 992 17564 1716 17592
rect 11333 17595 11391 17601
rect 992 17552 998 17564
rect 11333 17561 11345 17595
rect 11379 17592 11391 17595
rect 11701 17595 11759 17601
rect 11701 17592 11713 17595
rect 11379 17564 11713 17592
rect 11379 17561 11391 17564
rect 11333 17555 11391 17561
rect 11701 17561 11713 17564
rect 11747 17561 11759 17595
rect 13170 17592 13176 17604
rect 12926 17564 13176 17592
rect 11701 17555 11759 17561
rect 13170 17552 13176 17564
rect 13228 17552 13234 17604
rect 1857 17527 1915 17533
rect 1857 17493 1869 17527
rect 1903 17524 1915 17527
rect 3510 17524 3516 17536
rect 1903 17496 3516 17524
rect 1903 17493 1915 17496
rect 1857 17487 1915 17493
rect 3510 17484 3516 17496
rect 3568 17484 3574 17536
rect 8481 17527 8539 17533
rect 8481 17493 8493 17527
rect 8527 17524 8539 17527
rect 8754 17524 8760 17536
rect 8527 17496 8760 17524
rect 8527 17493 8539 17496
rect 8481 17487 8539 17493
rect 8754 17484 8760 17496
rect 8812 17484 8818 17536
rect 9306 17484 9312 17536
rect 9364 17484 9370 17536
rect 1104 17434 29048 17456
rect 1104 17382 7896 17434
rect 7948 17382 7960 17434
rect 8012 17382 8024 17434
rect 8076 17382 8088 17434
rect 8140 17382 8152 17434
rect 8204 17382 14842 17434
rect 14894 17382 14906 17434
rect 14958 17382 14970 17434
rect 15022 17382 15034 17434
rect 15086 17382 15098 17434
rect 15150 17382 21788 17434
rect 21840 17382 21852 17434
rect 21904 17382 21916 17434
rect 21968 17382 21980 17434
rect 22032 17382 22044 17434
rect 22096 17382 28734 17434
rect 28786 17382 28798 17434
rect 28850 17382 28862 17434
rect 28914 17382 28926 17434
rect 28978 17382 28990 17434
rect 29042 17382 29048 17434
rect 1104 17360 29048 17382
rect 1581 17323 1639 17329
rect 1581 17289 1593 17323
rect 1627 17320 1639 17323
rect 5258 17320 5264 17332
rect 1627 17292 5264 17320
rect 1627 17289 1639 17292
rect 1581 17283 1639 17289
rect 5258 17280 5264 17292
rect 5316 17280 5322 17332
rect 8846 17280 8852 17332
rect 8904 17280 8910 17332
rect 9309 17323 9367 17329
rect 9309 17289 9321 17323
rect 9355 17320 9367 17323
rect 9858 17320 9864 17332
rect 9355 17292 9864 17320
rect 9355 17289 9367 17292
rect 9309 17283 9367 17289
rect 9858 17280 9864 17292
rect 9916 17280 9922 17332
rect 10042 17280 10048 17332
rect 10100 17280 10106 17332
rect 10505 17323 10563 17329
rect 10505 17289 10517 17323
rect 10551 17320 10563 17323
rect 10686 17320 10692 17332
rect 10551 17292 10692 17320
rect 10551 17289 10563 17292
rect 10505 17283 10563 17289
rect 10686 17280 10692 17292
rect 10744 17280 10750 17332
rect 10870 17280 10876 17332
rect 10928 17280 10934 17332
rect 11790 17280 11796 17332
rect 11848 17280 11854 17332
rect 12710 17320 12716 17332
rect 11992 17292 12716 17320
rect 1854 17212 1860 17264
rect 1912 17252 1918 17264
rect 8864 17252 8892 17280
rect 1912 17224 8892 17252
rect 9677 17255 9735 17261
rect 1912 17212 1918 17224
rect 9677 17221 9689 17255
rect 9723 17252 9735 17255
rect 10137 17255 10195 17261
rect 10137 17252 10149 17255
rect 9723 17224 10149 17252
rect 9723 17221 9735 17224
rect 9677 17215 9735 17221
rect 10137 17221 10149 17224
rect 10183 17252 10195 17255
rect 11808 17252 11836 17280
rect 11992 17261 12020 17292
rect 12710 17280 12716 17292
rect 12768 17280 12774 17332
rect 10183 17224 11836 17252
rect 11977 17255 12035 17261
rect 10183 17221 10195 17224
rect 10137 17215 10195 17221
rect 11977 17221 11989 17255
rect 12023 17221 12035 17255
rect 14645 17255 14703 17261
rect 14645 17252 14657 17255
rect 13202 17224 14657 17252
rect 11977 17215 12035 17221
rect 14645 17221 14657 17224
rect 14691 17221 14703 17255
rect 14645 17215 14703 17221
rect 934 17144 940 17196
rect 992 17184 998 17196
rect 1397 17187 1455 17193
rect 1397 17184 1409 17187
rect 992 17156 1409 17184
rect 992 17144 998 17156
rect 1397 17153 1409 17156
rect 1443 17153 1455 17187
rect 1397 17147 1455 17153
rect 1673 17187 1731 17193
rect 1673 17153 1685 17187
rect 1719 17153 1731 17187
rect 1673 17147 1731 17153
rect 1026 17076 1032 17128
rect 1084 17116 1090 17128
rect 1688 17116 1716 17147
rect 5534 17144 5540 17196
rect 5592 17184 5598 17196
rect 5592 17156 7328 17184
rect 5592 17144 5598 17156
rect 1084 17088 1716 17116
rect 1084 17076 1090 17088
rect 7190 17076 7196 17128
rect 7248 17076 7254 17128
rect 7300 17116 7328 17156
rect 7374 17144 7380 17196
rect 7432 17184 7438 17196
rect 7561 17187 7619 17193
rect 7561 17184 7573 17187
rect 7432 17156 7573 17184
rect 7432 17144 7438 17156
rect 7561 17153 7573 17156
rect 7607 17153 7619 17187
rect 7561 17147 7619 17153
rect 7650 17144 7656 17196
rect 7708 17184 7714 17196
rect 8113 17187 8171 17193
rect 8113 17184 8125 17187
rect 7708 17156 8125 17184
rect 7708 17144 7714 17156
rect 8113 17153 8125 17156
rect 8159 17153 8171 17187
rect 8113 17147 8171 17153
rect 8297 17187 8355 17193
rect 8297 17153 8309 17187
rect 8343 17153 8355 17187
rect 8297 17147 8355 17153
rect 8481 17187 8539 17193
rect 8481 17153 8493 17187
rect 8527 17184 8539 17187
rect 8849 17187 8907 17193
rect 8849 17184 8861 17187
rect 8527 17156 8861 17184
rect 8527 17153 8539 17156
rect 8481 17147 8539 17153
rect 8849 17153 8861 17156
rect 8895 17153 8907 17187
rect 8849 17147 8907 17153
rect 8941 17187 8999 17193
rect 8941 17153 8953 17187
rect 8987 17184 8999 17187
rect 9766 17184 9772 17196
rect 8987 17156 9772 17184
rect 8987 17153 8999 17156
rect 8941 17147 8999 17153
rect 7745 17119 7803 17125
rect 7745 17116 7757 17119
rect 7300 17088 7757 17116
rect 7745 17085 7757 17088
rect 7791 17085 7803 17119
rect 7745 17079 7803 17085
rect 1302 17008 1308 17060
rect 1360 17048 1366 17060
rect 1360 17020 1900 17048
rect 1360 17008 1366 17020
rect 1872 16989 1900 17020
rect 7558 17008 7564 17060
rect 7616 17048 7622 17060
rect 8312 17048 8340 17147
rect 9766 17144 9772 17156
rect 9824 17144 9830 17196
rect 10962 17144 10968 17196
rect 11020 17144 11026 17196
rect 13722 17144 13728 17196
rect 13780 17144 13786 17196
rect 14734 17144 14740 17196
rect 14792 17184 14798 17196
rect 15013 17187 15071 17193
rect 15013 17184 15025 17187
rect 14792 17156 15025 17184
rect 14792 17144 14798 17156
rect 15013 17153 15025 17156
rect 15059 17153 15071 17187
rect 15013 17147 15071 17153
rect 16574 17144 16580 17196
rect 16632 17184 16638 17196
rect 27157 17187 27215 17193
rect 27157 17184 27169 17187
rect 16632 17156 27169 17184
rect 16632 17144 16638 17156
rect 27157 17153 27169 17156
rect 27203 17153 27215 17187
rect 27157 17147 27215 17153
rect 8754 17076 8760 17128
rect 8812 17076 8818 17128
rect 9953 17119 10011 17125
rect 9953 17085 9965 17119
rect 9999 17116 10011 17119
rect 10502 17116 10508 17128
rect 9999 17088 10508 17116
rect 9999 17085 10011 17088
rect 9953 17079 10011 17085
rect 7616 17020 8340 17048
rect 7616 17008 7622 17020
rect 1857 16983 1915 16989
rect 1857 16949 1869 16983
rect 1903 16949 1915 16983
rect 1857 16943 1915 16949
rect 6454 16940 6460 16992
rect 6512 16980 6518 16992
rect 6641 16983 6699 16989
rect 6641 16980 6653 16983
rect 6512 16952 6653 16980
rect 6512 16940 6518 16952
rect 6641 16949 6653 16952
rect 6687 16949 6699 16983
rect 6641 16943 6699 16949
rect 7374 16940 7380 16992
rect 7432 16940 7438 16992
rect 7742 16940 7748 16992
rect 7800 16980 7806 16992
rect 9968 16980 9996 17079
rect 10502 17076 10508 17088
rect 10560 17116 10566 17128
rect 10689 17119 10747 17125
rect 10689 17116 10701 17119
rect 10560 17088 10701 17116
rect 10560 17076 10566 17088
rect 10689 17085 10701 17088
rect 10735 17116 10747 17119
rect 11146 17116 11152 17128
rect 10735 17088 11152 17116
rect 10735 17085 10747 17088
rect 10689 17079 10747 17085
rect 11146 17076 11152 17088
rect 11204 17076 11210 17128
rect 11698 17076 11704 17128
rect 11756 17076 11762 17128
rect 14369 17119 14427 17125
rect 14369 17085 14381 17119
rect 14415 17085 14427 17119
rect 14369 17079 14427 17085
rect 14384 17048 14412 17079
rect 28350 17076 28356 17128
rect 28408 17076 28414 17128
rect 13372 17020 14412 17048
rect 7800 16952 9996 16980
rect 11333 16983 11391 16989
rect 7800 16940 7806 16952
rect 11333 16949 11345 16983
rect 11379 16980 11391 16983
rect 13372 16980 13400 17020
rect 11379 16952 13400 16980
rect 11379 16949 11391 16952
rect 11333 16943 11391 16949
rect 13814 16940 13820 16992
rect 13872 16940 13878 16992
rect 1104 16890 28888 16912
rect 1104 16838 4423 16890
rect 4475 16838 4487 16890
rect 4539 16838 4551 16890
rect 4603 16838 4615 16890
rect 4667 16838 4679 16890
rect 4731 16838 11369 16890
rect 11421 16838 11433 16890
rect 11485 16838 11497 16890
rect 11549 16838 11561 16890
rect 11613 16838 11625 16890
rect 11677 16838 18315 16890
rect 18367 16838 18379 16890
rect 18431 16838 18443 16890
rect 18495 16838 18507 16890
rect 18559 16838 18571 16890
rect 18623 16838 25261 16890
rect 25313 16838 25325 16890
rect 25377 16838 25389 16890
rect 25441 16838 25453 16890
rect 25505 16838 25517 16890
rect 25569 16838 28888 16890
rect 1104 16816 28888 16838
rect 8757 16779 8815 16785
rect 8757 16745 8769 16779
rect 8803 16776 8815 16779
rect 8803 16748 10916 16776
rect 8803 16745 8815 16748
rect 8757 16739 8815 16745
rect 10888 16708 10916 16748
rect 10962 16736 10968 16788
rect 11020 16776 11026 16788
rect 11241 16779 11299 16785
rect 11241 16776 11253 16779
rect 11020 16748 11253 16776
rect 11020 16736 11026 16748
rect 11241 16745 11253 16748
rect 11287 16776 11299 16779
rect 13630 16776 13636 16788
rect 11287 16748 13636 16776
rect 11287 16745 11299 16748
rect 11241 16739 11299 16745
rect 13630 16736 13636 16748
rect 13688 16736 13694 16788
rect 13814 16736 13820 16788
rect 13872 16736 13878 16788
rect 11054 16708 11060 16720
rect 10888 16680 11060 16708
rect 11054 16668 11060 16680
rect 11112 16668 11118 16720
rect 6365 16643 6423 16649
rect 6365 16609 6377 16643
rect 6411 16640 6423 16643
rect 6454 16640 6460 16652
rect 6411 16612 6460 16640
rect 6411 16609 6423 16612
rect 6365 16603 6423 16609
rect 6454 16600 6460 16612
rect 6512 16600 6518 16652
rect 8113 16643 8171 16649
rect 8113 16609 8125 16643
rect 8159 16640 8171 16643
rect 8294 16640 8300 16652
rect 8159 16612 8300 16640
rect 8159 16609 8171 16612
rect 8113 16603 8171 16609
rect 8294 16600 8300 16612
rect 8352 16600 8358 16652
rect 8386 16600 8392 16652
rect 8444 16600 8450 16652
rect 9217 16643 9275 16649
rect 9217 16609 9229 16643
rect 9263 16640 9275 16643
rect 9306 16640 9312 16652
rect 9263 16612 9312 16640
rect 9263 16609 9275 16612
rect 9217 16603 9275 16609
rect 9306 16600 9312 16612
rect 9364 16600 9370 16652
rect 10778 16600 10784 16652
rect 10836 16640 10842 16652
rect 11977 16643 12035 16649
rect 10836 16612 11008 16640
rect 10836 16600 10842 16612
rect 934 16532 940 16584
rect 992 16572 998 16584
rect 1397 16575 1455 16581
rect 1397 16572 1409 16575
rect 992 16544 1409 16572
rect 992 16532 998 16544
rect 1397 16541 1409 16544
rect 1443 16541 1455 16575
rect 1397 16535 1455 16541
rect 1857 16575 1915 16581
rect 1857 16541 1869 16575
rect 1903 16541 1915 16575
rect 1857 16535 1915 16541
rect 1026 16464 1032 16516
rect 1084 16504 1090 16516
rect 1872 16504 1900 16535
rect 5718 16532 5724 16584
rect 5776 16572 5782 16584
rect 6089 16575 6147 16581
rect 6089 16572 6101 16575
rect 5776 16544 6101 16572
rect 5776 16532 5782 16544
rect 6089 16541 6101 16544
rect 6135 16541 6147 16575
rect 6089 16535 6147 16541
rect 1084 16476 1900 16504
rect 1084 16464 1090 16476
rect 658 16396 664 16448
rect 716 16436 722 16448
rect 1581 16439 1639 16445
rect 1581 16436 1593 16439
rect 716 16408 1593 16436
rect 716 16396 722 16408
rect 1581 16405 1593 16408
rect 1627 16405 1639 16439
rect 1581 16399 1639 16405
rect 1670 16396 1676 16448
rect 1728 16396 1734 16448
rect 6104 16436 6132 16535
rect 8570 16532 8576 16584
rect 8628 16532 8634 16584
rect 10980 16581 11008 16612
rect 11977 16609 11989 16643
rect 12023 16640 12035 16643
rect 13832 16640 13860 16736
rect 12023 16612 13860 16640
rect 12023 16609 12035 16612
rect 11977 16603 12035 16609
rect 8941 16575 8999 16581
rect 8941 16541 8953 16575
rect 8987 16541 8999 16575
rect 8941 16535 8999 16541
rect 10965 16575 11023 16581
rect 10965 16541 10977 16575
rect 11011 16541 11023 16575
rect 11425 16575 11483 16581
rect 11425 16572 11437 16575
rect 10965 16535 11023 16541
rect 11348 16544 11437 16572
rect 6638 16464 6644 16516
rect 6696 16504 6702 16516
rect 8956 16504 8984 16535
rect 6696 16476 6854 16504
rect 8312 16476 8984 16504
rect 6696 16464 6702 16476
rect 8312 16448 8340 16476
rect 9858 16464 9864 16516
rect 9916 16464 9922 16516
rect 11348 16448 11376 16544
rect 11425 16541 11437 16544
rect 11471 16541 11483 16575
rect 11425 16535 11483 16541
rect 11698 16532 11704 16584
rect 11756 16532 11762 16584
rect 13630 16532 13636 16584
rect 13688 16572 13694 16584
rect 13725 16575 13783 16581
rect 13725 16572 13737 16575
rect 13688 16544 13737 16572
rect 13688 16532 13694 16544
rect 13725 16541 13737 16544
rect 13771 16572 13783 16575
rect 14642 16572 14648 16584
rect 13771 16544 14648 16572
rect 13771 16541 13783 16544
rect 13725 16535 13783 16541
rect 14642 16532 14648 16544
rect 14700 16532 14706 16584
rect 23474 16532 23480 16584
rect 23532 16572 23538 16584
rect 27157 16575 27215 16581
rect 27157 16572 27169 16575
rect 23532 16544 27169 16572
rect 23532 16532 23538 16544
rect 27157 16541 27169 16544
rect 27203 16541 27215 16575
rect 27157 16535 27215 16541
rect 13262 16504 13268 16516
rect 13202 16476 13268 16504
rect 13262 16464 13268 16476
rect 13320 16464 13326 16516
rect 28350 16464 28356 16516
rect 28408 16464 28414 16516
rect 8294 16436 8300 16448
rect 6104 16408 8300 16436
rect 8294 16396 8300 16408
rect 8352 16396 8358 16448
rect 11330 16396 11336 16448
rect 11388 16396 11394 16448
rect 11514 16396 11520 16448
rect 11572 16396 11578 16448
rect 1104 16346 29048 16368
rect 1104 16294 7896 16346
rect 7948 16294 7960 16346
rect 8012 16294 8024 16346
rect 8076 16294 8088 16346
rect 8140 16294 8152 16346
rect 8204 16294 14842 16346
rect 14894 16294 14906 16346
rect 14958 16294 14970 16346
rect 15022 16294 15034 16346
rect 15086 16294 15098 16346
rect 15150 16294 21788 16346
rect 21840 16294 21852 16346
rect 21904 16294 21916 16346
rect 21968 16294 21980 16346
rect 22032 16294 22044 16346
rect 22096 16294 28734 16346
rect 28786 16294 28798 16346
rect 28850 16294 28862 16346
rect 28914 16294 28926 16346
rect 28978 16294 28990 16346
rect 29042 16294 29048 16346
rect 1104 16272 29048 16294
rect 382 16192 388 16244
rect 440 16232 446 16244
rect 1670 16232 1676 16244
rect 440 16204 1676 16232
rect 440 16192 446 16204
rect 1670 16192 1676 16204
rect 1728 16192 1734 16244
rect 6638 16192 6644 16244
rect 6696 16192 6702 16244
rect 6825 16235 6883 16241
rect 6825 16201 6837 16235
rect 6871 16232 6883 16235
rect 7190 16232 7196 16244
rect 6871 16204 7196 16232
rect 6871 16201 6883 16204
rect 6825 16195 6883 16201
rect 7190 16192 7196 16204
rect 7248 16192 7254 16244
rect 7285 16235 7343 16241
rect 7285 16201 7297 16235
rect 7331 16232 7343 16235
rect 7374 16232 7380 16244
rect 7331 16204 7380 16232
rect 7331 16201 7343 16204
rect 7285 16195 7343 16201
rect 7374 16192 7380 16204
rect 7432 16192 7438 16244
rect 8386 16192 8392 16244
rect 8444 16192 8450 16244
rect 11514 16192 11520 16244
rect 11572 16232 11578 16244
rect 11572 16204 11928 16232
rect 11572 16192 11578 16204
rect 8404 16164 8432 16192
rect 11241 16167 11299 16173
rect 11241 16164 11253 16167
rect 7208 16136 8432 16164
rect 9798 16136 11253 16164
rect 934 16056 940 16108
rect 992 16096 998 16108
rect 7208 16105 7236 16136
rect 11241 16133 11253 16136
rect 11287 16133 11299 16167
rect 11698 16164 11704 16176
rect 11241 16127 11299 16133
rect 11532 16136 11704 16164
rect 1397 16099 1455 16105
rect 1397 16096 1409 16099
rect 992 16068 1409 16096
rect 992 16056 998 16068
rect 1397 16065 1409 16068
rect 1443 16065 1455 16099
rect 1397 16059 1455 16065
rect 1673 16099 1731 16105
rect 1673 16065 1685 16099
rect 1719 16065 1731 16099
rect 1673 16059 1731 16065
rect 6549 16099 6607 16105
rect 6549 16065 6561 16099
rect 6595 16096 6607 16099
rect 7193 16099 7251 16105
rect 6595 16068 6914 16096
rect 6595 16065 6607 16068
rect 6549 16059 6607 16065
rect 1026 15988 1032 16040
rect 1084 16028 1090 16040
rect 1688 16028 1716 16059
rect 1084 16000 1716 16028
rect 1084 15988 1090 16000
rect 6886 15960 6914 16068
rect 7193 16065 7205 16099
rect 7239 16065 7251 16099
rect 8021 16099 8079 16105
rect 8021 16096 8033 16099
rect 7193 16059 7251 16065
rect 7300 16068 8033 16096
rect 7006 15988 7012 16040
rect 7064 16028 7070 16040
rect 7300 16028 7328 16068
rect 8021 16065 8033 16068
rect 8067 16065 8079 16099
rect 8021 16059 8079 16065
rect 8294 16056 8300 16108
rect 8352 16056 8358 16108
rect 11330 16056 11336 16108
rect 11388 16056 11394 16108
rect 11532 16105 11560 16136
rect 11698 16124 11704 16136
rect 11756 16124 11762 16176
rect 11900 16164 11928 16204
rect 13262 16192 13268 16244
rect 13320 16232 13326 16244
rect 13725 16235 13783 16241
rect 13725 16232 13737 16235
rect 13320 16204 13737 16232
rect 13320 16192 13326 16204
rect 13725 16201 13737 16204
rect 13771 16201 13783 16235
rect 13725 16195 13783 16201
rect 11900 16136 12282 16164
rect 13078 16124 13084 16176
rect 13136 16164 13142 16176
rect 13541 16167 13599 16173
rect 13541 16164 13553 16167
rect 13136 16136 13553 16164
rect 13136 16124 13142 16136
rect 13541 16133 13553 16136
rect 13587 16164 13599 16167
rect 15194 16164 15200 16176
rect 13587 16136 15200 16164
rect 13587 16133 13599 16136
rect 13541 16127 13599 16133
rect 15194 16124 15200 16136
rect 15252 16164 15258 16176
rect 15746 16164 15752 16176
rect 15252 16136 15752 16164
rect 15252 16124 15258 16136
rect 15746 16124 15752 16136
rect 15804 16124 15810 16176
rect 11517 16099 11575 16105
rect 11517 16065 11529 16099
rect 11563 16065 11575 16099
rect 13817 16099 13875 16105
rect 13817 16096 13829 16099
rect 11517 16059 11575 16065
rect 13280 16068 13829 16096
rect 7064 16000 7328 16028
rect 7064 15988 7070 16000
rect 7374 15988 7380 16040
rect 7432 15988 7438 16040
rect 7466 15988 7472 16040
rect 7524 16028 7530 16040
rect 7837 16031 7895 16037
rect 7837 16028 7849 16031
rect 7524 16000 7849 16028
rect 7524 15988 7530 16000
rect 7837 15997 7849 16000
rect 7883 15997 7895 16031
rect 7837 15991 7895 15997
rect 8573 16031 8631 16037
rect 8573 15997 8585 16031
rect 8619 16028 8631 16031
rect 8619 16000 9628 16028
rect 8619 15997 8631 16000
rect 8573 15991 8631 15997
rect 7650 15960 7656 15972
rect 6886 15932 7656 15960
rect 7650 15920 7656 15932
rect 7708 15920 7714 15972
rect 7742 15920 7748 15972
rect 7800 15920 7806 15972
rect 9600 15960 9628 16000
rect 10318 15988 10324 16040
rect 10376 15988 10382 16040
rect 10962 15988 10968 16040
rect 11020 15988 11026 16040
rect 10413 15963 10471 15969
rect 10413 15960 10425 15963
rect 9600 15932 10425 15960
rect 10413 15929 10425 15932
rect 10459 15929 10471 15963
rect 10413 15923 10471 15929
rect 1581 15895 1639 15901
rect 1581 15861 1593 15895
rect 1627 15892 1639 15895
rect 1670 15892 1676 15904
rect 1627 15864 1676 15892
rect 1627 15861 1639 15864
rect 1581 15855 1639 15861
rect 1670 15852 1676 15864
rect 1728 15852 1734 15904
rect 1857 15895 1915 15901
rect 1857 15861 1869 15895
rect 1903 15892 1915 15895
rect 3234 15892 3240 15904
rect 1903 15864 3240 15892
rect 1903 15861 1915 15864
rect 1857 15855 1915 15861
rect 3234 15852 3240 15864
rect 3292 15852 3298 15904
rect 7374 15852 7380 15904
rect 7432 15892 7438 15904
rect 7760 15892 7788 15920
rect 7432 15864 7788 15892
rect 7432 15852 7438 15864
rect 8202 15852 8208 15904
rect 8260 15852 8266 15904
rect 9674 15852 9680 15904
rect 9732 15892 9738 15904
rect 11348 15892 11376 16056
rect 11790 15988 11796 16040
rect 11848 15988 11854 16040
rect 13280 15904 13308 16068
rect 13817 16065 13829 16068
rect 13863 16065 13875 16099
rect 13817 16059 13875 16065
rect 13262 15892 13268 15904
rect 9732 15864 13268 15892
rect 9732 15852 9738 15864
rect 13262 15852 13268 15864
rect 13320 15852 13326 15904
rect 1104 15802 28888 15824
rect 1104 15750 4423 15802
rect 4475 15750 4487 15802
rect 4539 15750 4551 15802
rect 4603 15750 4615 15802
rect 4667 15750 4679 15802
rect 4731 15750 11369 15802
rect 11421 15750 11433 15802
rect 11485 15750 11497 15802
rect 11549 15750 11561 15802
rect 11613 15750 11625 15802
rect 11677 15750 18315 15802
rect 18367 15750 18379 15802
rect 18431 15750 18443 15802
rect 18495 15750 18507 15802
rect 18559 15750 18571 15802
rect 18623 15750 25261 15802
rect 25313 15750 25325 15802
rect 25377 15750 25389 15802
rect 25441 15750 25453 15802
rect 25505 15750 25517 15802
rect 25569 15750 28888 15802
rect 1104 15728 28888 15750
rect 8202 15648 8208 15700
rect 8260 15648 8266 15700
rect 9858 15648 9864 15700
rect 9916 15648 9922 15700
rect 10962 15648 10968 15700
rect 11020 15648 11026 15700
rect 11146 15648 11152 15700
rect 11204 15648 11210 15700
rect 11790 15648 11796 15700
rect 11848 15688 11854 15700
rect 11977 15691 12035 15697
rect 11977 15688 11989 15691
rect 11848 15660 11989 15688
rect 11848 15648 11854 15660
rect 11977 15657 11989 15660
rect 12023 15657 12035 15691
rect 11977 15651 12035 15657
rect 13078 15648 13084 15700
rect 13136 15648 13142 15700
rect 13170 15648 13176 15700
rect 13228 15688 13234 15700
rect 13541 15691 13599 15697
rect 13541 15688 13553 15691
rect 13228 15660 13553 15688
rect 13228 15648 13234 15660
rect 13541 15657 13553 15660
rect 13587 15657 13599 15691
rect 13541 15651 13599 15657
rect 14274 15648 14280 15700
rect 14332 15648 14338 15700
rect 934 15580 940 15632
rect 992 15620 998 15632
rect 1673 15623 1731 15629
rect 1673 15620 1685 15623
rect 992 15592 1685 15620
rect 992 15580 998 15592
rect 1673 15589 1685 15592
rect 1719 15589 1731 15623
rect 8220 15620 8248 15648
rect 9677 15623 9735 15629
rect 8220 15592 9260 15620
rect 1673 15583 1731 15589
rect 7745 15555 7803 15561
rect 7745 15521 7757 15555
rect 7791 15552 7803 15555
rect 8386 15552 8392 15564
rect 7791 15524 8392 15552
rect 7791 15521 7803 15524
rect 7745 15515 7803 15521
rect 8386 15512 8392 15524
rect 8444 15512 8450 15564
rect 9232 15561 9260 15592
rect 9677 15589 9689 15623
rect 9723 15620 9735 15623
rect 10980 15620 11008 15648
rect 9723 15592 11008 15620
rect 9723 15589 9735 15592
rect 9677 15583 9735 15589
rect 9033 15555 9091 15561
rect 9033 15552 9045 15555
rect 8772 15524 9045 15552
rect 934 15444 940 15496
rect 992 15484 998 15496
rect 1397 15487 1455 15493
rect 1397 15484 1409 15487
rect 992 15456 1409 15484
rect 992 15444 998 15456
rect 1397 15453 1409 15456
rect 1443 15453 1455 15487
rect 1397 15447 1455 15453
rect 1578 15444 1584 15496
rect 1636 15444 1642 15496
rect 1854 15444 1860 15496
rect 1912 15444 1918 15496
rect 1596 15416 1624 15444
rect 7742 15416 7748 15428
rect 1596 15388 7748 15416
rect 7742 15376 7748 15388
rect 7800 15376 7806 15428
rect 8772 15360 8800 15524
rect 9033 15521 9045 15524
rect 9079 15521 9091 15555
rect 9033 15515 9091 15521
rect 9217 15555 9275 15561
rect 9217 15521 9229 15555
rect 9263 15521 9275 15555
rect 9217 15515 9275 15521
rect 11054 15512 11060 15564
rect 11112 15512 11118 15564
rect 11164 15552 11192 15648
rect 11885 15623 11943 15629
rect 11885 15589 11897 15623
rect 11931 15620 11943 15623
rect 11931 15592 12434 15620
rect 11931 15589 11943 15592
rect 11885 15583 11943 15589
rect 11241 15555 11299 15561
rect 11241 15552 11253 15555
rect 11164 15524 11253 15552
rect 11241 15521 11253 15524
rect 11287 15552 11299 15555
rect 12250 15552 12256 15564
rect 11287 15524 12256 15552
rect 11287 15521 11299 15524
rect 11241 15515 11299 15521
rect 12250 15512 12256 15524
rect 12308 15512 12314 15564
rect 12406 15552 12434 15592
rect 12529 15555 12587 15561
rect 12529 15552 12541 15555
rect 12406 15524 12541 15552
rect 12529 15521 12541 15524
rect 12575 15521 12587 15555
rect 12529 15515 12587 15521
rect 9769 15487 9827 15493
rect 9769 15484 9781 15487
rect 9692 15456 9781 15484
rect 9692 15428 9720 15456
rect 9769 15453 9781 15456
rect 9815 15453 9827 15487
rect 11072 15484 11100 15512
rect 11425 15487 11483 15493
rect 11425 15484 11437 15487
rect 11072 15456 11437 15484
rect 9769 15447 9827 15453
rect 11425 15453 11437 15456
rect 11471 15453 11483 15487
rect 13096 15484 13124 15648
rect 13262 15580 13268 15632
rect 13320 15580 13326 15632
rect 13280 15552 13308 15580
rect 13280 15524 13676 15552
rect 11425 15447 11483 15453
rect 11532 15456 13124 15484
rect 9674 15376 9680 15428
rect 9732 15376 9738 15428
rect 11532 15425 11560 15456
rect 13262 15444 13268 15496
rect 13320 15444 13326 15496
rect 13648 15493 13676 15524
rect 13633 15487 13691 15493
rect 13633 15453 13645 15487
rect 13679 15453 13691 15487
rect 13633 15447 13691 15453
rect 27157 15487 27215 15493
rect 27157 15453 27169 15487
rect 27203 15453 27215 15487
rect 27157 15447 27215 15453
rect 11057 15419 11115 15425
rect 11057 15385 11069 15419
rect 11103 15416 11115 15419
rect 11517 15419 11575 15425
rect 11517 15416 11529 15419
rect 11103 15388 11529 15416
rect 11103 15385 11115 15388
rect 11057 15379 11115 15385
rect 11517 15385 11529 15388
rect 11563 15385 11575 15419
rect 16206 15416 16212 15428
rect 11517 15379 11575 15385
rect 11624 15388 16212 15416
rect 474 15308 480 15360
rect 532 15348 538 15360
rect 1581 15351 1639 15357
rect 1581 15348 1593 15351
rect 532 15320 1593 15348
rect 532 15308 538 15320
rect 1581 15317 1593 15320
rect 1627 15317 1639 15351
rect 1581 15311 1639 15317
rect 8754 15308 8760 15360
rect 8812 15308 8818 15360
rect 9309 15351 9367 15357
rect 9309 15317 9321 15351
rect 9355 15348 9367 15351
rect 10318 15348 10324 15360
rect 9355 15320 10324 15348
rect 9355 15317 9367 15320
rect 9309 15311 9367 15317
rect 10318 15308 10324 15320
rect 10376 15348 10382 15360
rect 11624 15348 11652 15388
rect 16206 15376 16212 15388
rect 16264 15376 16270 15428
rect 10376 15320 11652 15348
rect 10376 15308 10382 15320
rect 12342 15308 12348 15360
rect 12400 15348 12406 15360
rect 12713 15351 12771 15357
rect 12713 15348 12725 15351
rect 12400 15320 12725 15348
rect 12400 15308 12406 15320
rect 12713 15317 12725 15320
rect 12759 15317 12771 15351
rect 12713 15311 12771 15317
rect 26970 15308 26976 15360
rect 27028 15348 27034 15360
rect 27172 15348 27200 15447
rect 28350 15376 28356 15428
rect 28408 15376 28414 15428
rect 27028 15320 27200 15348
rect 27028 15308 27034 15320
rect 1104 15258 29048 15280
rect 1104 15206 7896 15258
rect 7948 15206 7960 15258
rect 8012 15206 8024 15258
rect 8076 15206 8088 15258
rect 8140 15206 8152 15258
rect 8204 15206 14842 15258
rect 14894 15206 14906 15258
rect 14958 15206 14970 15258
rect 15022 15206 15034 15258
rect 15086 15206 15098 15258
rect 15150 15206 21788 15258
rect 21840 15206 21852 15258
rect 21904 15206 21916 15258
rect 21968 15206 21980 15258
rect 22032 15206 22044 15258
rect 22096 15206 28734 15258
rect 28786 15206 28798 15258
rect 28850 15206 28862 15258
rect 28914 15206 28926 15258
rect 28978 15206 28990 15258
rect 29042 15206 29048 15258
rect 1104 15184 29048 15206
rect 1581 15147 1639 15153
rect 1581 15113 1593 15147
rect 1627 15144 1639 15147
rect 12897 15147 12955 15153
rect 1627 15116 12848 15144
rect 1627 15113 1639 15116
rect 1581 15107 1639 15113
rect 1762 15036 1768 15088
rect 1820 15076 1826 15088
rect 1820 15048 9812 15076
rect 1820 15036 1826 15048
rect 934 14968 940 15020
rect 992 15008 998 15020
rect 1397 15011 1455 15017
rect 1397 15008 1409 15011
rect 992 14980 1409 15008
rect 992 14968 998 14980
rect 1397 14977 1409 14980
rect 1443 14977 1455 15011
rect 1397 14971 1455 14977
rect 5626 14968 5632 15020
rect 5684 15008 5690 15020
rect 5684 14980 7052 15008
rect 5684 14968 5690 14980
rect 6914 14900 6920 14952
rect 6972 14900 6978 14952
rect 7024 14940 7052 14980
rect 7282 14968 7288 15020
rect 7340 14968 7346 15020
rect 7650 14968 7656 15020
rect 7708 15008 7714 15020
rect 7745 15011 7803 15017
rect 7745 15008 7757 15011
rect 7708 14980 7757 15008
rect 7708 14968 7714 14980
rect 7745 14977 7757 14980
rect 7791 15008 7803 15011
rect 9674 15008 9680 15020
rect 7791 14980 9680 15008
rect 7791 14977 7803 14980
rect 7745 14971 7803 14977
rect 9674 14968 9680 14980
rect 9732 14968 9738 15020
rect 7469 14943 7527 14949
rect 7469 14940 7481 14943
rect 7024 14912 7481 14940
rect 7469 14909 7481 14912
rect 7515 14909 7527 14943
rect 7469 14903 7527 14909
rect 9784 14884 9812 15048
rect 11882 15036 11888 15088
rect 11940 15076 11946 15088
rect 12437 15079 12495 15085
rect 12437 15076 12449 15079
rect 11940 15048 12449 15076
rect 11940 15036 11946 15048
rect 12437 15045 12449 15048
rect 12483 15045 12495 15079
rect 12820 15076 12848 15116
rect 12897 15113 12909 15147
rect 12943 15144 12955 15147
rect 13262 15144 13268 15156
rect 12943 15116 13268 15144
rect 12943 15113 12955 15116
rect 12897 15107 12955 15113
rect 13262 15104 13268 15116
rect 13320 15104 13326 15156
rect 13357 15147 13415 15153
rect 13357 15113 13369 15147
rect 13403 15144 13415 15147
rect 14274 15144 14280 15156
rect 13403 15116 14280 15144
rect 13403 15113 13415 15116
rect 13357 15107 13415 15113
rect 14274 15104 14280 15116
rect 14332 15104 14338 15156
rect 14645 15147 14703 15153
rect 14645 15113 14657 15147
rect 14691 15144 14703 15147
rect 14734 15144 14740 15156
rect 14691 15116 14740 15144
rect 14691 15113 14703 15116
rect 14645 15107 14703 15113
rect 14734 15104 14740 15116
rect 14792 15104 14798 15156
rect 12820 15048 15792 15076
rect 12437 15039 12495 15045
rect 12069 15011 12127 15017
rect 12069 14977 12081 15011
rect 12115 15008 12127 15011
rect 12529 15011 12587 15017
rect 12529 15008 12541 15011
rect 12115 14980 12541 15008
rect 12115 14977 12127 14980
rect 12069 14971 12127 14977
rect 12529 14977 12541 14980
rect 12575 15008 12587 15011
rect 12575 14980 13584 15008
rect 12575 14977 12587 14980
rect 12529 14971 12587 14977
rect 12250 14940 12256 14952
rect 12211 14912 12256 14940
rect 12250 14900 12256 14912
rect 12308 14940 12314 14952
rect 13081 14943 13139 14949
rect 13081 14940 13093 14943
rect 12308 14912 13093 14940
rect 12308 14900 12314 14912
rect 13081 14909 13093 14912
rect 13127 14909 13139 14943
rect 13265 14943 13323 14949
rect 13265 14940 13277 14943
rect 13081 14903 13139 14909
rect 13188 14912 13277 14940
rect 1578 14832 1584 14884
rect 1636 14872 1642 14884
rect 1636 14844 7788 14872
rect 1636 14832 1642 14844
rect 6270 14764 6276 14816
rect 6328 14804 6334 14816
rect 6365 14807 6423 14813
rect 6365 14804 6377 14807
rect 6328 14776 6377 14804
rect 6328 14764 6334 14776
rect 6365 14773 6377 14776
rect 6411 14773 6423 14807
rect 6365 14767 6423 14773
rect 7098 14764 7104 14816
rect 7156 14764 7162 14816
rect 7650 14764 7656 14816
rect 7708 14764 7714 14816
rect 7760 14804 7788 14844
rect 9766 14832 9772 14884
rect 9824 14832 9830 14884
rect 10962 14832 10968 14884
rect 11020 14872 11026 14884
rect 13188 14872 13216 14912
rect 13265 14909 13277 14912
rect 13311 14909 13323 14943
rect 13265 14903 13323 14909
rect 13556 14884 13584 14980
rect 13722 14968 13728 15020
rect 13780 14968 13786 15020
rect 14277 15011 14335 15017
rect 14277 14977 14289 15011
rect 14323 15008 14335 15011
rect 14734 15008 14740 15020
rect 14323 14980 14740 15008
rect 14323 14977 14335 14980
rect 14277 14971 14335 14977
rect 14734 14968 14740 14980
rect 14792 14968 14798 15020
rect 13740 14940 13768 14968
rect 15286 14940 15292 14952
rect 13740 14912 15292 14940
rect 15286 14900 15292 14912
rect 15344 14900 15350 14952
rect 11020 14844 13216 14872
rect 11020 14832 11026 14844
rect 13538 14832 13544 14884
rect 13596 14832 13602 14884
rect 13648 14844 15516 14872
rect 13648 14804 13676 14844
rect 15488 14816 15516 14844
rect 15764 14816 15792 15048
rect 27157 15011 27215 15017
rect 27157 15008 27169 15011
rect 26712 14980 27169 15008
rect 7760 14776 13676 14804
rect 13722 14764 13728 14816
rect 13780 14764 13786 14816
rect 14182 14764 14188 14816
rect 14240 14764 14246 14816
rect 15470 14764 15476 14816
rect 15528 14764 15534 14816
rect 15746 14764 15752 14816
rect 15804 14764 15810 14816
rect 15930 14764 15936 14816
rect 15988 14804 15994 14816
rect 26712 14813 26740 14980
rect 27157 14977 27169 14980
rect 27203 14977 27215 15011
rect 27157 14971 27215 14977
rect 28350 14900 28356 14952
rect 28408 14900 28414 14952
rect 26697 14807 26755 14813
rect 26697 14804 26709 14807
rect 15988 14776 26709 14804
rect 15988 14764 15994 14776
rect 26697 14773 26709 14776
rect 26743 14773 26755 14807
rect 26697 14767 26755 14773
rect 1104 14714 28888 14736
rect 1104 14662 4423 14714
rect 4475 14662 4487 14714
rect 4539 14662 4551 14714
rect 4603 14662 4615 14714
rect 4667 14662 4679 14714
rect 4731 14662 11369 14714
rect 11421 14662 11433 14714
rect 11485 14662 11497 14714
rect 11549 14662 11561 14714
rect 11613 14662 11625 14714
rect 11677 14662 18315 14714
rect 18367 14662 18379 14714
rect 18431 14662 18443 14714
rect 18495 14662 18507 14714
rect 18559 14662 18571 14714
rect 18623 14662 25261 14714
rect 25313 14662 25325 14714
rect 25377 14662 25389 14714
rect 25441 14662 25453 14714
rect 25505 14662 25517 14714
rect 25569 14662 28888 14714
rect 1104 14640 28888 14662
rect 1581 14603 1639 14609
rect 1581 14569 1593 14603
rect 1627 14600 1639 14603
rect 1627 14572 7604 14600
rect 1627 14569 1639 14572
rect 1581 14563 1639 14569
rect 7576 14532 7604 14572
rect 8294 14560 8300 14612
rect 8352 14600 8358 14612
rect 11425 14603 11483 14609
rect 8352 14572 11284 14600
rect 8352 14560 8358 14572
rect 7576 14504 11192 14532
rect 6181 14467 6239 14473
rect 6181 14433 6193 14467
rect 6227 14464 6239 14467
rect 6270 14464 6276 14476
rect 6227 14436 6276 14464
rect 6227 14433 6239 14436
rect 6181 14427 6239 14433
rect 6270 14424 6276 14436
rect 6328 14424 6334 14476
rect 9766 14424 9772 14476
rect 9824 14464 9830 14476
rect 11057 14467 11115 14473
rect 11057 14464 11069 14467
rect 9824 14436 11069 14464
rect 9824 14424 9830 14436
rect 11057 14433 11069 14436
rect 11103 14433 11115 14467
rect 11057 14427 11115 14433
rect 934 14356 940 14408
rect 992 14396 998 14408
rect 1397 14399 1455 14405
rect 1397 14396 1409 14399
rect 992 14368 1409 14396
rect 992 14356 998 14368
rect 1397 14365 1409 14368
rect 1443 14365 1455 14399
rect 1397 14359 1455 14365
rect 1673 14399 1731 14405
rect 1673 14365 1685 14399
rect 1719 14365 1731 14399
rect 1673 14359 1731 14365
rect 1026 14288 1032 14340
rect 1084 14328 1090 14340
rect 1688 14328 1716 14359
rect 5718 14356 5724 14408
rect 5776 14396 5782 14408
rect 5905 14399 5963 14405
rect 5905 14396 5917 14399
rect 5776 14368 5917 14396
rect 5776 14356 5782 14368
rect 5905 14365 5917 14368
rect 5951 14365 5963 14399
rect 7650 14396 7656 14408
rect 7314 14368 7656 14396
rect 5905 14359 5963 14365
rect 7650 14356 7656 14368
rect 7708 14356 7714 14408
rect 9585 14399 9643 14405
rect 9585 14365 9597 14399
rect 9631 14396 9643 14399
rect 9674 14396 9680 14408
rect 9631 14368 9680 14396
rect 9631 14365 9643 14368
rect 9585 14359 9643 14365
rect 9674 14356 9680 14368
rect 9732 14396 9738 14408
rect 10318 14396 10324 14408
rect 9732 14368 10324 14396
rect 9732 14356 9738 14368
rect 10318 14356 10324 14368
rect 10376 14356 10382 14408
rect 10410 14356 10416 14408
rect 10468 14356 10474 14408
rect 10597 14399 10655 14405
rect 10597 14365 10609 14399
rect 10643 14365 10655 14399
rect 10597 14359 10655 14365
rect 1084 14300 1716 14328
rect 1084 14288 1090 14300
rect 7466 14288 7472 14340
rect 7524 14328 7530 14340
rect 7929 14331 7987 14337
rect 7929 14328 7941 14331
rect 7524 14300 7941 14328
rect 7524 14288 7530 14300
rect 7929 14297 7941 14300
rect 7975 14297 7987 14331
rect 10612 14328 10640 14359
rect 10778 14356 10784 14408
rect 10836 14356 10842 14408
rect 10962 14356 10968 14408
rect 11020 14356 11026 14408
rect 7929 14291 7987 14297
rect 8036 14300 10640 14328
rect 11164 14328 11192 14504
rect 11256 14464 11284 14572
rect 11425 14569 11437 14603
rect 11471 14600 11483 14603
rect 11882 14600 11888 14612
rect 11471 14572 11888 14600
rect 11471 14569 11483 14572
rect 11425 14563 11483 14569
rect 11882 14560 11888 14572
rect 11940 14560 11946 14612
rect 12148 14603 12206 14609
rect 12148 14569 12160 14603
rect 12194 14600 12206 14603
rect 12342 14600 12348 14612
rect 12194 14572 12348 14600
rect 12194 14569 12206 14572
rect 12148 14563 12206 14569
rect 12342 14560 12348 14572
rect 12400 14560 12406 14612
rect 13722 14560 13728 14612
rect 13780 14600 13786 14612
rect 13780 14572 14688 14600
rect 13780 14560 13786 14572
rect 14182 14492 14188 14544
rect 14240 14492 14246 14544
rect 14200 14464 14228 14492
rect 14660 14473 14688 14572
rect 11256 14436 13216 14464
rect 13188 14408 13216 14436
rect 13280 14436 14228 14464
rect 14645 14467 14703 14473
rect 11238 14356 11244 14408
rect 11296 14356 11302 14408
rect 11882 14356 11888 14408
rect 11940 14356 11946 14408
rect 13170 14356 13176 14408
rect 13228 14356 13234 14408
rect 13280 14382 13308 14436
rect 14645 14433 14657 14467
rect 14691 14433 14703 14467
rect 14645 14427 14703 14433
rect 14734 14424 14740 14476
rect 14792 14464 14798 14476
rect 15473 14467 15531 14473
rect 14792 14436 15056 14464
rect 14792 14424 14798 14436
rect 15028 14405 15056 14436
rect 15473 14433 15485 14467
rect 15519 14464 15531 14467
rect 15565 14467 15623 14473
rect 15565 14464 15577 14467
rect 15519 14436 15577 14464
rect 15519 14433 15531 14436
rect 15473 14427 15531 14433
rect 15565 14433 15577 14436
rect 15611 14464 15623 14467
rect 22738 14464 22744 14476
rect 15611 14436 22744 14464
rect 15611 14433 15623 14436
rect 15565 14427 15623 14433
rect 15013 14399 15071 14405
rect 15013 14365 15025 14399
rect 15059 14365 15071 14399
rect 15013 14359 15071 14365
rect 11164 14300 12388 14328
rect 1854 14220 1860 14272
rect 1912 14220 1918 14272
rect 1946 14220 1952 14272
rect 2004 14260 2010 14272
rect 8036 14260 8064 14300
rect 12360 14272 12388 14300
rect 13538 14288 13544 14340
rect 13596 14328 13602 14340
rect 13909 14331 13967 14337
rect 13909 14328 13921 14331
rect 13596 14300 13921 14328
rect 13596 14288 13602 14300
rect 13909 14297 13921 14300
rect 13955 14328 13967 14331
rect 15488 14328 15516 14427
rect 22738 14424 22744 14436
rect 22796 14424 22802 14476
rect 15746 14356 15752 14408
rect 15804 14356 15810 14408
rect 13955 14300 15516 14328
rect 13955 14297 13967 14300
rect 13909 14291 13967 14297
rect 2004 14232 8064 14260
rect 2004 14220 2010 14232
rect 9766 14220 9772 14272
rect 9824 14260 9830 14272
rect 9861 14263 9919 14269
rect 9861 14260 9873 14263
rect 9824 14232 9873 14260
rect 9824 14220 9830 14232
rect 9861 14229 9873 14232
rect 9907 14229 9919 14263
rect 9861 14223 9919 14229
rect 12342 14220 12348 14272
rect 12400 14220 12406 14272
rect 12434 14220 12440 14272
rect 12492 14260 12498 14272
rect 14093 14263 14151 14269
rect 14093 14260 14105 14263
rect 12492 14232 14105 14260
rect 12492 14220 12498 14232
rect 14093 14229 14105 14232
rect 14139 14229 14151 14263
rect 14093 14223 14151 14229
rect 14182 14220 14188 14272
rect 14240 14260 14246 14272
rect 14921 14263 14979 14269
rect 14921 14260 14933 14263
rect 14240 14232 14933 14260
rect 14240 14220 14246 14232
rect 14921 14229 14933 14232
rect 14967 14229 14979 14263
rect 14921 14223 14979 14229
rect 15933 14263 15991 14269
rect 15933 14229 15945 14263
rect 15979 14260 15991 14263
rect 16298 14260 16304 14272
rect 15979 14232 16304 14260
rect 15979 14229 15991 14232
rect 15933 14223 15991 14229
rect 16298 14220 16304 14232
rect 16356 14220 16362 14272
rect 1104 14170 29048 14192
rect 1104 14118 7896 14170
rect 7948 14118 7960 14170
rect 8012 14118 8024 14170
rect 8076 14118 8088 14170
rect 8140 14118 8152 14170
rect 8204 14118 14842 14170
rect 14894 14118 14906 14170
rect 14958 14118 14970 14170
rect 15022 14118 15034 14170
rect 15086 14118 15098 14170
rect 15150 14118 21788 14170
rect 21840 14118 21852 14170
rect 21904 14118 21916 14170
rect 21968 14118 21980 14170
rect 22032 14118 22044 14170
rect 22096 14118 28734 14170
rect 28786 14118 28798 14170
rect 28850 14118 28862 14170
rect 28914 14118 28926 14170
rect 28978 14118 28990 14170
rect 29042 14118 29048 14170
rect 1104 14096 29048 14118
rect 1578 14016 1584 14068
rect 1636 14016 1642 14068
rect 1854 14016 1860 14068
rect 1912 14016 1918 14068
rect 6549 14059 6607 14065
rect 6549 14025 6561 14059
rect 6595 14056 6607 14059
rect 6914 14056 6920 14068
rect 6595 14028 6920 14056
rect 6595 14025 6607 14028
rect 6549 14019 6607 14025
rect 6914 14016 6920 14028
rect 6972 14016 6978 14068
rect 7009 14059 7067 14065
rect 7009 14025 7021 14059
rect 7055 14056 7067 14059
rect 7098 14056 7104 14068
rect 7055 14028 7104 14056
rect 7055 14025 7067 14028
rect 7009 14019 7067 14025
rect 7098 14016 7104 14028
rect 7156 14016 7162 14068
rect 9033 14059 9091 14065
rect 9033 14025 9045 14059
rect 9079 14056 9091 14059
rect 9674 14056 9680 14068
rect 9079 14028 9680 14056
rect 9079 14025 9091 14028
rect 9033 14019 9091 14025
rect 9674 14016 9680 14028
rect 9732 14016 9738 14068
rect 9953 14059 10011 14065
rect 9953 14025 9965 14059
rect 9999 14056 10011 14059
rect 10410 14056 10416 14068
rect 9999 14028 10416 14056
rect 9999 14025 10011 14028
rect 9953 14019 10011 14025
rect 10410 14016 10416 14028
rect 10468 14016 10474 14068
rect 11149 14059 11207 14065
rect 11149 14025 11161 14059
rect 11195 14056 11207 14059
rect 12526 14056 12532 14068
rect 11195 14028 12532 14056
rect 11195 14025 11207 14028
rect 11149 14019 11207 14025
rect 12526 14016 12532 14028
rect 12584 14016 12590 14068
rect 13170 14016 13176 14068
rect 13228 14056 13234 14068
rect 26697 14059 26755 14065
rect 26697 14056 26709 14059
rect 13228 14028 26709 14056
rect 13228 14016 13234 14028
rect 26697 14025 26709 14028
rect 26743 14025 26755 14059
rect 26697 14019 26755 14025
rect 7466 13988 7472 14000
rect 6932 13960 7472 13988
rect 1394 13880 1400 13932
rect 1452 13880 1458 13932
rect 1670 13880 1676 13932
rect 1728 13880 1734 13932
rect 6932 13929 6960 13960
rect 7466 13948 7472 13960
rect 7524 13988 7530 14000
rect 7653 13991 7711 13997
rect 7653 13988 7665 13991
rect 7524 13960 7665 13988
rect 7524 13948 7530 13960
rect 7653 13957 7665 13960
rect 7699 13988 7711 13991
rect 10042 13988 10048 14000
rect 7699 13960 10048 13988
rect 7699 13957 7711 13960
rect 7653 13951 7711 13957
rect 10042 13948 10048 13960
rect 10100 13948 10106 14000
rect 10321 13991 10379 13997
rect 10321 13957 10333 13991
rect 10367 13988 10379 13991
rect 11054 13988 11060 14000
rect 10367 13960 11060 13988
rect 10367 13957 10379 13960
rect 10321 13951 10379 13957
rect 11054 13948 11060 13960
rect 11112 13988 11118 14000
rect 11701 13991 11759 13997
rect 11701 13988 11713 13991
rect 11112 13960 11713 13988
rect 11112 13948 11118 13960
rect 11701 13957 11713 13960
rect 11747 13957 11759 13991
rect 11701 13951 11759 13957
rect 12345 13991 12403 13997
rect 12345 13957 12357 13991
rect 12391 13988 12403 13991
rect 12434 13988 12440 14000
rect 12391 13960 12440 13988
rect 12391 13957 12403 13960
rect 12345 13951 12403 13957
rect 12434 13948 12440 13960
rect 12492 13948 12498 14000
rect 14182 13988 14188 14000
rect 13570 13960 14188 13988
rect 14182 13948 14188 13960
rect 14240 13948 14246 14000
rect 14734 13948 14740 14000
rect 14792 13948 14798 14000
rect 15565 13991 15623 13997
rect 15565 13957 15577 13991
rect 15611 13988 15623 13991
rect 17678 13988 17684 14000
rect 15611 13960 17684 13988
rect 15611 13957 15623 13960
rect 15565 13951 15623 13957
rect 17678 13948 17684 13960
rect 17736 13948 17742 14000
rect 6917 13923 6975 13929
rect 6917 13889 6929 13923
rect 6963 13889 6975 13923
rect 6917 13883 6975 13889
rect 8386 13880 8392 13932
rect 8444 13920 8450 13932
rect 9490 13920 9496 13932
rect 8444 13892 9496 13920
rect 8444 13880 8450 13892
rect 9490 13880 9496 13892
rect 9548 13880 9554 13932
rect 9582 13880 9588 13932
rect 9640 13920 9646 13932
rect 9677 13923 9735 13929
rect 9677 13920 9689 13923
rect 9640 13892 9689 13920
rect 9640 13880 9646 13892
rect 9677 13889 9689 13892
rect 9723 13889 9735 13923
rect 9677 13883 9735 13889
rect 7098 13812 7104 13864
rect 7156 13852 7162 13864
rect 7193 13855 7251 13861
rect 7193 13852 7205 13855
rect 7156 13824 7205 13852
rect 7156 13812 7162 13824
rect 7193 13821 7205 13824
rect 7239 13852 7251 13855
rect 7374 13852 7380 13864
rect 7239 13824 7380 13852
rect 7239 13821 7251 13824
rect 7193 13815 7251 13821
rect 7374 13812 7380 13824
rect 7432 13812 7438 13864
rect 9122 13812 9128 13864
rect 9180 13812 9186 13864
rect 9306 13812 9312 13864
rect 9364 13812 9370 13864
rect 2038 13744 2044 13796
rect 2096 13784 2102 13796
rect 6730 13784 6736 13796
rect 2096 13756 6736 13784
rect 2096 13744 2102 13756
rect 6730 13744 6736 13756
rect 6788 13744 6794 13796
rect 8573 13787 8631 13793
rect 8573 13753 8585 13787
rect 8619 13784 8631 13787
rect 8754 13784 8760 13796
rect 8619 13756 8760 13784
rect 8619 13753 8631 13756
rect 8573 13747 8631 13753
rect 8754 13744 8760 13756
rect 8812 13784 8818 13796
rect 9324 13784 9352 13812
rect 8812 13756 9352 13784
rect 9692 13784 9720 13883
rect 10134 13880 10140 13932
rect 10192 13920 10198 13932
rect 10781 13923 10839 13929
rect 10781 13920 10793 13923
rect 10192 13892 10793 13920
rect 10192 13880 10198 13892
rect 10781 13889 10793 13892
rect 10827 13889 10839 13923
rect 10781 13883 10839 13889
rect 10962 13880 10968 13932
rect 11020 13880 11026 13932
rect 15381 13923 15439 13929
rect 15381 13920 15393 13923
rect 13924 13892 15393 13920
rect 10410 13812 10416 13864
rect 10468 13812 10474 13864
rect 10597 13855 10655 13861
rect 10597 13821 10609 13855
rect 10643 13852 10655 13855
rect 10643 13824 11284 13852
rect 10643 13821 10655 13824
rect 10597 13815 10655 13821
rect 11256 13784 11284 13824
rect 11882 13812 11888 13864
rect 11940 13852 11946 13864
rect 12069 13855 12127 13861
rect 12069 13852 12081 13855
rect 11940 13824 12081 13852
rect 11940 13812 11946 13824
rect 12069 13821 12081 13824
rect 12115 13821 12127 13855
rect 12069 13815 12127 13821
rect 12342 13812 12348 13864
rect 12400 13852 12406 13864
rect 13924 13852 13952 13892
rect 15381 13889 15393 13892
rect 15427 13889 15439 13923
rect 15381 13883 15439 13889
rect 15470 13880 15476 13932
rect 15528 13920 15534 13932
rect 15933 13923 15991 13929
rect 15933 13920 15945 13923
rect 15528 13892 15945 13920
rect 15528 13880 15534 13892
rect 15933 13889 15945 13892
rect 15979 13889 15991 13923
rect 16393 13923 16451 13929
rect 16393 13920 16405 13923
rect 15933 13883 15991 13889
rect 16040 13892 16405 13920
rect 12400 13824 13952 13852
rect 14093 13855 14151 13861
rect 12400 13812 12406 13824
rect 14093 13821 14105 13855
rect 14139 13852 14151 13855
rect 14274 13852 14280 13864
rect 14139 13824 14280 13852
rect 14139 13821 14151 13824
rect 14093 13815 14151 13821
rect 14274 13812 14280 13824
rect 14332 13852 14338 13864
rect 15013 13855 15071 13861
rect 15013 13852 15025 13855
rect 14332 13824 15025 13852
rect 14332 13812 14338 13824
rect 15013 13821 15025 13824
rect 15059 13852 15071 13855
rect 15197 13855 15255 13861
rect 15197 13852 15209 13855
rect 15059 13824 15209 13852
rect 15059 13821 15071 13824
rect 15013 13815 15071 13821
rect 15197 13821 15209 13824
rect 15243 13821 15255 13855
rect 15197 13815 15255 13821
rect 15286 13812 15292 13864
rect 15344 13852 15350 13864
rect 15749 13855 15807 13861
rect 15749 13852 15761 13855
rect 15344 13824 15761 13852
rect 15344 13812 15350 13824
rect 15749 13821 15761 13824
rect 15795 13852 15807 13855
rect 16040 13852 16068 13892
rect 16393 13889 16405 13892
rect 16439 13889 16451 13923
rect 26712 13920 26740 14019
rect 27157 13923 27215 13929
rect 27157 13920 27169 13923
rect 26712 13892 27169 13920
rect 16393 13883 16451 13889
rect 27157 13889 27169 13892
rect 27203 13889 27215 13923
rect 27157 13883 27215 13889
rect 15795 13824 16068 13852
rect 16117 13855 16175 13861
rect 15795 13821 15807 13824
rect 15749 13815 15807 13821
rect 16117 13821 16129 13855
rect 16163 13852 16175 13855
rect 16482 13852 16488 13864
rect 16163 13824 16488 13852
rect 16163 13821 16175 13824
rect 16117 13815 16175 13821
rect 16482 13812 16488 13824
rect 16540 13812 16546 13864
rect 28350 13812 28356 13864
rect 28408 13812 28414 13864
rect 9692 13756 11192 13784
rect 11256 13756 12204 13784
rect 8812 13744 8818 13756
rect 11164 13728 11192 13756
rect 12176 13728 12204 13756
rect 8110 13676 8116 13728
rect 8168 13676 8174 13728
rect 8662 13676 8668 13728
rect 8720 13676 8726 13728
rect 9585 13719 9643 13725
rect 9585 13685 9597 13719
rect 9631 13716 9643 13719
rect 9674 13716 9680 13728
rect 9631 13688 9680 13716
rect 9631 13685 9643 13688
rect 9585 13679 9643 13685
rect 9674 13676 9680 13688
rect 9732 13676 9738 13728
rect 11146 13676 11152 13728
rect 11204 13676 11210 13728
rect 12158 13676 12164 13728
rect 12216 13716 12222 13728
rect 12434 13716 12440 13728
rect 12216 13688 12440 13716
rect 12216 13676 12222 13688
rect 12434 13676 12440 13688
rect 12492 13676 12498 13728
rect 1104 13626 28888 13648
rect 1104 13574 4423 13626
rect 4475 13574 4487 13626
rect 4539 13574 4551 13626
rect 4603 13574 4615 13626
rect 4667 13574 4679 13626
rect 4731 13574 11369 13626
rect 11421 13574 11433 13626
rect 11485 13574 11497 13626
rect 11549 13574 11561 13626
rect 11613 13574 11625 13626
rect 11677 13574 18315 13626
rect 18367 13574 18379 13626
rect 18431 13574 18443 13626
rect 18495 13574 18507 13626
rect 18559 13574 18571 13626
rect 18623 13574 25261 13626
rect 25313 13574 25325 13626
rect 25377 13574 25389 13626
rect 25441 13574 25453 13626
rect 25505 13574 25517 13626
rect 25569 13574 28888 13626
rect 1104 13552 28888 13574
rect 6730 13472 6736 13524
rect 6788 13512 6794 13524
rect 8754 13512 8760 13524
rect 6788 13484 8760 13512
rect 6788 13472 6794 13484
rect 8754 13472 8760 13484
rect 8812 13472 8818 13524
rect 9122 13472 9128 13524
rect 9180 13512 9186 13524
rect 9309 13515 9367 13521
rect 9309 13512 9321 13515
rect 9180 13484 9321 13512
rect 9180 13472 9186 13484
rect 9309 13481 9321 13484
rect 9355 13481 9367 13515
rect 26973 13515 27031 13521
rect 26973 13512 26985 13515
rect 9309 13475 9367 13481
rect 9416 13484 26985 13512
rect 1854 13404 1860 13456
rect 1912 13404 1918 13456
rect 7650 13404 7656 13456
rect 7708 13444 7714 13456
rect 8110 13444 8116 13456
rect 7708 13416 8116 13444
rect 7708 13404 7714 13416
rect 8110 13404 8116 13416
rect 8168 13444 8174 13456
rect 9416 13444 9444 13484
rect 26973 13481 26985 13484
rect 27019 13481 27031 13515
rect 26973 13475 27031 13481
rect 8168 13416 9444 13444
rect 8168 13404 8174 13416
rect 3970 13336 3976 13388
rect 4028 13376 4034 13388
rect 5261 13379 5319 13385
rect 5261 13376 5273 13379
rect 4028 13348 5273 13376
rect 4028 13336 4034 13348
rect 5261 13345 5273 13348
rect 5307 13345 5319 13379
rect 5261 13339 5319 13345
rect 6730 13336 6736 13388
rect 6788 13376 6794 13388
rect 7745 13379 7803 13385
rect 7745 13376 7757 13379
rect 6788 13348 7757 13376
rect 6788 13336 6794 13348
rect 7745 13345 7757 13348
rect 7791 13376 7803 13379
rect 8294 13376 8300 13388
rect 7791 13348 8300 13376
rect 7791 13345 7803 13348
rect 7745 13339 7803 13345
rect 8294 13336 8300 13348
rect 8352 13336 8358 13388
rect 8662 13336 8668 13388
rect 8720 13336 8726 13388
rect 9030 13336 9036 13388
rect 9088 13376 9094 13388
rect 9401 13379 9459 13385
rect 9401 13376 9413 13379
rect 9088 13348 9413 13376
rect 9088 13336 9094 13348
rect 9401 13345 9413 13348
rect 9447 13345 9459 13379
rect 9401 13339 9459 13345
rect 9677 13379 9735 13385
rect 9677 13345 9689 13379
rect 9723 13376 9735 13379
rect 9766 13376 9772 13388
rect 9723 13348 9772 13376
rect 9723 13345 9735 13348
rect 9677 13339 9735 13345
rect 9766 13336 9772 13348
rect 9824 13336 9830 13388
rect 11054 13336 11060 13388
rect 11112 13376 11118 13388
rect 11422 13376 11428 13388
rect 11112 13348 11428 13376
rect 11112 13336 11118 13348
rect 11422 13336 11428 13348
rect 11480 13336 11486 13388
rect 13722 13336 13728 13388
rect 13780 13376 13786 13388
rect 13780 13348 15700 13376
rect 13780 13336 13786 13348
rect 934 13268 940 13320
rect 992 13308 998 13320
rect 1397 13311 1455 13317
rect 1397 13308 1409 13311
rect 992 13280 1409 13308
rect 992 13268 998 13280
rect 1397 13277 1409 13280
rect 1443 13277 1455 13311
rect 1397 13271 1455 13277
rect 1673 13311 1731 13317
rect 1673 13277 1685 13311
rect 1719 13277 1731 13311
rect 1673 13271 1731 13277
rect 5445 13311 5503 13317
rect 5445 13277 5457 13311
rect 5491 13308 5503 13311
rect 5626 13308 5632 13320
rect 5491 13280 5632 13308
rect 5491 13277 5503 13280
rect 5445 13271 5503 13277
rect 1026 13200 1032 13252
rect 1084 13240 1090 13252
rect 1688 13240 1716 13271
rect 5626 13268 5632 13280
rect 5684 13268 5690 13320
rect 5718 13268 5724 13320
rect 5776 13268 5782 13320
rect 8386 13268 8392 13320
rect 8444 13308 8450 13320
rect 8941 13311 8999 13317
rect 8941 13308 8953 13311
rect 8444 13280 8953 13308
rect 8444 13268 8450 13280
rect 8941 13277 8953 13280
rect 8987 13277 8999 13311
rect 8941 13271 8999 13277
rect 9122 13268 9128 13320
rect 9180 13268 9186 13320
rect 11882 13268 11888 13320
rect 11940 13268 11946 13320
rect 15672 13317 15700 13348
rect 16022 13336 16028 13388
rect 16080 13376 16086 13388
rect 16669 13379 16727 13385
rect 16669 13376 16681 13379
rect 16080 13348 16681 13376
rect 16080 13336 16086 13348
rect 16669 13345 16681 13348
rect 16715 13345 16727 13379
rect 16669 13339 16727 13345
rect 15565 13311 15623 13317
rect 15565 13277 15577 13311
rect 15611 13277 15623 13311
rect 15565 13271 15623 13277
rect 15657 13311 15715 13317
rect 15657 13277 15669 13311
rect 15703 13277 15715 13311
rect 15657 13271 15715 13277
rect 1084 13212 1716 13240
rect 1084 13200 1090 13212
rect 5994 13200 6000 13252
rect 6052 13200 6058 13252
rect 7374 13240 7380 13252
rect 7222 13212 7380 13240
rect 7374 13200 7380 13212
rect 7432 13200 7438 13252
rect 10686 13200 10692 13252
rect 10744 13200 10750 13252
rect 12158 13200 12164 13252
rect 12216 13200 12222 13252
rect 13446 13240 13452 13252
rect 13386 13212 13452 13240
rect 13446 13200 13452 13212
rect 13504 13200 13510 13252
rect 13909 13243 13967 13249
rect 13909 13209 13921 13243
rect 13955 13240 13967 13243
rect 15381 13243 15439 13249
rect 15381 13240 15393 13243
rect 13955 13212 15393 13240
rect 13955 13209 13967 13212
rect 13909 13203 13967 13209
rect 15381 13209 15393 13212
rect 15427 13240 15439 13243
rect 15580 13240 15608 13271
rect 15746 13268 15752 13320
rect 15804 13308 15810 13320
rect 16209 13311 16267 13317
rect 16209 13308 16221 13311
rect 15804 13280 16221 13308
rect 15804 13268 15810 13280
rect 16209 13277 16221 13280
rect 16255 13277 16267 13311
rect 26988 13308 27016 13475
rect 27157 13311 27215 13317
rect 27157 13308 27169 13311
rect 26988 13280 27169 13308
rect 16209 13271 16267 13277
rect 27157 13277 27169 13280
rect 27203 13277 27215 13311
rect 27157 13271 27215 13277
rect 25682 13240 25688 13252
rect 15427 13212 25688 13240
rect 15427 13209 15439 13212
rect 15381 13203 15439 13209
rect 1578 13132 1584 13184
rect 1636 13132 1642 13184
rect 5629 13175 5687 13181
rect 5629 13141 5641 13175
rect 5675 13172 5687 13175
rect 6822 13172 6828 13184
rect 5675 13144 6828 13172
rect 5675 13141 5687 13144
rect 5629 13135 5687 13141
rect 6822 13132 6828 13144
rect 6880 13132 6886 13184
rect 8113 13175 8171 13181
rect 8113 13141 8125 13175
rect 8159 13172 8171 13175
rect 8662 13172 8668 13184
rect 8159 13144 8668 13172
rect 8159 13141 8171 13144
rect 8113 13135 8171 13141
rect 8662 13132 8668 13144
rect 8720 13132 8726 13184
rect 12894 13132 12900 13184
rect 12952 13172 12958 13184
rect 13924 13172 13952 13203
rect 25682 13200 25688 13212
rect 25740 13200 25746 13252
rect 28350 13200 28356 13252
rect 28408 13200 28414 13252
rect 12952 13144 13952 13172
rect 12952 13132 12958 13144
rect 15838 13132 15844 13184
rect 15896 13132 15902 13184
rect 16390 13132 16396 13184
rect 16448 13132 16454 13184
rect 1104 13082 29048 13104
rect 1104 13030 7896 13082
rect 7948 13030 7960 13082
rect 8012 13030 8024 13082
rect 8076 13030 8088 13082
rect 8140 13030 8152 13082
rect 8204 13030 14842 13082
rect 14894 13030 14906 13082
rect 14958 13030 14970 13082
rect 15022 13030 15034 13082
rect 15086 13030 15098 13082
rect 15150 13030 21788 13082
rect 21840 13030 21852 13082
rect 21904 13030 21916 13082
rect 21968 13030 21980 13082
rect 22032 13030 22044 13082
rect 22096 13030 28734 13082
rect 28786 13030 28798 13082
rect 28850 13030 28862 13082
rect 28914 13030 28926 13082
rect 28978 13030 28990 13082
rect 29042 13030 29048 13082
rect 1104 13008 29048 13030
rect 1581 12971 1639 12977
rect 1581 12937 1593 12971
rect 1627 12968 1639 12971
rect 5537 12971 5595 12977
rect 1627 12940 2774 12968
rect 1627 12937 1639 12940
rect 1581 12931 1639 12937
rect 934 12792 940 12844
rect 992 12832 998 12844
rect 1397 12835 1455 12841
rect 1397 12832 1409 12835
rect 992 12804 1409 12832
rect 992 12792 998 12804
rect 1397 12801 1409 12804
rect 1443 12801 1455 12835
rect 1397 12795 1455 12801
rect 1670 12792 1676 12844
rect 1728 12792 1734 12844
rect 1854 12656 1860 12708
rect 1912 12656 1918 12708
rect 2746 12696 2774 12940
rect 5537 12937 5549 12971
rect 5583 12968 5595 12971
rect 5994 12968 6000 12980
rect 5583 12940 6000 12968
rect 5583 12937 5595 12940
rect 5537 12931 5595 12937
rect 5994 12928 6000 12940
rect 6052 12928 6058 12980
rect 6730 12928 6736 12980
rect 6788 12928 6794 12980
rect 6822 12928 6828 12980
rect 6880 12928 6886 12980
rect 7374 12928 7380 12980
rect 7432 12928 7438 12980
rect 7466 12928 7472 12980
rect 7524 12968 7530 12980
rect 7561 12971 7619 12977
rect 7561 12968 7573 12971
rect 7524 12940 7573 12968
rect 7524 12928 7530 12940
rect 7561 12937 7573 12940
rect 7607 12968 7619 12971
rect 7650 12968 7656 12980
rect 7607 12940 7656 12968
rect 7607 12937 7619 12940
rect 7561 12931 7619 12937
rect 7650 12928 7656 12940
rect 7708 12928 7714 12980
rect 7834 12928 7840 12980
rect 7892 12968 7898 12980
rect 7892 12940 8340 12968
rect 7892 12928 7898 12940
rect 5626 12860 5632 12912
rect 5684 12900 5690 12912
rect 5902 12900 5908 12912
rect 5684 12872 5908 12900
rect 5684 12860 5690 12872
rect 5902 12860 5908 12872
rect 5960 12860 5966 12912
rect 6748 12900 6776 12928
rect 6012 12872 6776 12900
rect 7392 12900 7420 12928
rect 8113 12903 8171 12909
rect 8113 12900 8125 12903
rect 7392 12872 8125 12900
rect 5445 12835 5503 12841
rect 5445 12801 5457 12835
rect 5491 12832 5503 12835
rect 6012 12832 6040 12872
rect 8113 12869 8125 12872
rect 8159 12869 8171 12903
rect 8113 12863 8171 12869
rect 5491 12804 6040 12832
rect 6104 12804 7604 12832
rect 5491 12801 5503 12804
rect 5445 12795 5503 12801
rect 6104 12696 6132 12804
rect 6181 12767 6239 12773
rect 6181 12733 6193 12767
rect 6227 12733 6239 12767
rect 6181 12727 6239 12733
rect 7009 12767 7067 12773
rect 7009 12733 7021 12767
rect 7055 12764 7067 12767
rect 7098 12764 7104 12776
rect 7055 12736 7104 12764
rect 7055 12733 7067 12736
rect 7009 12727 7067 12733
rect 2746 12668 6132 12696
rect 6196 12696 6224 12727
rect 7098 12724 7104 12736
rect 7156 12764 7162 12776
rect 7285 12767 7343 12773
rect 7285 12764 7297 12767
rect 7156 12736 7297 12764
rect 7156 12724 7162 12736
rect 7285 12733 7297 12736
rect 7331 12764 7343 12767
rect 7374 12764 7380 12776
rect 7331 12736 7380 12764
rect 7331 12733 7343 12736
rect 7285 12727 7343 12733
rect 7374 12724 7380 12736
rect 7432 12724 7438 12776
rect 7469 12767 7527 12773
rect 7469 12733 7481 12767
rect 7515 12733 7527 12767
rect 7469 12727 7527 12733
rect 6365 12699 6423 12705
rect 6365 12696 6377 12699
rect 6196 12668 6377 12696
rect 6365 12665 6377 12668
rect 6411 12665 6423 12699
rect 6365 12659 6423 12665
rect 5994 12588 6000 12640
rect 6052 12628 6058 12640
rect 7484 12628 7512 12727
rect 6052 12600 7512 12628
rect 7576 12628 7604 12804
rect 8018 12792 8024 12844
rect 8076 12832 8082 12844
rect 8312 12841 8340 12940
rect 8754 12928 8760 12980
rect 8812 12968 8818 12980
rect 8812 12940 10364 12968
rect 8812 12928 8818 12940
rect 8573 12903 8631 12909
rect 8573 12869 8585 12903
rect 8619 12900 8631 12903
rect 8662 12900 8668 12912
rect 8619 12872 8668 12900
rect 8619 12869 8631 12872
rect 8573 12863 8631 12869
rect 8662 12860 8668 12872
rect 8720 12860 8726 12912
rect 10336 12900 10364 12940
rect 10410 12928 10416 12980
rect 10468 12928 10474 12980
rect 10686 12928 10692 12980
rect 10744 12968 10750 12980
rect 10965 12971 11023 12977
rect 10965 12968 10977 12971
rect 10744 12940 10977 12968
rect 10744 12928 10750 12940
rect 10965 12937 10977 12940
rect 11011 12937 11023 12971
rect 10965 12931 11023 12937
rect 12158 12928 12164 12980
rect 12216 12968 12222 12980
rect 13081 12971 13139 12977
rect 13081 12968 13093 12971
rect 12216 12940 13093 12968
rect 12216 12928 12222 12940
rect 13081 12937 13093 12940
rect 13127 12937 13139 12971
rect 13081 12931 13139 12937
rect 13446 12928 13452 12980
rect 13504 12968 13510 12980
rect 13909 12971 13967 12977
rect 13909 12968 13921 12971
rect 13504 12940 13921 12968
rect 13504 12928 13510 12940
rect 13909 12937 13921 12940
rect 13955 12937 13967 12971
rect 13909 12931 13967 12937
rect 14369 12971 14427 12977
rect 14369 12937 14381 12971
rect 14415 12968 14427 12971
rect 14734 12968 14740 12980
rect 14415 12940 14740 12968
rect 14415 12937 14427 12940
rect 14369 12931 14427 12937
rect 10336 12872 10732 12900
rect 8197 12835 8255 12841
rect 8076 12830 8156 12832
rect 8197 12830 8209 12835
rect 8076 12804 8209 12830
rect 8076 12792 8082 12804
rect 8128 12802 8209 12804
rect 8197 12801 8209 12802
rect 8243 12801 8255 12835
rect 8197 12795 8255 12801
rect 8297 12835 8355 12841
rect 8297 12801 8309 12835
rect 8343 12801 8355 12835
rect 8297 12795 8355 12801
rect 9674 12792 9680 12844
rect 9732 12792 9738 12844
rect 10594 12792 10600 12844
rect 10652 12792 10658 12844
rect 10704 12841 10732 12872
rect 10796 12872 13768 12900
rect 10689 12835 10747 12841
rect 10689 12801 10701 12835
rect 10735 12801 10747 12835
rect 10689 12795 10747 12801
rect 10318 12724 10324 12776
rect 10376 12764 10382 12776
rect 10796 12764 10824 12872
rect 11054 12792 11060 12844
rect 11112 12792 11118 12844
rect 12161 12835 12219 12841
rect 12161 12801 12173 12835
rect 12207 12832 12219 12835
rect 12452 12832 12572 12838
rect 12621 12835 12679 12841
rect 12621 12832 12633 12835
rect 12207 12810 12633 12832
rect 12207 12804 12480 12810
rect 12544 12804 12633 12810
rect 12207 12801 12219 12804
rect 12161 12795 12219 12801
rect 12621 12801 12633 12804
rect 12667 12832 12679 12835
rect 12667 12804 12721 12832
rect 12667 12801 12679 12804
rect 12621 12795 12679 12801
rect 10376 12736 10824 12764
rect 10376 12724 10382 12736
rect 12434 12724 12440 12776
rect 12492 12724 12498 12776
rect 12526 12724 12532 12776
rect 12584 12724 12590 12776
rect 12636 12764 12664 12795
rect 12894 12764 12900 12776
rect 12636 12736 12900 12764
rect 12894 12724 12900 12736
rect 12952 12724 12958 12776
rect 13633 12767 13691 12773
rect 13633 12764 13645 12767
rect 13004 12736 13645 12764
rect 7926 12656 7932 12708
rect 7984 12656 7990 12708
rect 9766 12656 9772 12708
rect 9824 12656 9830 12708
rect 13004 12705 13032 12736
rect 13633 12733 13645 12736
rect 13679 12733 13691 12767
rect 13740 12764 13768 12872
rect 13814 12792 13820 12844
rect 13872 12832 13878 12844
rect 14001 12835 14059 12841
rect 14001 12832 14013 12835
rect 13872 12804 14013 12832
rect 13872 12792 13878 12804
rect 14001 12801 14013 12804
rect 14047 12832 14059 12835
rect 14384 12832 14412 12931
rect 14734 12928 14740 12940
rect 14792 12928 14798 12980
rect 16390 12928 16396 12980
rect 16448 12968 16454 12980
rect 22830 12968 22836 12980
rect 16448 12940 22836 12968
rect 16448 12928 16454 12940
rect 22830 12928 22836 12940
rect 22888 12928 22894 12980
rect 14642 12860 14648 12912
rect 14700 12900 14706 12912
rect 14921 12903 14979 12909
rect 14921 12900 14933 12903
rect 14700 12872 14933 12900
rect 14700 12860 14706 12872
rect 14921 12869 14933 12872
rect 14967 12869 14979 12903
rect 17770 12900 17776 12912
rect 14921 12863 14979 12869
rect 15212 12872 17776 12900
rect 14047 12804 14412 12832
rect 14936 12832 14964 12863
rect 15105 12835 15163 12841
rect 15105 12832 15117 12835
rect 14936 12804 15117 12832
rect 14047 12801 14059 12804
rect 14001 12795 14059 12801
rect 15105 12801 15117 12804
rect 15151 12801 15163 12835
rect 15105 12795 15163 12801
rect 15212 12764 15240 12872
rect 17770 12860 17776 12872
rect 17828 12860 17834 12912
rect 15286 12792 15292 12844
rect 15344 12792 15350 12844
rect 16114 12792 16120 12844
rect 16172 12792 16178 12844
rect 13740 12736 15240 12764
rect 15841 12767 15899 12773
rect 13633 12727 13691 12733
rect 15841 12733 15853 12767
rect 15887 12764 15899 12767
rect 15933 12767 15991 12773
rect 15933 12764 15945 12767
rect 15887 12736 15945 12764
rect 15887 12733 15899 12736
rect 15841 12727 15899 12733
rect 15933 12733 15945 12736
rect 15979 12764 15991 12767
rect 25774 12764 25780 12776
rect 15979 12736 25780 12764
rect 15979 12733 15991 12736
rect 15933 12727 15991 12733
rect 12989 12699 13047 12705
rect 12989 12665 13001 12699
rect 13035 12665 13047 12699
rect 15856 12696 15884 12727
rect 25774 12724 25780 12736
rect 25832 12724 25838 12776
rect 12989 12659 13047 12665
rect 14200 12668 15884 12696
rect 9784 12628 9812 12656
rect 7576 12600 9812 12628
rect 6052 12588 6058 12600
rect 11422 12588 11428 12640
rect 11480 12628 11486 12640
rect 14200 12628 14228 12668
rect 11480 12600 14228 12628
rect 11480 12588 11486 12600
rect 15470 12588 15476 12640
rect 15528 12588 15534 12640
rect 16301 12631 16359 12637
rect 16301 12597 16313 12631
rect 16347 12628 16359 12631
rect 17218 12628 17224 12640
rect 16347 12600 17224 12628
rect 16347 12597 16359 12600
rect 16301 12591 16359 12597
rect 17218 12588 17224 12600
rect 17276 12588 17282 12640
rect 1104 12538 28888 12560
rect 1104 12486 4423 12538
rect 4475 12486 4487 12538
rect 4539 12486 4551 12538
rect 4603 12486 4615 12538
rect 4667 12486 4679 12538
rect 4731 12486 11369 12538
rect 11421 12486 11433 12538
rect 11485 12486 11497 12538
rect 11549 12486 11561 12538
rect 11613 12486 11625 12538
rect 11677 12486 18315 12538
rect 18367 12486 18379 12538
rect 18431 12486 18443 12538
rect 18495 12486 18507 12538
rect 18559 12486 18571 12538
rect 18623 12486 25261 12538
rect 25313 12486 25325 12538
rect 25377 12486 25389 12538
rect 25441 12486 25453 12538
rect 25505 12486 25517 12538
rect 25569 12486 28888 12538
rect 1104 12464 28888 12486
rect 2746 12396 9996 12424
rect 1581 12359 1639 12365
rect 1581 12325 1593 12359
rect 1627 12356 1639 12359
rect 2746 12356 2774 12396
rect 1627 12328 2774 12356
rect 1627 12325 1639 12328
rect 1581 12319 1639 12325
rect 5718 12316 5724 12368
rect 5776 12356 5782 12368
rect 7834 12356 7840 12368
rect 5776 12328 7840 12356
rect 5776 12316 5782 12328
rect 7834 12316 7840 12328
rect 7892 12356 7898 12368
rect 9030 12356 9036 12368
rect 7892 12328 9036 12356
rect 7892 12316 7898 12328
rect 9030 12316 9036 12328
rect 9088 12316 9094 12368
rect 7006 12248 7012 12300
rect 7064 12288 7070 12300
rect 7374 12288 7380 12300
rect 7064 12260 7380 12288
rect 7064 12248 7070 12260
rect 7374 12248 7380 12260
rect 7432 12248 7438 12300
rect 7484 12260 8240 12288
rect 934 12180 940 12232
rect 992 12220 998 12232
rect 1397 12223 1455 12229
rect 1397 12220 1409 12223
rect 992 12192 1409 12220
rect 992 12180 998 12192
rect 1397 12189 1409 12192
rect 1443 12189 1455 12223
rect 1397 12183 1455 12189
rect 1673 12223 1731 12229
rect 1673 12189 1685 12223
rect 1719 12189 1731 12223
rect 1673 12183 1731 12189
rect 1026 12112 1032 12164
rect 1084 12152 1090 12164
rect 1688 12152 1716 12183
rect 6638 12180 6644 12232
rect 6696 12220 6702 12232
rect 7484 12220 7512 12260
rect 8113 12223 8171 12229
rect 8113 12220 8125 12223
rect 6696 12192 7512 12220
rect 8036 12192 8125 12220
rect 6696 12180 6702 12192
rect 1084 12124 1716 12152
rect 7009 12155 7067 12161
rect 1084 12112 1090 12124
rect 7009 12121 7021 12155
rect 7055 12152 7067 12155
rect 7742 12152 7748 12164
rect 7055 12124 7748 12152
rect 7055 12121 7067 12124
rect 7009 12115 7067 12121
rect 7742 12112 7748 12124
rect 7800 12112 7806 12164
rect 1854 12044 1860 12096
rect 1912 12044 1918 12096
rect 5166 12044 5172 12096
rect 5224 12044 5230 12096
rect 6822 12044 6828 12096
rect 6880 12084 6886 12096
rect 7561 12087 7619 12093
rect 7561 12084 7573 12087
rect 6880 12056 7573 12084
rect 6880 12044 6886 12056
rect 7561 12053 7573 12056
rect 7607 12053 7619 12087
rect 7561 12047 7619 12053
rect 7653 12087 7711 12093
rect 7653 12053 7665 12087
rect 7699 12084 7711 12087
rect 7926 12084 7932 12096
rect 7699 12056 7932 12084
rect 7699 12053 7711 12056
rect 7653 12047 7711 12053
rect 7926 12044 7932 12056
rect 7984 12044 7990 12096
rect 8036 12093 8064 12192
rect 8113 12189 8125 12192
rect 8159 12189 8171 12223
rect 8113 12183 8171 12189
rect 8212 12152 8240 12260
rect 8754 12248 8760 12300
rect 8812 12288 8818 12300
rect 9493 12291 9551 12297
rect 9493 12288 9505 12291
rect 8812 12260 9505 12288
rect 8812 12248 8818 12260
rect 9493 12257 9505 12260
rect 9539 12257 9551 12291
rect 9493 12251 9551 12257
rect 8941 12223 8999 12229
rect 8941 12189 8953 12223
rect 8987 12189 8999 12223
rect 8941 12183 8999 12189
rect 8956 12152 8984 12183
rect 9858 12180 9864 12232
rect 9916 12180 9922 12232
rect 9968 12229 9996 12396
rect 15194 12384 15200 12436
rect 15252 12384 15258 12436
rect 16206 12384 16212 12436
rect 16264 12424 16270 12436
rect 16301 12427 16359 12433
rect 16301 12424 16313 12427
rect 16264 12396 16313 12424
rect 16264 12384 16270 12396
rect 16301 12393 16313 12396
rect 16347 12424 16359 12427
rect 16347 12396 16528 12424
rect 16347 12393 16359 12396
rect 16301 12387 16359 12393
rect 10137 12359 10195 12365
rect 10137 12325 10149 12359
rect 10183 12356 10195 12359
rect 10594 12356 10600 12368
rect 10183 12328 10600 12356
rect 10183 12325 10195 12328
rect 10137 12319 10195 12325
rect 10594 12316 10600 12328
rect 10652 12316 10658 12368
rect 11425 12359 11483 12365
rect 11425 12325 11437 12359
rect 11471 12325 11483 12359
rect 11425 12319 11483 12325
rect 10781 12291 10839 12297
rect 10781 12257 10793 12291
rect 10827 12288 10839 12291
rect 11440 12288 11468 12319
rect 11790 12316 11796 12368
rect 11848 12356 11854 12368
rect 12989 12359 13047 12365
rect 11848 12328 12020 12356
rect 11848 12316 11854 12328
rect 10827 12260 11468 12288
rect 10827 12257 10839 12260
rect 10781 12251 10839 12257
rect 11514 12248 11520 12300
rect 11572 12288 11578 12300
rect 11992 12297 12020 12328
rect 12360 12328 12664 12356
rect 12360 12300 12388 12328
rect 11885 12291 11943 12297
rect 11885 12288 11897 12291
rect 11572 12260 11897 12288
rect 11572 12248 11578 12260
rect 11885 12257 11897 12260
rect 11931 12257 11943 12291
rect 11885 12251 11943 12257
rect 11977 12291 12035 12297
rect 11977 12257 11989 12291
rect 12023 12257 12035 12291
rect 11977 12251 12035 12257
rect 12342 12248 12348 12300
rect 12400 12248 12406 12300
rect 12434 12248 12440 12300
rect 12492 12248 12498 12300
rect 9953 12223 10011 12229
rect 9953 12189 9965 12223
rect 9999 12189 10011 12223
rect 9953 12183 10011 12189
rect 10505 12223 10563 12229
rect 10505 12189 10517 12223
rect 10551 12220 10563 12223
rect 11054 12220 11060 12232
rect 10551 12192 11060 12220
rect 10551 12189 10563 12192
rect 10505 12183 10563 12189
rect 11054 12180 11060 12192
rect 11112 12180 11118 12232
rect 11333 12223 11391 12229
rect 11333 12189 11345 12223
rect 11379 12220 11391 12223
rect 11422 12220 11428 12232
rect 11379 12192 11428 12220
rect 11379 12189 11391 12192
rect 11333 12183 11391 12189
rect 11422 12180 11428 12192
rect 11480 12180 11486 12232
rect 12529 12223 12587 12229
rect 12529 12220 12541 12223
rect 11532 12192 12541 12220
rect 8212 12124 8984 12152
rect 9306 12112 9312 12164
rect 9364 12152 9370 12164
rect 11532 12152 11560 12192
rect 12529 12189 12541 12192
rect 12575 12189 12587 12223
rect 12636 12220 12664 12328
rect 12989 12325 13001 12359
rect 13035 12325 13047 12359
rect 12989 12319 13047 12325
rect 13004 12288 13032 12319
rect 13633 12291 13691 12297
rect 13633 12288 13645 12291
rect 13004 12260 13645 12288
rect 13633 12257 13645 12260
rect 13679 12257 13691 12291
rect 15212 12288 15240 12384
rect 16500 12297 16528 12396
rect 16666 12384 16672 12436
rect 16724 12424 16730 12436
rect 23474 12424 23480 12436
rect 16724 12396 23480 12424
rect 16724 12384 16730 12396
rect 23474 12384 23480 12396
rect 23532 12384 23538 12436
rect 15381 12291 15439 12297
rect 15381 12288 15393 12291
rect 15212 12260 15393 12288
rect 13633 12251 13691 12257
rect 15381 12257 15393 12260
rect 15427 12257 15439 12291
rect 15381 12251 15439 12257
rect 16485 12291 16543 12297
rect 16485 12257 16497 12291
rect 16531 12257 16543 12291
rect 16485 12251 16543 12257
rect 14093 12223 14151 12229
rect 14093 12220 14105 12223
rect 12636 12192 14105 12220
rect 12529 12183 12587 12189
rect 14093 12189 14105 12192
rect 14139 12189 14151 12223
rect 14093 12183 14151 12189
rect 15562 12180 15568 12232
rect 15620 12180 15626 12232
rect 16669 12223 16727 12229
rect 16669 12220 16681 12223
rect 15672 12192 16681 12220
rect 9364 12124 11560 12152
rect 11793 12155 11851 12161
rect 9364 12112 9370 12124
rect 11793 12121 11805 12155
rect 11839 12152 11851 12155
rect 12621 12155 12679 12161
rect 11839 12124 12572 12152
rect 11839 12121 11851 12124
rect 11793 12115 11851 12121
rect 8021 12087 8079 12093
rect 8021 12053 8033 12087
rect 8067 12053 8079 12087
rect 8021 12047 8079 12053
rect 8662 12044 8668 12096
rect 8720 12084 8726 12096
rect 8757 12087 8815 12093
rect 8757 12084 8769 12087
rect 8720 12056 8769 12084
rect 8720 12044 8726 12056
rect 8757 12053 8769 12056
rect 8803 12053 8815 12087
rect 8757 12047 8815 12053
rect 8846 12044 8852 12096
rect 8904 12084 8910 12096
rect 9582 12084 9588 12096
rect 8904 12056 9588 12084
rect 8904 12044 8910 12056
rect 9582 12044 9588 12056
rect 9640 12044 9646 12096
rect 10410 12044 10416 12096
rect 10468 12044 10474 12096
rect 11238 12044 11244 12096
rect 11296 12084 11302 12096
rect 12434 12084 12440 12096
rect 11296 12056 12440 12084
rect 11296 12044 11302 12056
rect 12434 12044 12440 12056
rect 12492 12044 12498 12096
rect 12544 12084 12572 12124
rect 12621 12121 12633 12155
rect 12667 12152 12679 12155
rect 12667 12124 13676 12152
rect 12667 12121 12679 12124
rect 12621 12115 12679 12121
rect 13648 12096 13676 12124
rect 13722 12112 13728 12164
rect 13780 12152 13786 12164
rect 15672 12152 15700 12192
rect 16669 12189 16681 12192
rect 16715 12189 16727 12223
rect 27157 12223 27215 12229
rect 27157 12220 27169 12223
rect 16669 12183 16727 12189
rect 22066 12192 27169 12220
rect 13780 12124 15700 12152
rect 15749 12155 15807 12161
rect 13780 12112 13786 12124
rect 15749 12121 15761 12155
rect 15795 12152 15807 12155
rect 20070 12152 20076 12164
rect 15795 12124 20076 12152
rect 15795 12121 15807 12124
rect 15749 12115 15807 12121
rect 20070 12112 20076 12124
rect 20128 12112 20134 12164
rect 20162 12112 20168 12164
rect 20220 12152 20226 12164
rect 22066 12152 22094 12192
rect 27157 12189 27169 12192
rect 27203 12189 27215 12223
rect 27157 12183 27215 12189
rect 20220 12124 22094 12152
rect 20220 12112 20226 12124
rect 28350 12112 28356 12164
rect 28408 12112 28414 12164
rect 12986 12084 12992 12096
rect 12544 12056 12992 12084
rect 12986 12044 12992 12056
rect 13044 12044 13050 12096
rect 13078 12044 13084 12096
rect 13136 12044 13142 12096
rect 13630 12044 13636 12096
rect 13688 12044 13694 12096
rect 14182 12044 14188 12096
rect 14240 12044 14246 12096
rect 16853 12087 16911 12093
rect 16853 12053 16865 12087
rect 16899 12084 16911 12087
rect 18874 12084 18880 12096
rect 16899 12056 18880 12084
rect 16899 12053 16911 12056
rect 16853 12047 16911 12053
rect 18874 12044 18880 12056
rect 18932 12044 18938 12096
rect 1104 11994 29048 12016
rect 1104 11942 7896 11994
rect 7948 11942 7960 11994
rect 8012 11942 8024 11994
rect 8076 11942 8088 11994
rect 8140 11942 8152 11994
rect 8204 11942 14842 11994
rect 14894 11942 14906 11994
rect 14958 11942 14970 11994
rect 15022 11942 15034 11994
rect 15086 11942 15098 11994
rect 15150 11942 21788 11994
rect 21840 11942 21852 11994
rect 21904 11942 21916 11994
rect 21968 11942 21980 11994
rect 22032 11942 22044 11994
rect 22096 11942 28734 11994
rect 28786 11942 28798 11994
rect 28850 11942 28862 11994
rect 28914 11942 28926 11994
rect 28978 11942 28990 11994
rect 29042 11942 29048 11994
rect 1104 11920 29048 11942
rect 5994 11840 6000 11892
rect 6052 11840 6058 11892
rect 6822 11840 6828 11892
rect 6880 11840 6886 11892
rect 8018 11880 8024 11892
rect 7392 11852 8024 11880
rect 7392 11824 7420 11852
rect 8018 11840 8024 11852
rect 8076 11840 8082 11892
rect 8846 11880 8852 11892
rect 8312 11852 8852 11880
rect 3602 11772 3608 11824
rect 3660 11812 3666 11824
rect 6914 11812 6920 11824
rect 3660 11784 6500 11812
rect 3660 11772 3666 11784
rect 934 11704 940 11756
rect 992 11744 998 11756
rect 1397 11747 1455 11753
rect 1397 11744 1409 11747
rect 992 11716 1409 11744
rect 992 11704 998 11716
rect 1397 11713 1409 11716
rect 1443 11713 1455 11747
rect 1397 11707 1455 11713
rect 1673 11747 1731 11753
rect 1673 11713 1685 11747
rect 1719 11713 1731 11747
rect 1673 11707 1731 11713
rect 1026 11636 1032 11688
rect 1084 11676 1090 11688
rect 1688 11676 1716 11707
rect 3786 11704 3792 11756
rect 3844 11744 3850 11756
rect 5629 11747 5687 11753
rect 5629 11744 5641 11747
rect 3844 11716 5641 11744
rect 3844 11704 3850 11716
rect 5629 11713 5641 11716
rect 5675 11713 5687 11747
rect 5629 11707 5687 11713
rect 5813 11747 5871 11753
rect 5813 11713 5825 11747
rect 5859 11744 5871 11747
rect 6362 11744 6368 11756
rect 5859 11716 6368 11744
rect 5859 11713 5871 11716
rect 5813 11707 5871 11713
rect 6362 11704 6368 11716
rect 6420 11704 6426 11756
rect 6472 11753 6500 11784
rect 6656 11784 6920 11812
rect 6656 11753 6684 11784
rect 6914 11772 6920 11784
rect 6972 11772 6978 11824
rect 7374 11772 7380 11824
rect 7432 11772 7438 11824
rect 8312 11812 8340 11852
rect 8846 11840 8852 11852
rect 8904 11840 8910 11892
rect 9861 11883 9919 11889
rect 8956 11852 9444 11880
rect 8234 11784 8340 11812
rect 8754 11772 8760 11824
rect 8812 11812 8818 11824
rect 8956 11812 8984 11852
rect 8812 11784 8984 11812
rect 8812 11772 8818 11784
rect 6457 11747 6515 11753
rect 6457 11713 6469 11747
rect 6503 11713 6515 11747
rect 6457 11707 6515 11713
rect 6641 11747 6699 11753
rect 6641 11713 6653 11747
rect 6687 11713 6699 11747
rect 6641 11707 6699 11713
rect 9217 11748 9275 11753
rect 9416 11748 9444 11852
rect 9861 11849 9873 11883
rect 9907 11880 9919 11883
rect 10042 11880 10048 11892
rect 9907 11852 10048 11880
rect 9907 11849 9919 11852
rect 9861 11843 9919 11849
rect 10042 11840 10048 11852
rect 10100 11840 10106 11892
rect 10410 11840 10416 11892
rect 10468 11840 10474 11892
rect 11514 11840 11520 11892
rect 11572 11840 11578 11892
rect 13078 11880 13084 11892
rect 12406 11852 13084 11880
rect 9582 11772 9588 11824
rect 9640 11812 9646 11824
rect 10428 11812 10456 11840
rect 11532 11812 11560 11840
rect 9640 11784 10456 11812
rect 10796 11784 11560 11812
rect 12253 11815 12311 11821
rect 9640 11772 9646 11784
rect 9217 11747 9444 11748
rect 9217 11713 9229 11747
rect 9263 11720 9444 11747
rect 9263 11713 9275 11720
rect 9217 11707 9275 11713
rect 9490 11704 9496 11756
rect 9548 11704 9554 11756
rect 9858 11704 9864 11756
rect 9916 11744 9922 11756
rect 10321 11747 10379 11753
rect 10321 11744 10333 11747
rect 9916 11716 10333 11744
rect 9916 11704 9922 11716
rect 10321 11713 10333 11716
rect 10367 11713 10379 11747
rect 10321 11707 10379 11713
rect 1084 11648 1716 11676
rect 6917 11679 6975 11685
rect 1084 11636 1090 11648
rect 6917 11645 6929 11679
rect 6963 11676 6975 11679
rect 7926 11676 7932 11688
rect 6963 11648 7932 11676
rect 6963 11645 6975 11648
rect 6917 11639 6975 11645
rect 7926 11636 7932 11648
rect 7984 11676 7990 11688
rect 8202 11676 8208 11688
rect 7984 11648 8208 11676
rect 7984 11636 7990 11648
rect 8202 11636 8208 11648
rect 8260 11636 8266 11688
rect 8662 11636 8668 11688
rect 8720 11636 8726 11688
rect 8941 11679 8999 11685
rect 8941 11645 8953 11679
rect 8987 11645 8999 11679
rect 8941 11639 8999 11645
rect 9033 11679 9091 11685
rect 9033 11645 9045 11679
rect 9079 11676 9091 11679
rect 9508 11676 9536 11704
rect 10689 11679 10747 11685
rect 10689 11676 10701 11679
rect 9079 11648 9168 11676
rect 9079 11645 9091 11648
rect 9033 11639 9091 11645
rect 1581 11611 1639 11617
rect 1581 11577 1593 11611
rect 1627 11608 1639 11611
rect 1627 11580 7696 11608
rect 1627 11577 1639 11580
rect 1581 11571 1639 11577
rect 1854 11500 1860 11552
rect 1912 11500 1918 11552
rect 7668 11540 7696 11580
rect 8662 11540 8668 11552
rect 7668 11512 8668 11540
rect 8662 11500 8668 11512
rect 8720 11500 8726 11552
rect 8956 11540 8984 11639
rect 9140 11608 9168 11648
rect 9508 11648 10701 11676
rect 9508 11608 9536 11648
rect 10689 11645 10701 11648
rect 10735 11645 10747 11679
rect 10689 11639 10747 11645
rect 9140 11580 9536 11608
rect 9582 11568 9588 11620
rect 9640 11608 9646 11620
rect 10796 11608 10824 11784
rect 12253 11781 12265 11815
rect 12299 11812 12311 11815
rect 12406 11812 12434 11852
rect 13078 11840 13084 11852
rect 13136 11840 13142 11892
rect 16666 11840 16672 11892
rect 16724 11840 16730 11892
rect 17681 11883 17739 11889
rect 17681 11849 17693 11883
rect 17727 11880 17739 11883
rect 17770 11880 17776 11892
rect 17727 11852 17776 11880
rect 17727 11849 17739 11852
rect 17681 11843 17739 11849
rect 14182 11812 14188 11824
rect 12299 11784 12434 11812
rect 13478 11784 14188 11812
rect 12299 11781 12311 11784
rect 12253 11775 12311 11781
rect 14182 11772 14188 11784
rect 14240 11772 14246 11824
rect 11054 11704 11060 11756
rect 11112 11744 11118 11756
rect 11701 11747 11759 11753
rect 11701 11744 11713 11747
rect 11112 11716 11713 11744
rect 11112 11704 11118 11716
rect 11701 11713 11713 11716
rect 11747 11713 11759 11747
rect 11701 11707 11759 11713
rect 11422 11636 11428 11688
rect 11480 11636 11486 11688
rect 11716 11676 11744 11707
rect 11974 11704 11980 11756
rect 12032 11704 12038 11756
rect 13722 11704 13728 11756
rect 13780 11744 13786 11756
rect 14001 11747 14059 11753
rect 14001 11744 14013 11747
rect 13780 11716 14013 11744
rect 13780 11704 13786 11716
rect 14001 11713 14013 11716
rect 14047 11744 14059 11747
rect 16684 11744 16712 11840
rect 17696 11812 17724 11843
rect 17770 11840 17776 11852
rect 17828 11840 17834 11892
rect 20162 11840 20168 11892
rect 20220 11840 20226 11892
rect 17052 11784 17724 11812
rect 17052 11753 17080 11784
rect 14047 11716 16712 11744
rect 17037 11747 17095 11753
rect 14047 11713 14059 11716
rect 14001 11707 14059 11713
rect 17037 11713 17049 11747
rect 17083 11713 17095 11747
rect 17037 11707 17095 11713
rect 17126 11704 17132 11756
rect 17184 11704 17190 11756
rect 12342 11676 12348 11688
rect 11716 11648 12348 11676
rect 12342 11636 12348 11648
rect 12400 11636 12406 11688
rect 13538 11636 13544 11688
rect 13596 11676 13602 11688
rect 20180 11676 20208 11840
rect 27157 11747 27215 11753
rect 27157 11744 27169 11747
rect 13596 11648 20208 11676
rect 26712 11716 27169 11744
rect 13596 11636 13602 11648
rect 9640 11580 10824 11608
rect 11440 11608 11468 11636
rect 11882 11608 11888 11620
rect 11440 11580 11888 11608
rect 9640 11568 9646 11580
rect 11882 11568 11888 11580
rect 11940 11568 11946 11620
rect 26712 11552 26740 11716
rect 27157 11713 27169 11716
rect 27203 11713 27215 11747
rect 27157 11707 27215 11713
rect 28350 11636 28356 11688
rect 28408 11636 28414 11688
rect 9030 11540 9036 11552
rect 8956 11512 9036 11540
rect 9030 11500 9036 11512
rect 9088 11500 9094 11552
rect 9401 11543 9459 11549
rect 9401 11509 9413 11543
rect 9447 11540 9459 11543
rect 9490 11540 9496 11552
rect 9447 11512 9496 11540
rect 9447 11509 9459 11512
rect 9401 11503 9459 11509
rect 9490 11500 9496 11512
rect 9548 11500 9554 11552
rect 11333 11543 11391 11549
rect 11333 11509 11345 11543
rect 11379 11540 11391 11543
rect 11698 11540 11704 11552
rect 11379 11512 11704 11540
rect 11379 11509 11391 11512
rect 11333 11503 11391 11509
rect 11698 11500 11704 11512
rect 11756 11500 11762 11552
rect 11793 11543 11851 11549
rect 11793 11509 11805 11543
rect 11839 11540 11851 11543
rect 12250 11540 12256 11552
rect 11839 11512 12256 11540
rect 11839 11509 11851 11512
rect 11793 11503 11851 11509
rect 12250 11500 12256 11512
rect 12308 11500 12314 11552
rect 17313 11543 17371 11549
rect 17313 11509 17325 11543
rect 17359 11540 17371 11543
rect 19242 11540 19248 11552
rect 17359 11512 19248 11540
rect 17359 11509 17371 11512
rect 17313 11503 17371 11509
rect 19242 11500 19248 11512
rect 19300 11500 19306 11552
rect 26694 11500 26700 11552
rect 26752 11500 26758 11552
rect 1104 11450 28888 11472
rect 1104 11398 4423 11450
rect 4475 11398 4487 11450
rect 4539 11398 4551 11450
rect 4603 11398 4615 11450
rect 4667 11398 4679 11450
rect 4731 11398 11369 11450
rect 11421 11398 11433 11450
rect 11485 11398 11497 11450
rect 11549 11398 11561 11450
rect 11613 11398 11625 11450
rect 11677 11398 18315 11450
rect 18367 11398 18379 11450
rect 18431 11398 18443 11450
rect 18495 11398 18507 11450
rect 18559 11398 18571 11450
rect 18623 11398 25261 11450
rect 25313 11398 25325 11450
rect 25377 11398 25389 11450
rect 25441 11398 25453 11450
rect 25505 11398 25517 11450
rect 25569 11398 28888 11450
rect 1104 11376 28888 11398
rect 1854 11296 1860 11348
rect 1912 11336 1918 11348
rect 11425 11339 11483 11345
rect 1912 11308 10916 11336
rect 1912 11296 1918 11308
rect 1581 11271 1639 11277
rect 1581 11237 1593 11271
rect 1627 11268 1639 11271
rect 5718 11268 5724 11280
rect 1627 11240 5724 11268
rect 1627 11237 1639 11240
rect 1581 11231 1639 11237
rect 5718 11228 5724 11240
rect 5776 11228 5782 11280
rect 7374 11228 7380 11280
rect 7432 11268 7438 11280
rect 7432 11240 10180 11268
rect 7432 11228 7438 11240
rect 3326 11160 3332 11212
rect 3384 11200 3390 11212
rect 4893 11203 4951 11209
rect 4893 11200 4905 11203
rect 3384 11172 4905 11200
rect 3384 11160 3390 11172
rect 4893 11169 4905 11172
rect 4939 11169 4951 11203
rect 4893 11163 4951 11169
rect 5261 11203 5319 11209
rect 5261 11169 5273 11203
rect 5307 11200 5319 11203
rect 5307 11172 7604 11200
rect 5307 11169 5319 11172
rect 5261 11163 5319 11169
rect 1394 11092 1400 11144
rect 1452 11092 1458 11144
rect 1670 11092 1676 11144
rect 1728 11092 1734 11144
rect 5077 11135 5135 11141
rect 5077 11101 5089 11135
rect 5123 11101 5135 11135
rect 5077 11095 5135 11101
rect 4890 11024 4896 11076
rect 4948 11064 4954 11076
rect 5092 11064 5120 11095
rect 5902 11092 5908 11144
rect 5960 11092 5966 11144
rect 5994 11092 6000 11144
rect 6052 11132 6058 11144
rect 6089 11135 6147 11141
rect 6089 11132 6101 11135
rect 6052 11104 6101 11132
rect 6052 11092 6058 11104
rect 6089 11101 6101 11104
rect 6135 11101 6147 11135
rect 6089 11095 6147 11101
rect 7466 11092 7472 11144
rect 7524 11092 7530 11144
rect 7576 11132 7604 11172
rect 7650 11160 7656 11212
rect 7708 11200 7714 11212
rect 8205 11203 8263 11209
rect 8205 11200 8217 11203
rect 7708 11172 8217 11200
rect 7708 11160 7714 11172
rect 8205 11169 8217 11172
rect 8251 11169 8263 11203
rect 8205 11163 8263 11169
rect 8573 11203 8631 11209
rect 8573 11169 8585 11203
rect 8619 11200 8631 11203
rect 8846 11200 8852 11212
rect 8619 11172 8852 11200
rect 8619 11169 8631 11172
rect 8573 11163 8631 11169
rect 8846 11160 8852 11172
rect 8904 11160 8910 11212
rect 8938 11160 8944 11212
rect 8996 11160 9002 11212
rect 9306 11160 9312 11212
rect 9364 11160 9370 11212
rect 9677 11203 9735 11209
rect 9677 11169 9689 11203
rect 9723 11200 9735 11203
rect 10042 11200 10048 11212
rect 9723 11172 10048 11200
rect 9723 11169 9735 11172
rect 9677 11163 9735 11169
rect 10042 11160 10048 11172
rect 10100 11160 10106 11212
rect 7576 11104 8240 11132
rect 6365 11067 6423 11073
rect 4948 11036 5120 11064
rect 5276 11036 6316 11064
rect 4948 11024 4954 11036
rect 1857 10999 1915 11005
rect 1857 10965 1869 10999
rect 1903 10996 1915 10999
rect 5276 10996 5304 11036
rect 1903 10968 5304 10996
rect 1903 10965 1915 10968
rect 1857 10959 1915 10965
rect 5350 10956 5356 11008
rect 5408 10956 5414 11008
rect 6288 10996 6316 11036
rect 6365 11033 6377 11067
rect 6411 11064 6423 11067
rect 6638 11064 6644 11076
rect 6411 11036 6644 11064
rect 6411 11033 6423 11036
rect 6365 11027 6423 11033
rect 6638 11024 6644 11036
rect 6696 11024 6702 11076
rect 8018 11024 8024 11076
rect 8076 11064 8082 11076
rect 8113 11067 8171 11073
rect 8113 11064 8125 11067
rect 8076 11036 8125 11064
rect 8076 11024 8082 11036
rect 8113 11033 8125 11036
rect 8159 11033 8171 11067
rect 8212 11064 8240 11104
rect 8386 11092 8392 11144
rect 8444 11092 8450 11144
rect 9125 11135 9183 11141
rect 9125 11101 9137 11135
rect 9171 11132 9183 11135
rect 9582 11132 9588 11144
rect 9171 11104 9588 11132
rect 9171 11101 9183 11104
rect 9125 11095 9183 11101
rect 9582 11092 9588 11104
rect 9640 11092 9646 11144
rect 9861 11135 9919 11141
rect 9861 11101 9873 11135
rect 9907 11132 9919 11135
rect 10152 11132 10180 11240
rect 10781 11203 10839 11209
rect 10781 11169 10793 11203
rect 10827 11169 10839 11203
rect 10888 11200 10916 11308
rect 11425 11305 11437 11339
rect 11471 11336 11483 11339
rect 12434 11336 12440 11348
rect 11471 11308 12440 11336
rect 11471 11305 11483 11308
rect 11425 11299 11483 11305
rect 12434 11296 12440 11308
rect 12492 11296 12498 11348
rect 16574 11200 16580 11212
rect 10888 11172 14320 11200
rect 10781 11163 10839 11169
rect 9907 11104 10180 11132
rect 10796 11132 10824 11163
rect 11238 11132 11244 11144
rect 10796 11104 11244 11132
rect 9907 11101 9919 11104
rect 9861 11095 9919 11101
rect 11238 11092 11244 11104
rect 11296 11092 11302 11144
rect 11514 11092 11520 11144
rect 11572 11092 11578 11144
rect 13078 11092 13084 11144
rect 13136 11132 13142 11144
rect 14292 11141 14320 11172
rect 14384 11172 16580 11200
rect 13541 11135 13599 11141
rect 13541 11132 13553 11135
rect 13136 11104 13553 11132
rect 13136 11092 13142 11104
rect 13541 11101 13553 11104
rect 13587 11132 13599 11135
rect 14185 11135 14243 11141
rect 14185 11132 14197 11135
rect 13587 11104 14197 11132
rect 13587 11101 13599 11104
rect 13541 11095 13599 11101
rect 14185 11101 14197 11104
rect 14231 11101 14243 11135
rect 14185 11095 14243 11101
rect 14277 11135 14335 11141
rect 14277 11101 14289 11135
rect 14323 11101 14335 11135
rect 14277 11095 14335 11101
rect 10965 11067 11023 11073
rect 10965 11064 10977 11067
rect 8212 11036 10977 11064
rect 8113 11027 8171 11033
rect 10965 11033 10977 11036
rect 11011 11033 11023 11067
rect 10965 11027 11023 11033
rect 11057 11067 11115 11073
rect 11057 11033 11069 11067
rect 11103 11064 11115 11067
rect 11793 11067 11851 11073
rect 11103 11036 11560 11064
rect 11103 11033 11115 11036
rect 11057 11027 11115 11033
rect 7374 10996 7380 11008
rect 6288 10968 7380 10996
rect 7374 10956 7380 10968
rect 7432 10956 7438 11008
rect 8128 10996 8156 11027
rect 9766 10996 9772 11008
rect 8128 10968 9772 10996
rect 9766 10956 9772 10968
rect 9824 10956 9830 11008
rect 10045 10999 10103 11005
rect 10045 10965 10057 10999
rect 10091 10996 10103 10999
rect 10226 10996 10232 11008
rect 10091 10968 10232 10996
rect 10091 10965 10103 10968
rect 10045 10959 10103 10965
rect 10226 10956 10232 10968
rect 10284 10956 10290 11008
rect 11532 10996 11560 11036
rect 11793 11033 11805 11067
rect 11839 11064 11851 11067
rect 11882 11064 11888 11076
rect 11839 11036 11888 11064
rect 11839 11033 11851 11036
rect 11793 11027 11851 11033
rect 11882 11024 11888 11036
rect 11940 11024 11946 11076
rect 12250 11024 12256 11076
rect 12308 11024 12314 11076
rect 14200 11064 14228 11095
rect 14384 11064 14412 11172
rect 16574 11160 16580 11172
rect 16632 11160 16638 11212
rect 14200 11036 14412 11064
rect 14458 11024 14464 11076
rect 14516 11024 14522 11076
rect 13538 10996 13544 11008
rect 11532 10968 13544 10996
rect 13538 10956 13544 10968
rect 13596 10956 13602 11008
rect 1104 10906 29048 10928
rect 1104 10854 7896 10906
rect 7948 10854 7960 10906
rect 8012 10854 8024 10906
rect 8076 10854 8088 10906
rect 8140 10854 8152 10906
rect 8204 10854 14842 10906
rect 14894 10854 14906 10906
rect 14958 10854 14970 10906
rect 15022 10854 15034 10906
rect 15086 10854 15098 10906
rect 15150 10854 21788 10906
rect 21840 10854 21852 10906
rect 21904 10854 21916 10906
rect 21968 10854 21980 10906
rect 22032 10854 22044 10906
rect 22096 10854 28734 10906
rect 28786 10854 28798 10906
rect 28850 10854 28862 10906
rect 28914 10854 28926 10906
rect 28978 10854 28990 10906
rect 29042 10854 29048 10906
rect 1104 10832 29048 10854
rect 5445 10795 5503 10801
rect 5445 10761 5457 10795
rect 5491 10792 5503 10795
rect 5902 10792 5908 10804
rect 5491 10764 5908 10792
rect 5491 10761 5503 10764
rect 5445 10755 5503 10761
rect 5902 10752 5908 10764
rect 5960 10752 5966 10804
rect 6178 10752 6184 10804
rect 6236 10792 6242 10804
rect 7006 10792 7012 10804
rect 6236 10764 7012 10792
rect 6236 10752 6242 10764
rect 7006 10752 7012 10764
rect 7064 10752 7070 10804
rect 7466 10752 7472 10804
rect 7524 10792 7530 10804
rect 7561 10795 7619 10801
rect 7561 10792 7573 10795
rect 7524 10764 7573 10792
rect 7524 10752 7530 10764
rect 7561 10761 7573 10764
rect 7607 10761 7619 10795
rect 7561 10755 7619 10761
rect 10502 10752 10508 10804
rect 10560 10752 10566 10804
rect 26694 10792 26700 10804
rect 10612 10764 13860 10792
rect 4893 10727 4951 10733
rect 4893 10693 4905 10727
rect 4939 10724 4951 10727
rect 5074 10724 5080 10736
rect 4939 10696 5080 10724
rect 4939 10693 4951 10696
rect 4893 10687 4951 10693
rect 5074 10684 5080 10696
rect 5132 10724 5138 10736
rect 5132 10696 5396 10724
rect 5132 10684 5138 10696
rect 934 10616 940 10668
rect 992 10656 998 10668
rect 1397 10659 1455 10665
rect 1397 10656 1409 10659
rect 992 10628 1409 10656
rect 992 10616 998 10628
rect 1397 10625 1409 10628
rect 1443 10625 1455 10659
rect 1397 10619 1455 10625
rect 1673 10659 1731 10665
rect 1673 10625 1685 10659
rect 1719 10625 1731 10659
rect 1673 10619 1731 10625
rect 1026 10548 1032 10600
rect 1084 10588 1090 10600
rect 1688 10588 1716 10619
rect 4154 10616 4160 10668
rect 4212 10656 4218 10668
rect 4985 10659 5043 10665
rect 4985 10656 4997 10659
rect 4212 10628 4997 10656
rect 4212 10616 4218 10628
rect 4985 10625 4997 10628
rect 5031 10625 5043 10659
rect 4985 10619 5043 10625
rect 5169 10659 5227 10665
rect 5169 10625 5181 10659
rect 5215 10625 5227 10659
rect 5368 10656 5396 10696
rect 5718 10684 5724 10736
rect 5776 10724 5782 10736
rect 5776 10696 7972 10724
rect 5776 10684 5782 10696
rect 5813 10659 5871 10665
rect 5813 10656 5825 10659
rect 5368 10628 5825 10656
rect 5169 10619 5227 10625
rect 5813 10625 5825 10628
rect 5859 10656 5871 10659
rect 5859 10628 6316 10656
rect 5859 10625 5871 10628
rect 5813 10619 5871 10625
rect 1084 10560 1716 10588
rect 1084 10548 1090 10560
rect 4338 10548 4344 10600
rect 4396 10588 4402 10600
rect 5184 10588 5212 10619
rect 4396 10560 5212 10588
rect 5353 10591 5411 10597
rect 4396 10548 4402 10560
rect 5353 10557 5365 10591
rect 5399 10588 5411 10591
rect 5905 10591 5963 10597
rect 5905 10588 5917 10591
rect 5399 10560 5917 10588
rect 5399 10557 5411 10560
rect 5353 10551 5411 10557
rect 5905 10557 5917 10560
rect 5951 10557 5963 10591
rect 5905 10551 5963 10557
rect 6089 10591 6147 10597
rect 6089 10557 6101 10591
rect 6135 10588 6147 10591
rect 6178 10588 6184 10600
rect 6135 10560 6184 10588
rect 6135 10557 6147 10560
rect 6089 10551 6147 10557
rect 6178 10548 6184 10560
rect 6236 10548 6242 10600
rect 6288 10588 6316 10628
rect 6546 10616 6552 10668
rect 6604 10616 6610 10668
rect 6638 10616 6644 10668
rect 6696 10616 6702 10668
rect 6822 10616 6828 10668
rect 6880 10656 6886 10668
rect 7193 10659 7251 10665
rect 7193 10656 7205 10659
rect 6880 10628 7205 10656
rect 6880 10616 6886 10628
rect 7193 10625 7205 10628
rect 7239 10656 7251 10659
rect 7653 10659 7711 10665
rect 7653 10656 7665 10659
rect 7239 10628 7665 10656
rect 7239 10625 7251 10628
rect 7193 10619 7251 10625
rect 7653 10625 7665 10628
rect 7699 10625 7711 10659
rect 7653 10619 7711 10625
rect 6656 10588 6684 10616
rect 6288 10560 6684 10588
rect 7668 10588 7696 10619
rect 7742 10616 7748 10668
rect 7800 10656 7806 10668
rect 7837 10659 7895 10665
rect 7837 10656 7849 10659
rect 7800 10628 7849 10656
rect 7800 10616 7806 10628
rect 7837 10625 7849 10628
rect 7883 10625 7895 10659
rect 7944 10656 7972 10696
rect 9674 10684 9680 10736
rect 9732 10724 9738 10736
rect 10410 10724 10416 10736
rect 9732 10696 10416 10724
rect 9732 10684 9738 10696
rect 10410 10684 10416 10696
rect 10468 10684 10474 10736
rect 10612 10656 10640 10764
rect 12802 10684 12808 10736
rect 12860 10684 12866 10736
rect 13538 10684 13544 10736
rect 13596 10684 13602 10736
rect 7944 10628 10640 10656
rect 7837 10619 7895 10625
rect 13722 10616 13728 10668
rect 13780 10616 13786 10668
rect 13832 10665 13860 10764
rect 13924 10764 26700 10792
rect 13817 10659 13875 10665
rect 13817 10625 13829 10659
rect 13863 10625 13875 10659
rect 13817 10619 13875 10625
rect 8294 10588 8300 10600
rect 7668 10560 8300 10588
rect 8294 10548 8300 10560
rect 8352 10548 8358 10600
rect 9585 10591 9643 10597
rect 9585 10557 9597 10591
rect 9631 10557 9643 10591
rect 9585 10551 9643 10557
rect 1578 10480 1584 10532
rect 1636 10480 1642 10532
rect 6454 10520 6460 10532
rect 1872 10492 6460 10520
rect 1872 10461 1900 10492
rect 6454 10480 6460 10492
rect 6512 10480 6518 10532
rect 6546 10480 6552 10532
rect 6604 10480 6610 10532
rect 9600 10520 9628 10551
rect 10318 10548 10324 10600
rect 10376 10548 10382 10600
rect 10870 10548 10876 10600
rect 10928 10588 10934 10600
rect 11057 10591 11115 10597
rect 11057 10588 11069 10591
rect 10928 10560 11069 10588
rect 10928 10548 10934 10560
rect 11057 10557 11069 10560
rect 11103 10557 11115 10591
rect 11057 10551 11115 10557
rect 11514 10548 11520 10600
rect 11572 10548 11578 10600
rect 11790 10548 11796 10600
rect 11848 10548 11854 10600
rect 9950 10520 9956 10532
rect 9600 10492 9956 10520
rect 9950 10480 9956 10492
rect 10008 10520 10014 10532
rect 11532 10520 11560 10548
rect 10008 10492 11560 10520
rect 10008 10480 10014 10492
rect 1857 10455 1915 10461
rect 1857 10421 1869 10455
rect 1903 10421 1915 10455
rect 1857 10415 1915 10421
rect 4154 10412 4160 10464
rect 4212 10452 4218 10464
rect 4525 10455 4583 10461
rect 4525 10452 4537 10455
rect 4212 10424 4537 10452
rect 4212 10412 4218 10424
rect 4525 10421 4537 10424
rect 4571 10452 4583 10455
rect 6564 10452 6592 10480
rect 4571 10424 6592 10452
rect 9769 10455 9827 10461
rect 4571 10421 4583 10424
rect 4525 10415 4583 10421
rect 9769 10421 9781 10455
rect 9815 10452 9827 10455
rect 10042 10452 10048 10464
rect 9815 10424 10048 10452
rect 9815 10421 9827 10424
rect 9769 10415 9827 10421
rect 10042 10412 10048 10424
rect 10100 10412 10106 10464
rect 10134 10412 10140 10464
rect 10192 10452 10198 10464
rect 13924 10452 13952 10764
rect 26694 10752 26700 10764
rect 26752 10752 26758 10804
rect 15657 10727 15715 10733
rect 15657 10693 15669 10727
rect 15703 10724 15715 10727
rect 16022 10724 16028 10736
rect 15703 10696 16028 10724
rect 15703 10693 15715 10696
rect 15657 10687 15715 10693
rect 15764 10665 15792 10696
rect 16022 10684 16028 10696
rect 16080 10684 16086 10736
rect 15749 10659 15807 10665
rect 15749 10625 15761 10659
rect 15795 10656 15807 10659
rect 15795 10628 15829 10656
rect 15795 10625 15807 10628
rect 15749 10619 15807 10625
rect 15930 10616 15936 10668
rect 15988 10616 15994 10668
rect 17126 10616 17132 10668
rect 17184 10656 17190 10668
rect 27157 10659 27215 10665
rect 27157 10656 27169 10659
rect 17184 10628 27169 10656
rect 17184 10616 17190 10628
rect 27157 10625 27169 10628
rect 27203 10625 27215 10659
rect 27157 10619 27215 10625
rect 28350 10548 28356 10600
rect 28408 10548 28414 10600
rect 10192 10424 13952 10452
rect 10192 10412 10198 10424
rect 13998 10412 14004 10464
rect 14056 10412 14062 10464
rect 16114 10412 16120 10464
rect 16172 10412 16178 10464
rect 1104 10362 28888 10384
rect 1104 10310 4423 10362
rect 4475 10310 4487 10362
rect 4539 10310 4551 10362
rect 4603 10310 4615 10362
rect 4667 10310 4679 10362
rect 4731 10310 11369 10362
rect 11421 10310 11433 10362
rect 11485 10310 11497 10362
rect 11549 10310 11561 10362
rect 11613 10310 11625 10362
rect 11677 10310 18315 10362
rect 18367 10310 18379 10362
rect 18431 10310 18443 10362
rect 18495 10310 18507 10362
rect 18559 10310 18571 10362
rect 18623 10310 25261 10362
rect 25313 10310 25325 10362
rect 25377 10310 25389 10362
rect 25441 10310 25453 10362
rect 25505 10310 25517 10362
rect 25569 10310 28888 10362
rect 1104 10288 28888 10310
rect 290 10208 296 10260
rect 348 10248 354 10260
rect 658 10248 664 10260
rect 348 10220 664 10248
rect 348 10208 354 10220
rect 658 10208 664 10220
rect 716 10208 722 10260
rect 4908 10220 6316 10248
rect 1857 10183 1915 10189
rect 1857 10149 1869 10183
rect 1903 10149 1915 10183
rect 1857 10143 1915 10149
rect 1872 10112 1900 10143
rect 4908 10112 4936 10220
rect 6288 10180 6316 10220
rect 6454 10208 6460 10260
rect 6512 10248 6518 10260
rect 7374 10248 7380 10260
rect 6512 10220 7380 10248
rect 6512 10208 6518 10220
rect 7374 10208 7380 10220
rect 7432 10208 7438 10260
rect 8478 10208 8484 10260
rect 8536 10248 8542 10260
rect 8665 10251 8723 10257
rect 8665 10248 8677 10251
rect 8536 10220 8677 10248
rect 8536 10208 8542 10220
rect 8665 10217 8677 10220
rect 8711 10217 8723 10251
rect 8665 10211 8723 10217
rect 9858 10208 9864 10260
rect 9916 10208 9922 10260
rect 10042 10208 10048 10260
rect 10100 10208 10106 10260
rect 11790 10208 11796 10260
rect 11848 10248 11854 10260
rect 11885 10251 11943 10257
rect 11885 10248 11897 10251
rect 11848 10220 11897 10248
rect 11848 10208 11854 10220
rect 11885 10217 11897 10220
rect 11931 10217 11943 10251
rect 11885 10211 11943 10217
rect 12713 10251 12771 10257
rect 12713 10217 12725 10251
rect 12759 10248 12771 10251
rect 12802 10248 12808 10260
rect 12759 10220 12808 10248
rect 12759 10217 12771 10220
rect 12713 10211 12771 10217
rect 12802 10208 12808 10220
rect 12860 10208 12866 10260
rect 17126 10208 17132 10260
rect 17184 10208 17190 10260
rect 17218 10208 17224 10260
rect 17276 10248 17282 10260
rect 26973 10251 27031 10257
rect 26973 10248 26985 10251
rect 17276 10220 26985 10248
rect 17276 10208 17282 10220
rect 26973 10217 26985 10220
rect 27019 10217 27031 10251
rect 26973 10211 27031 10217
rect 9674 10180 9680 10192
rect 6288 10152 9680 10180
rect 9674 10140 9680 10152
rect 9732 10140 9738 10192
rect 1872 10084 4936 10112
rect 4985 10115 5043 10121
rect 4985 10081 4997 10115
rect 5031 10112 5043 10115
rect 5994 10112 6000 10124
rect 5031 10084 6000 10112
rect 5031 10081 5043 10084
rect 4985 10075 5043 10081
rect 5994 10072 6000 10084
rect 6052 10072 6058 10124
rect 7006 10072 7012 10124
rect 7064 10112 7070 10124
rect 7285 10115 7343 10121
rect 7285 10112 7297 10115
rect 7064 10084 7297 10112
rect 7064 10072 7070 10084
rect 7285 10081 7297 10084
rect 7331 10081 7343 10115
rect 7285 10075 7343 10081
rect 9950 10072 9956 10124
rect 10008 10072 10014 10124
rect 10060 10112 10088 10208
rect 11701 10183 11759 10189
rect 11701 10149 11713 10183
rect 11747 10180 11759 10183
rect 12066 10180 12072 10192
rect 11747 10152 12072 10180
rect 11747 10149 11759 10152
rect 11701 10143 11759 10149
rect 12066 10140 12072 10152
rect 12124 10180 12130 10192
rect 17144 10180 17172 10208
rect 12124 10152 17172 10180
rect 12124 10140 12130 10152
rect 10229 10115 10287 10121
rect 10229 10112 10241 10115
rect 10060 10084 10241 10112
rect 10229 10081 10241 10084
rect 10275 10081 10287 10115
rect 10229 10075 10287 10081
rect 12434 10072 12440 10124
rect 12492 10072 12498 10124
rect 934 10004 940 10056
rect 992 10044 998 10056
rect 1397 10047 1455 10053
rect 1397 10044 1409 10047
rect 992 10016 1409 10044
rect 992 10004 998 10016
rect 1397 10013 1409 10016
rect 1443 10013 1455 10047
rect 1397 10007 1455 10013
rect 1670 10004 1676 10056
rect 1728 10004 1734 10056
rect 6638 10004 6644 10056
rect 6696 10044 6702 10056
rect 8113 10047 8171 10053
rect 6696 10016 7052 10044
rect 6696 10004 6702 10016
rect 5261 9979 5319 9985
rect 1596 9948 5212 9976
rect 1596 9917 1624 9948
rect 1581 9911 1639 9917
rect 1581 9877 1593 9911
rect 1627 9877 1639 9911
rect 1581 9871 1639 9877
rect 2225 9911 2283 9917
rect 2225 9877 2237 9911
rect 2271 9908 2283 9911
rect 3142 9908 3148 9920
rect 2271 9880 3148 9908
rect 2271 9877 2283 9880
rect 2225 9871 2283 9877
rect 3142 9868 3148 9880
rect 3200 9868 3206 9920
rect 4798 9868 4804 9920
rect 4856 9868 4862 9920
rect 5184 9908 5212 9948
rect 5261 9945 5273 9979
rect 5307 9976 5319 9979
rect 5350 9976 5356 9988
rect 5307 9948 5356 9976
rect 5307 9945 5319 9948
rect 5261 9939 5319 9945
rect 5350 9936 5356 9948
rect 5408 9936 5414 9988
rect 5718 9936 5724 9988
rect 5776 9936 5782 9988
rect 7024 9985 7052 10016
rect 8113 10013 8125 10047
rect 8159 10044 8171 10047
rect 8662 10044 8668 10056
rect 8159 10016 8668 10044
rect 8159 10013 8171 10016
rect 8113 10007 8171 10013
rect 8662 10004 8668 10016
rect 8720 10044 8726 10056
rect 9214 10044 9220 10056
rect 8720 10016 9220 10044
rect 8720 10004 8726 10016
rect 9214 10004 9220 10016
rect 9272 10004 9278 10056
rect 9309 10047 9367 10053
rect 9309 10013 9321 10047
rect 9355 10044 9367 10047
rect 9858 10044 9864 10056
rect 9355 10016 9864 10044
rect 9355 10013 9367 10016
rect 9309 10007 9367 10013
rect 9858 10004 9864 10016
rect 9916 10004 9922 10056
rect 12342 10004 12348 10056
rect 12400 10044 12406 10056
rect 12805 10047 12863 10053
rect 12805 10044 12817 10047
rect 12400 10016 12817 10044
rect 12400 10004 12406 10016
rect 12805 10013 12817 10016
rect 12851 10013 12863 10047
rect 26988 10044 27016 10211
rect 27157 10047 27215 10053
rect 27157 10044 27169 10047
rect 26988 10016 27169 10044
rect 12805 10007 12863 10013
rect 27157 10013 27169 10016
rect 27203 10013 27215 10047
rect 27157 10007 27215 10013
rect 7009 9979 7067 9985
rect 7009 9945 7021 9979
rect 7055 9976 7067 9979
rect 10134 9976 10140 9988
rect 7055 9948 10140 9976
rect 7055 9945 7067 9948
rect 7009 9939 7067 9945
rect 10134 9936 10140 9948
rect 10192 9936 10198 9988
rect 11514 9976 11520 9988
rect 11454 9948 11520 9976
rect 11514 9936 11520 9948
rect 11572 9936 11578 9988
rect 28350 9936 28356 9988
rect 28408 9936 28414 9988
rect 11054 9908 11060 9920
rect 5184 9880 11060 9908
rect 11054 9868 11060 9880
rect 11112 9868 11118 9920
rect 1104 9818 29048 9840
rect 1104 9766 7896 9818
rect 7948 9766 7960 9818
rect 8012 9766 8024 9818
rect 8076 9766 8088 9818
rect 8140 9766 8152 9818
rect 8204 9766 14842 9818
rect 14894 9766 14906 9818
rect 14958 9766 14970 9818
rect 15022 9766 15034 9818
rect 15086 9766 15098 9818
rect 15150 9766 21788 9818
rect 21840 9766 21852 9818
rect 21904 9766 21916 9818
rect 21968 9766 21980 9818
rect 22032 9766 22044 9818
rect 22096 9766 28734 9818
rect 28786 9766 28798 9818
rect 28850 9766 28862 9818
rect 28914 9766 28926 9818
rect 28978 9766 28990 9818
rect 29042 9766 29048 9818
rect 1104 9744 29048 9766
rect 1857 9707 1915 9713
rect 1857 9673 1869 9707
rect 1903 9704 1915 9707
rect 5902 9704 5908 9716
rect 1903 9676 5908 9704
rect 1903 9673 1915 9676
rect 1857 9667 1915 9673
rect 5902 9664 5908 9676
rect 5960 9664 5966 9716
rect 6822 9664 6828 9716
rect 6880 9704 6886 9716
rect 6880 9676 6960 9704
rect 6880 9664 6886 9676
rect 4614 9596 4620 9648
rect 4672 9596 4678 9648
rect 4706 9596 4712 9648
rect 4764 9636 4770 9648
rect 4801 9639 4859 9645
rect 4801 9636 4813 9639
rect 4764 9608 4813 9636
rect 4764 9596 4770 9608
rect 4801 9605 4813 9608
rect 4847 9605 4859 9639
rect 6932 9636 6960 9676
rect 7834 9664 7840 9716
rect 7892 9704 7898 9716
rect 17218 9704 17224 9716
rect 7892 9676 17224 9704
rect 7892 9664 7898 9676
rect 17218 9664 17224 9676
rect 17276 9664 17282 9716
rect 4801 9599 4859 9605
rect 5000 9608 6960 9636
rect 7009 9639 7067 9645
rect 934 9528 940 9580
rect 992 9568 998 9580
rect 1397 9571 1455 9577
rect 1397 9568 1409 9571
rect 992 9540 1409 9568
rect 992 9528 998 9540
rect 1397 9537 1409 9540
rect 1443 9537 1455 9571
rect 1397 9531 1455 9537
rect 1673 9571 1731 9577
rect 1673 9537 1685 9571
rect 1719 9537 1731 9571
rect 1673 9531 1731 9537
rect 1026 9460 1032 9512
rect 1084 9500 1090 9512
rect 1688 9500 1716 9531
rect 1762 9528 1768 9580
rect 1820 9568 1826 9580
rect 1949 9571 2007 9577
rect 1949 9568 1961 9571
rect 1820 9540 1961 9568
rect 1820 9528 1826 9540
rect 1949 9537 1961 9540
rect 1995 9537 2007 9571
rect 1949 9531 2007 9537
rect 2038 9528 2044 9580
rect 2096 9568 2102 9580
rect 2225 9571 2283 9577
rect 2225 9568 2237 9571
rect 2096 9540 2237 9568
rect 2096 9528 2102 9540
rect 2225 9537 2237 9540
rect 2271 9537 2283 9571
rect 2225 9531 2283 9537
rect 4893 9571 4951 9577
rect 4893 9537 4905 9571
rect 4939 9568 4951 9571
rect 5000 9568 5028 9608
rect 7009 9605 7021 9639
rect 7055 9636 7067 9639
rect 7190 9636 7196 9648
rect 7055 9608 7196 9636
rect 7055 9605 7067 9608
rect 7009 9599 7067 9605
rect 7190 9596 7196 9608
rect 7248 9596 7254 9648
rect 7374 9596 7380 9648
rect 7432 9636 7438 9648
rect 7432 9608 9260 9636
rect 7432 9596 7438 9608
rect 4939 9540 5028 9568
rect 4939 9537 4951 9540
rect 4893 9531 4951 9537
rect 5074 9528 5080 9580
rect 5132 9528 5138 9580
rect 5166 9528 5172 9580
rect 5224 9566 5230 9580
rect 5224 9538 5267 9566
rect 5224 9528 5230 9538
rect 6178 9528 6184 9580
rect 6236 9528 6242 9580
rect 6365 9571 6423 9577
rect 6365 9537 6377 9571
rect 6411 9568 6423 9571
rect 6454 9568 6460 9580
rect 6411 9540 6460 9568
rect 6411 9537 6423 9540
rect 6365 9531 6423 9537
rect 6454 9528 6460 9540
rect 6512 9528 6518 9580
rect 6546 9528 6552 9580
rect 6604 9568 6610 9580
rect 7101 9571 7159 9577
rect 7101 9568 7113 9571
rect 6604 9540 7113 9568
rect 6604 9528 6610 9540
rect 7101 9537 7113 9540
rect 7147 9537 7159 9571
rect 7101 9531 7159 9537
rect 8478 9528 8484 9580
rect 8536 9568 8542 9580
rect 9232 9577 9260 9608
rect 9398 9596 9404 9648
rect 9456 9636 9462 9648
rect 9585 9639 9643 9645
rect 9585 9636 9597 9639
rect 9456 9608 9597 9636
rect 9456 9596 9462 9608
rect 9585 9605 9597 9608
rect 9631 9605 9643 9639
rect 9585 9599 9643 9605
rect 10134 9596 10140 9648
rect 10192 9636 10198 9648
rect 10689 9639 10747 9645
rect 10192 9608 10272 9636
rect 10192 9596 10198 9608
rect 10244 9577 10272 9608
rect 10689 9605 10701 9639
rect 10735 9636 10747 9639
rect 12066 9636 12072 9648
rect 10735 9608 12072 9636
rect 10735 9605 10747 9608
rect 10689 9599 10747 9605
rect 12066 9596 12072 9608
rect 12124 9596 12130 9648
rect 9033 9571 9091 9577
rect 9033 9568 9045 9571
rect 8536 9540 9045 9568
rect 8536 9528 8542 9540
rect 9033 9537 9045 9540
rect 9079 9537 9091 9571
rect 9033 9531 9091 9537
rect 9217 9571 9275 9577
rect 9217 9537 9229 9571
rect 9263 9537 9275 9571
rect 9217 9531 9275 9537
rect 10229 9571 10287 9577
rect 10229 9537 10241 9571
rect 10275 9537 10287 9571
rect 10229 9531 10287 9537
rect 11333 9571 11391 9577
rect 11333 9537 11345 9571
rect 11379 9568 11391 9571
rect 11379 9540 11468 9568
rect 11379 9537 11391 9540
rect 11333 9531 11391 9537
rect 1084 9472 1716 9500
rect 1084 9460 1090 9472
rect 5902 9460 5908 9512
rect 5960 9500 5966 9512
rect 9674 9500 9680 9512
rect 5960 9472 9680 9500
rect 5960 9460 5966 9472
rect 9674 9460 9680 9472
rect 9732 9460 9738 9512
rect 10502 9460 10508 9512
rect 10560 9500 10566 9512
rect 10781 9503 10839 9509
rect 10781 9500 10793 9503
rect 10560 9472 10793 9500
rect 10560 9460 10566 9472
rect 10781 9469 10793 9472
rect 10827 9469 10839 9503
rect 10781 9463 10839 9469
rect 10965 9503 11023 9509
rect 10965 9469 10977 9503
rect 11011 9469 11023 9503
rect 10965 9463 11023 9469
rect 11241 9503 11299 9509
rect 11241 9469 11253 9503
rect 11287 9500 11299 9503
rect 11440 9500 11468 9540
rect 11698 9528 11704 9580
rect 11756 9568 11762 9580
rect 12161 9571 12219 9577
rect 12161 9568 12173 9571
rect 11756 9540 12173 9568
rect 11756 9528 11762 9540
rect 12161 9537 12173 9540
rect 12207 9537 12219 9571
rect 12161 9531 12219 9537
rect 14182 9528 14188 9580
rect 14240 9528 14246 9580
rect 14001 9503 14059 9509
rect 11287 9472 11376 9500
rect 11440 9472 11836 9500
rect 11287 9469 11299 9472
rect 11241 9463 11299 9469
rect 1581 9435 1639 9441
rect 1581 9401 1593 9435
rect 1627 9432 1639 9435
rect 1627 9404 5028 9432
rect 1627 9401 1639 9404
rect 1581 9395 1639 9401
rect 2130 9324 2136 9376
rect 2188 9324 2194 9376
rect 2406 9324 2412 9376
rect 2464 9324 2470 9376
rect 2777 9367 2835 9373
rect 2777 9333 2789 9367
rect 2823 9364 2835 9367
rect 3145 9367 3203 9373
rect 3145 9364 3157 9367
rect 2823 9336 3157 9364
rect 2823 9333 2835 9336
rect 2777 9327 2835 9333
rect 3145 9333 3157 9336
rect 3191 9364 3203 9367
rect 3786 9364 3792 9376
rect 3191 9336 3792 9364
rect 3191 9333 3203 9336
rect 3145 9327 3203 9333
rect 3786 9324 3792 9336
rect 3844 9324 3850 9376
rect 4154 9324 4160 9376
rect 4212 9324 4218 9376
rect 5000 9364 5028 9404
rect 5626 9392 5632 9444
rect 5684 9432 5690 9444
rect 10042 9432 10048 9444
rect 5684 9404 10048 9432
rect 5684 9392 5690 9404
rect 10042 9392 10048 9404
rect 10100 9392 10106 9444
rect 10980 9432 11008 9463
rect 11348 9432 11376 9472
rect 11422 9432 11428 9444
rect 10980 9404 11284 9432
rect 11348 9404 11428 9432
rect 11256 9376 11284 9404
rect 11422 9392 11428 9404
rect 11480 9392 11486 9444
rect 11808 9376 11836 9472
rect 14001 9469 14013 9503
rect 14047 9469 14059 9503
rect 14001 9463 14059 9469
rect 13538 9392 13544 9444
rect 13596 9432 13602 9444
rect 14016 9432 14044 9463
rect 13596 9404 14044 9432
rect 13596 9392 13602 9404
rect 17218 9392 17224 9444
rect 17276 9432 17282 9444
rect 23842 9432 23848 9444
rect 17276 9404 23848 9432
rect 17276 9392 17282 9404
rect 23842 9392 23848 9404
rect 23900 9392 23906 9444
rect 5166 9364 5172 9376
rect 5000 9336 5172 9364
rect 5166 9324 5172 9336
rect 5224 9324 5230 9376
rect 5350 9324 5356 9376
rect 5408 9324 5414 9376
rect 5537 9367 5595 9373
rect 5537 9333 5549 9367
rect 5583 9364 5595 9367
rect 5810 9364 5816 9376
rect 5583 9336 5816 9364
rect 5583 9333 5595 9336
rect 5537 9327 5595 9333
rect 5810 9324 5816 9336
rect 5868 9324 5874 9376
rect 7098 9324 7104 9376
rect 7156 9364 7162 9376
rect 7742 9364 7748 9376
rect 7156 9336 7748 9364
rect 7156 9324 7162 9336
rect 7742 9324 7748 9336
rect 7800 9364 7806 9376
rect 8389 9367 8447 9373
rect 8389 9364 8401 9367
rect 7800 9336 8401 9364
rect 7800 9324 7806 9336
rect 8389 9333 8401 9336
rect 8435 9333 8447 9367
rect 8389 9327 8447 9333
rect 9401 9367 9459 9373
rect 9401 9333 9413 9367
rect 9447 9364 9459 9367
rect 9490 9364 9496 9376
rect 9447 9336 9496 9364
rect 9447 9333 9459 9336
rect 9401 9327 9459 9333
rect 9490 9324 9496 9336
rect 9548 9324 9554 9376
rect 10318 9324 10324 9376
rect 10376 9324 10382 9376
rect 11238 9324 11244 9376
rect 11296 9324 11302 9376
rect 11790 9324 11796 9376
rect 11848 9364 11854 9376
rect 13814 9364 13820 9376
rect 11848 9336 13820 9364
rect 11848 9324 11854 9336
rect 13814 9324 13820 9336
rect 13872 9324 13878 9376
rect 14369 9367 14427 9373
rect 14369 9333 14381 9367
rect 14415 9364 14427 9367
rect 25774 9364 25780 9376
rect 14415 9336 25780 9364
rect 14415 9333 14427 9336
rect 14369 9327 14427 9333
rect 25774 9324 25780 9336
rect 25832 9324 25838 9376
rect 1104 9274 28888 9296
rect 1104 9222 4423 9274
rect 4475 9222 4487 9274
rect 4539 9222 4551 9274
rect 4603 9222 4615 9274
rect 4667 9222 4679 9274
rect 4731 9222 11369 9274
rect 11421 9222 11433 9274
rect 11485 9222 11497 9274
rect 11549 9222 11561 9274
rect 11613 9222 11625 9274
rect 11677 9222 18315 9274
rect 18367 9222 18379 9274
rect 18431 9222 18443 9274
rect 18495 9222 18507 9274
rect 18559 9222 18571 9274
rect 18623 9222 25261 9274
rect 25313 9222 25325 9274
rect 25377 9222 25389 9274
rect 25441 9222 25453 9274
rect 25505 9222 25517 9274
rect 25569 9222 28888 9274
rect 1104 9200 28888 9222
rect 1857 9163 1915 9169
rect 1857 9129 1869 9163
rect 1903 9160 1915 9163
rect 1903 9132 5580 9160
rect 1903 9129 1915 9132
rect 1857 9123 1915 9129
rect 1578 9052 1584 9104
rect 1636 9052 1642 9104
rect 4709 9095 4767 9101
rect 4709 9061 4721 9095
rect 4755 9092 4767 9095
rect 5442 9092 5448 9104
rect 4755 9064 5448 9092
rect 4755 9061 4767 9064
rect 4709 9055 4767 9061
rect 5442 9052 5448 9064
rect 5500 9052 5506 9104
rect 5552 9092 5580 9132
rect 5626 9120 5632 9172
rect 5684 9120 5690 9172
rect 5810 9120 5816 9172
rect 5868 9120 5874 9172
rect 6454 9120 6460 9172
rect 6512 9160 6518 9172
rect 7466 9160 7472 9172
rect 6512 9132 7472 9160
rect 6512 9120 6518 9132
rect 7466 9120 7472 9132
rect 7524 9120 7530 9172
rect 7558 9120 7564 9172
rect 7616 9160 7622 9172
rect 8113 9163 8171 9169
rect 8113 9160 8125 9163
rect 7616 9132 8125 9160
rect 7616 9120 7622 9132
rect 8113 9129 8125 9132
rect 8159 9129 8171 9163
rect 9858 9160 9864 9172
rect 8113 9123 8171 9129
rect 9048 9132 9864 9160
rect 5552 9064 5764 9092
rect 1302 8984 1308 9036
rect 1360 9024 1366 9036
rect 1360 8996 2636 9024
rect 1360 8984 1366 8996
rect 934 8916 940 8968
rect 992 8956 998 8968
rect 1397 8959 1455 8965
rect 1397 8956 1409 8959
rect 992 8928 1409 8956
rect 992 8916 998 8928
rect 1397 8925 1409 8928
rect 1443 8925 1455 8959
rect 1397 8919 1455 8925
rect 1673 8959 1731 8965
rect 1673 8925 1685 8959
rect 1719 8925 1731 8959
rect 1673 8919 1731 8925
rect 1026 8848 1032 8900
rect 1084 8888 1090 8900
rect 1688 8888 1716 8919
rect 1854 8916 1860 8968
rect 1912 8956 1918 8968
rect 2133 8959 2191 8965
rect 2133 8956 2145 8959
rect 1912 8928 2145 8956
rect 1912 8916 1918 8928
rect 2133 8925 2145 8928
rect 2179 8925 2191 8959
rect 2133 8919 2191 8925
rect 2222 8916 2228 8968
rect 2280 8916 2286 8968
rect 2498 8956 2504 8968
rect 2424 8928 2504 8956
rect 2314 8888 2320 8900
rect 1084 8860 1716 8888
rect 1780 8860 2320 8888
rect 1084 8848 1090 8860
rect 842 8780 848 8832
rect 900 8820 906 8832
rect 1780 8820 1808 8860
rect 2314 8848 2320 8860
rect 2372 8848 2378 8900
rect 900 8792 1808 8820
rect 900 8780 906 8792
rect 1946 8780 1952 8832
rect 2004 8780 2010 8832
rect 2424 8829 2452 8928
rect 2498 8916 2504 8928
rect 2556 8916 2562 8968
rect 2608 8888 2636 8996
rect 2700 8996 3464 9024
rect 2700 8965 2728 8996
rect 2685 8959 2743 8965
rect 2685 8925 2697 8959
rect 2731 8925 2743 8959
rect 3436 8956 3464 8996
rect 3510 8984 3516 9036
rect 3568 9024 3574 9036
rect 4801 9027 4859 9033
rect 4801 9024 4813 9027
rect 3568 8996 4813 9024
rect 3568 8984 3574 8996
rect 4801 8993 4813 8996
rect 4847 8993 4859 9027
rect 4801 8987 4859 8993
rect 3602 8956 3608 8968
rect 3436 8928 3608 8956
rect 2685 8919 2743 8925
rect 3602 8916 3608 8928
rect 3660 8916 3666 8968
rect 4985 8959 5043 8965
rect 4985 8925 4997 8959
rect 5031 8956 5043 8959
rect 5166 8956 5172 8968
rect 5031 8928 5172 8956
rect 5031 8925 5043 8928
rect 4985 8919 5043 8925
rect 5166 8916 5172 8928
rect 5224 8916 5230 8968
rect 5353 8959 5411 8965
rect 5353 8925 5365 8959
rect 5399 8925 5411 8959
rect 5353 8919 5411 8925
rect 2774 8888 2780 8900
rect 2608 8860 2780 8888
rect 2774 8848 2780 8860
rect 2832 8848 2838 8900
rect 3418 8848 3424 8900
rect 3476 8888 3482 8900
rect 5368 8888 5396 8919
rect 5442 8916 5448 8968
rect 5500 8916 5506 8968
rect 3476 8860 5396 8888
rect 3476 8848 3482 8860
rect 2409 8823 2467 8829
rect 2409 8789 2421 8823
rect 2455 8789 2467 8823
rect 2409 8783 2467 8789
rect 2498 8780 2504 8832
rect 2556 8780 2562 8832
rect 3142 8780 3148 8832
rect 3200 8820 3206 8832
rect 3237 8823 3295 8829
rect 3237 8820 3249 8823
rect 3200 8792 3249 8820
rect 3200 8780 3206 8792
rect 3237 8789 3249 8792
rect 3283 8820 3295 8823
rect 3510 8820 3516 8832
rect 3283 8792 3516 8820
rect 3283 8789 3295 8792
rect 3237 8783 3295 8789
rect 3510 8780 3516 8792
rect 3568 8780 3574 8832
rect 3605 8823 3663 8829
rect 3605 8789 3617 8823
rect 3651 8820 3663 8823
rect 4341 8823 4399 8829
rect 4341 8820 4353 8823
rect 3651 8792 4353 8820
rect 3651 8789 3663 8792
rect 3605 8783 3663 8789
rect 4341 8789 4353 8792
rect 4387 8820 4399 8823
rect 4706 8820 4712 8832
rect 4387 8792 4712 8820
rect 4387 8789 4399 8792
rect 4341 8783 4399 8789
rect 4706 8780 4712 8792
rect 4764 8780 4770 8832
rect 5169 8823 5227 8829
rect 5169 8789 5181 8823
rect 5215 8820 5227 8823
rect 5534 8820 5540 8832
rect 5215 8792 5540 8820
rect 5215 8789 5227 8792
rect 5169 8783 5227 8789
rect 5534 8780 5540 8792
rect 5592 8780 5598 8832
rect 5736 8820 5764 9064
rect 5828 9024 5856 9120
rect 9048 9092 9076 9132
rect 9858 9120 9864 9132
rect 9916 9120 9922 9172
rect 10594 9120 10600 9172
rect 10652 9160 10658 9172
rect 23474 9160 23480 9172
rect 10652 9132 23480 9160
rect 10652 9120 10658 9132
rect 23474 9120 23480 9132
rect 23532 9120 23538 9172
rect 7208 9064 9076 9092
rect 6089 9027 6147 9033
rect 6089 9024 6101 9027
rect 5828 8996 6101 9024
rect 6089 8993 6101 8996
rect 6135 8993 6147 9027
rect 6089 8987 6147 8993
rect 5813 8959 5871 8965
rect 5813 8925 5825 8959
rect 5859 8925 5871 8959
rect 7208 8942 7236 9064
rect 10226 9052 10232 9104
rect 10284 9092 10290 9104
rect 10284 9064 19334 9092
rect 10284 9052 10290 9064
rect 7834 8984 7840 9036
rect 7892 8984 7898 9036
rect 8757 9027 8815 9033
rect 8757 8993 8769 9027
rect 8803 9024 8815 9027
rect 9306 9024 9312 9036
rect 8803 8996 9312 9024
rect 8803 8993 8815 8996
rect 8757 8987 8815 8993
rect 9306 8984 9312 8996
rect 9364 8984 9370 9036
rect 9674 8984 9680 9036
rect 9732 9024 9738 9036
rect 9732 8996 11192 9024
rect 9732 8984 9738 8996
rect 5813 8919 5871 8925
rect 5828 8888 5856 8919
rect 8938 8916 8944 8968
rect 8996 8916 9002 8968
rect 10594 8916 10600 8968
rect 10652 8956 10658 8968
rect 10873 8959 10931 8965
rect 10873 8956 10885 8959
rect 10652 8928 10885 8956
rect 10652 8916 10658 8928
rect 10873 8925 10885 8928
rect 10919 8925 10931 8959
rect 10873 8919 10931 8925
rect 5994 8888 6000 8900
rect 5828 8860 6000 8888
rect 5994 8848 6000 8860
rect 6052 8848 6058 8900
rect 9214 8848 9220 8900
rect 9272 8848 9278 8900
rect 9766 8848 9772 8900
rect 9824 8848 9830 8900
rect 10502 8820 10508 8832
rect 5736 8792 10508 8820
rect 10502 8780 10508 8792
rect 10560 8780 10566 8832
rect 10594 8780 10600 8832
rect 10652 8820 10658 8832
rect 10689 8823 10747 8829
rect 10689 8820 10701 8823
rect 10652 8792 10701 8820
rect 10652 8780 10658 8792
rect 10689 8789 10701 8792
rect 10735 8789 10747 8823
rect 10888 8820 10916 8919
rect 11054 8916 11060 8968
rect 11112 8916 11118 8968
rect 11164 8956 11192 8996
rect 12066 8984 12072 9036
rect 12124 8984 12130 9036
rect 19306 9024 19334 9064
rect 26602 9024 26608 9036
rect 19306 8996 26608 9024
rect 26602 8984 26608 8996
rect 26660 8984 26666 9036
rect 28353 9027 28411 9033
rect 28353 8993 28365 9027
rect 28399 9024 28411 9027
rect 28810 9024 28816 9036
rect 28399 8996 28816 9024
rect 28399 8993 28411 8996
rect 28353 8987 28411 8993
rect 28810 8984 28816 8996
rect 28868 8984 28874 9036
rect 12253 8959 12311 8965
rect 12253 8956 12265 8959
rect 11164 8928 12265 8956
rect 12253 8925 12265 8928
rect 12299 8925 12311 8959
rect 12253 8919 12311 8925
rect 27154 8916 27160 8968
rect 27212 8916 27218 8968
rect 11241 8891 11299 8897
rect 11241 8857 11253 8891
rect 11287 8888 11299 8891
rect 26878 8888 26884 8900
rect 11287 8860 26884 8888
rect 11287 8857 11299 8860
rect 11241 8851 11299 8857
rect 26878 8848 26884 8860
rect 26936 8848 26942 8900
rect 11609 8823 11667 8829
rect 11609 8820 11621 8823
rect 10888 8792 11621 8820
rect 10689 8783 10747 8789
rect 11609 8789 11621 8792
rect 11655 8789 11667 8823
rect 11609 8783 11667 8789
rect 12434 8780 12440 8832
rect 12492 8780 12498 8832
rect 1104 8730 29048 8752
rect 1104 8678 7896 8730
rect 7948 8678 7960 8730
rect 8012 8678 8024 8730
rect 8076 8678 8088 8730
rect 8140 8678 8152 8730
rect 8204 8678 14842 8730
rect 14894 8678 14906 8730
rect 14958 8678 14970 8730
rect 15022 8678 15034 8730
rect 15086 8678 15098 8730
rect 15150 8678 21788 8730
rect 21840 8678 21852 8730
rect 21904 8678 21916 8730
rect 21968 8678 21980 8730
rect 22032 8678 22044 8730
rect 22096 8678 28734 8730
rect 28786 8678 28798 8730
rect 28850 8678 28862 8730
rect 28914 8678 28926 8730
rect 28978 8678 28990 8730
rect 29042 8678 29048 8730
rect 1104 8656 29048 8678
rect 1578 8576 1584 8628
rect 1636 8576 1642 8628
rect 2409 8619 2467 8625
rect 2409 8616 2421 8619
rect 2148 8588 2421 8616
rect 1486 8508 1492 8560
rect 1544 8548 1550 8560
rect 2038 8548 2044 8560
rect 1544 8520 2044 8548
rect 1544 8508 1550 8520
rect 2038 8508 2044 8520
rect 2096 8508 2102 8560
rect 2148 8492 2176 8588
rect 2409 8585 2421 8588
rect 2455 8585 2467 8619
rect 2409 8579 2467 8585
rect 2774 8576 2780 8628
rect 2832 8576 2838 8628
rect 5902 8616 5908 8628
rect 3436 8588 5908 8616
rect 1394 8440 1400 8492
rect 1452 8440 1458 8492
rect 1670 8440 1676 8492
rect 1728 8440 1734 8492
rect 1949 8483 2007 8489
rect 1949 8480 1961 8483
rect 1780 8452 1961 8480
rect 750 8372 756 8424
rect 808 8412 814 8424
rect 1026 8412 1032 8424
rect 808 8384 1032 8412
rect 808 8372 814 8384
rect 1026 8372 1032 8384
rect 1084 8372 1090 8424
rect 1780 8412 1808 8452
rect 1949 8449 1961 8452
rect 1995 8449 2007 8483
rect 1949 8443 2007 8449
rect 2130 8440 2136 8492
rect 2188 8440 2194 8492
rect 2225 8483 2283 8489
rect 2225 8449 2237 8483
rect 2271 8480 2283 8483
rect 2314 8480 2320 8492
rect 2271 8452 2320 8480
rect 2271 8449 2283 8452
rect 2225 8443 2283 8449
rect 2314 8440 2320 8452
rect 2372 8440 2378 8492
rect 2685 8483 2743 8489
rect 2685 8449 2697 8483
rect 2731 8480 2743 8483
rect 2866 8480 2872 8492
rect 2731 8452 2872 8480
rect 2731 8449 2743 8452
rect 2685 8443 2743 8449
rect 2866 8440 2872 8452
rect 2924 8440 2930 8492
rect 2958 8440 2964 8492
rect 3016 8440 3022 8492
rect 3142 8440 3148 8492
rect 3200 8480 3206 8492
rect 3237 8483 3295 8489
rect 3237 8480 3249 8483
rect 3200 8452 3249 8480
rect 3200 8440 3206 8452
rect 3237 8449 3249 8452
rect 3283 8449 3295 8483
rect 3237 8443 3295 8449
rect 3326 8440 3332 8492
rect 3384 8440 3390 8492
rect 3436 8412 3464 8588
rect 5902 8576 5908 8588
rect 5960 8576 5966 8628
rect 6178 8576 6184 8628
rect 6236 8616 6242 8628
rect 6365 8619 6423 8625
rect 6365 8616 6377 8619
rect 6236 8588 6377 8616
rect 6236 8576 6242 8588
rect 6365 8585 6377 8588
rect 6411 8585 6423 8619
rect 6365 8579 6423 8585
rect 6733 8619 6791 8625
rect 6733 8585 6745 8619
rect 6779 8616 6791 8619
rect 7193 8619 7251 8625
rect 6779 8588 7144 8616
rect 6779 8585 6791 8588
rect 6733 8579 6791 8585
rect 4982 8508 4988 8560
rect 5040 8548 5046 8560
rect 5445 8551 5503 8557
rect 5445 8548 5457 8551
rect 5040 8520 5457 8548
rect 5040 8508 5046 8520
rect 5445 8517 5457 8520
rect 5491 8517 5503 8551
rect 5445 8511 5503 8517
rect 5534 8508 5540 8560
rect 5592 8548 5598 8560
rect 6825 8551 6883 8557
rect 6825 8548 6837 8551
rect 5592 8520 6837 8548
rect 5592 8508 5598 8520
rect 6825 8517 6837 8520
rect 6871 8517 6883 8551
rect 7116 8548 7144 8588
rect 7193 8585 7205 8619
rect 7239 8616 7251 8619
rect 7282 8616 7288 8628
rect 7239 8588 7288 8616
rect 7239 8585 7251 8588
rect 7193 8579 7251 8585
rect 7282 8576 7288 8588
rect 7340 8576 7346 8628
rect 7742 8576 7748 8628
rect 7800 8576 7806 8628
rect 8570 8576 8576 8628
rect 8628 8576 8634 8628
rect 9214 8576 9220 8628
rect 9272 8616 9278 8628
rect 9493 8619 9551 8625
rect 9493 8616 9505 8619
rect 9272 8588 9505 8616
rect 9272 8576 9278 8588
rect 9493 8585 9505 8588
rect 9539 8585 9551 8619
rect 9493 8579 9551 8585
rect 10594 8576 10600 8628
rect 10652 8576 10658 8628
rect 10689 8619 10747 8625
rect 10689 8585 10701 8619
rect 10735 8616 10747 8619
rect 10778 8616 10784 8628
rect 10735 8588 10784 8616
rect 10735 8585 10747 8588
rect 10689 8579 10747 8585
rect 10778 8576 10784 8588
rect 10836 8576 10842 8628
rect 11146 8576 11152 8628
rect 11204 8616 11210 8628
rect 11517 8619 11575 8625
rect 11517 8616 11529 8619
rect 11204 8588 11529 8616
rect 11204 8576 11210 8588
rect 11517 8585 11529 8588
rect 11563 8585 11575 8619
rect 27154 8616 27160 8628
rect 11517 8579 11575 8585
rect 12406 8588 27160 8616
rect 7760 8548 7788 8576
rect 7116 8520 7788 8548
rect 9033 8551 9091 8557
rect 6825 8511 6883 8517
rect 9033 8517 9045 8551
rect 9079 8548 9091 8551
rect 10612 8548 10640 8576
rect 12406 8548 12434 8588
rect 27154 8576 27160 8588
rect 27212 8576 27218 8628
rect 9079 8520 12434 8548
rect 9079 8517 9091 8520
rect 9033 8511 9091 8517
rect 3694 8440 3700 8492
rect 3752 8480 3758 8492
rect 4893 8483 4951 8489
rect 4893 8480 4905 8483
rect 3752 8452 4905 8480
rect 3752 8440 3758 8452
rect 4893 8449 4905 8452
rect 4939 8449 4951 8483
rect 4893 8443 4951 8449
rect 5077 8483 5135 8489
rect 5077 8449 5089 8483
rect 5123 8480 5135 8483
rect 5166 8480 5172 8492
rect 5123 8452 5172 8480
rect 5123 8449 5135 8452
rect 5077 8443 5135 8449
rect 5166 8440 5172 8452
rect 5224 8440 5230 8492
rect 7374 8480 7380 8492
rect 6012 8452 7380 8480
rect 6012 8412 6040 8452
rect 7374 8440 7380 8452
rect 7432 8440 7438 8492
rect 10336 8489 10364 8520
rect 17218 8508 17224 8560
rect 17276 8508 17282 8560
rect 8021 8483 8079 8489
rect 8021 8449 8033 8483
rect 8067 8480 8079 8483
rect 10321 8483 10379 8489
rect 8067 8452 10272 8480
rect 8067 8449 8079 8452
rect 8021 8443 8079 8449
rect 1136 8384 1808 8412
rect 2240 8384 3464 8412
rect 3528 8384 6040 8412
rect 1136 8344 1164 8384
rect 1044 8316 1164 8344
rect 1857 8347 1915 8353
rect 1044 8288 1072 8316
rect 1857 8313 1869 8347
rect 1903 8344 1915 8347
rect 2240 8344 2268 8384
rect 1903 8316 2268 8344
rect 1903 8313 1915 8316
rect 1857 8307 1915 8313
rect 2314 8304 2320 8356
rect 2372 8344 2378 8356
rect 2501 8347 2559 8353
rect 2501 8344 2513 8347
rect 2372 8316 2513 8344
rect 2372 8304 2378 8316
rect 2501 8313 2513 8316
rect 2547 8313 2559 8347
rect 2501 8307 2559 8313
rect 3050 8304 3056 8356
rect 3108 8304 3114 8356
rect 3528 8353 3556 8384
rect 6086 8372 6092 8424
rect 6144 8372 6150 8424
rect 6270 8372 6276 8424
rect 6328 8412 6334 8424
rect 6917 8415 6975 8421
rect 6917 8412 6929 8415
rect 6328 8384 6929 8412
rect 6328 8372 6334 8384
rect 6917 8381 6929 8384
rect 6963 8381 6975 8415
rect 6917 8375 6975 8381
rect 7742 8372 7748 8424
rect 7800 8372 7806 8424
rect 8570 8372 8576 8424
rect 8628 8412 8634 8424
rect 8757 8415 8815 8421
rect 8757 8412 8769 8415
rect 8628 8384 8769 8412
rect 8628 8372 8634 8384
rect 8757 8381 8769 8384
rect 8803 8381 8815 8415
rect 8757 8375 8815 8381
rect 8941 8415 8999 8421
rect 8941 8381 8953 8415
rect 8987 8381 8999 8415
rect 10045 8415 10103 8421
rect 10045 8412 10057 8415
rect 8941 8375 8999 8381
rect 9416 8384 10057 8412
rect 3513 8347 3571 8353
rect 3513 8313 3525 8347
rect 3559 8313 3571 8347
rect 3513 8307 3571 8313
rect 4065 8347 4123 8353
rect 4065 8313 4077 8347
rect 4111 8344 4123 8347
rect 4433 8347 4491 8353
rect 4111 8316 4292 8344
rect 4111 8313 4123 8316
rect 4065 8307 4123 8313
rect 4264 8288 4292 8316
rect 4433 8313 4445 8347
rect 4479 8344 4491 8347
rect 4706 8344 4712 8356
rect 4479 8316 4712 8344
rect 4479 8313 4491 8316
rect 4433 8307 4491 8313
rect 4706 8304 4712 8316
rect 4764 8304 4770 8356
rect 4801 8347 4859 8353
rect 4801 8313 4813 8347
rect 4847 8344 4859 8347
rect 5261 8347 5319 8353
rect 4847 8316 5212 8344
rect 4847 8313 4859 8316
rect 4801 8307 4859 8313
rect 1026 8236 1032 8288
rect 1084 8236 1090 8288
rect 1578 8236 1584 8288
rect 1636 8276 1642 8288
rect 1946 8276 1952 8288
rect 1636 8248 1952 8276
rect 1636 8236 1642 8248
rect 1946 8236 1952 8248
rect 2004 8236 2010 8288
rect 2038 8236 2044 8288
rect 2096 8276 2102 8288
rect 2133 8279 2191 8285
rect 2133 8276 2145 8279
rect 2096 8248 2145 8276
rect 2096 8236 2102 8248
rect 2133 8245 2145 8248
rect 2179 8245 2191 8279
rect 2133 8239 2191 8245
rect 4246 8236 4252 8288
rect 4304 8236 4310 8288
rect 5184 8276 5212 8316
rect 5261 8313 5273 8347
rect 5307 8344 5319 8347
rect 8956 8344 8984 8375
rect 9416 8353 9444 8384
rect 10045 8381 10057 8384
rect 10091 8381 10103 8415
rect 10244 8412 10272 8452
rect 10321 8449 10333 8483
rect 10367 8449 10379 8483
rect 10321 8443 10379 8449
rect 10413 8483 10471 8489
rect 10413 8449 10425 8483
rect 10459 8480 10471 8483
rect 10502 8480 10508 8492
rect 10459 8452 10508 8480
rect 10459 8449 10471 8452
rect 10413 8443 10471 8449
rect 10502 8440 10508 8452
rect 10560 8440 10566 8492
rect 10597 8483 10655 8489
rect 10597 8449 10609 8483
rect 10643 8480 10655 8483
rect 17236 8480 17264 8508
rect 27157 8483 27215 8489
rect 27157 8480 27169 8483
rect 10643 8452 17264 8480
rect 26712 8452 27169 8480
rect 10643 8449 10655 8452
rect 10597 8443 10655 8449
rect 11054 8412 11060 8424
rect 10244 8384 11060 8412
rect 10045 8375 10103 8381
rect 11054 8372 11060 8384
rect 11112 8372 11118 8424
rect 11238 8372 11244 8424
rect 11296 8372 11302 8424
rect 12158 8372 12164 8424
rect 12216 8372 12222 8424
rect 26712 8353 26740 8452
rect 27157 8449 27169 8452
rect 27203 8449 27215 8483
rect 27157 8443 27215 8449
rect 28350 8372 28356 8424
rect 28408 8372 28414 8424
rect 5307 8316 8984 8344
rect 9401 8347 9459 8353
rect 5307 8313 5319 8316
rect 5261 8307 5319 8313
rect 9401 8313 9413 8347
rect 9447 8313 9459 8347
rect 26697 8347 26755 8353
rect 26697 8344 26709 8347
rect 9401 8307 9459 8313
rect 23400 8316 26709 8344
rect 23400 8288 23428 8316
rect 26697 8313 26709 8316
rect 26743 8313 26755 8347
rect 26697 8307 26755 8313
rect 7650 8276 7656 8288
rect 5184 8248 7656 8276
rect 7650 8236 7656 8248
rect 7708 8236 7714 8288
rect 23382 8236 23388 8288
rect 23440 8236 23446 8288
rect 1104 8186 28888 8208
rect 1104 8134 4423 8186
rect 4475 8134 4487 8186
rect 4539 8134 4551 8186
rect 4603 8134 4615 8186
rect 4667 8134 4679 8186
rect 4731 8134 11369 8186
rect 11421 8134 11433 8186
rect 11485 8134 11497 8186
rect 11549 8134 11561 8186
rect 11613 8134 11625 8186
rect 11677 8134 18315 8186
rect 18367 8134 18379 8186
rect 18431 8134 18443 8186
rect 18495 8134 18507 8186
rect 18559 8134 18571 8186
rect 18623 8134 25261 8186
rect 25313 8134 25325 8186
rect 25377 8134 25389 8186
rect 25441 8134 25453 8186
rect 25505 8134 25517 8186
rect 25569 8134 28888 8186
rect 1104 8112 28888 8134
rect 1394 8032 1400 8084
rect 1452 8072 1458 8084
rect 1670 8072 1676 8084
rect 1452 8044 1676 8072
rect 1452 8032 1458 8044
rect 1670 8032 1676 8044
rect 1728 8032 1734 8084
rect 5074 8072 5080 8084
rect 4632 8044 5080 8072
rect 474 7964 480 8016
rect 532 8004 538 8016
rect 532 7976 3832 8004
rect 532 7964 538 7976
rect 768 7908 2544 7936
rect 768 7608 796 7908
rect 1394 7828 1400 7880
rect 1452 7828 1458 7880
rect 1578 7828 1584 7880
rect 1636 7868 1642 7880
rect 1765 7871 1823 7877
rect 1765 7868 1777 7871
rect 1636 7840 1777 7868
rect 1636 7828 1642 7840
rect 1765 7837 1777 7840
rect 1811 7837 1823 7871
rect 1765 7831 1823 7837
rect 2038 7828 2044 7880
rect 2096 7868 2102 7880
rect 2516 7877 2544 7908
rect 3234 7896 3240 7948
rect 3292 7896 3298 7948
rect 3804 7945 3832 7976
rect 3789 7939 3847 7945
rect 3789 7905 3801 7939
rect 3835 7905 3847 7939
rect 3789 7899 3847 7905
rect 3878 7896 3884 7948
rect 3936 7936 3942 7948
rect 4154 7936 4160 7948
rect 3936 7908 4160 7936
rect 3936 7896 3942 7908
rect 4154 7896 4160 7908
rect 4212 7936 4218 7948
rect 4632 7945 4660 8044
rect 5074 8032 5080 8044
rect 5132 8032 5138 8084
rect 5626 8072 5632 8084
rect 5276 8044 5632 8072
rect 5276 8004 5304 8044
rect 5626 8032 5632 8044
rect 5684 8032 5690 8084
rect 5902 8032 5908 8084
rect 5960 8072 5966 8084
rect 5960 8044 6500 8072
rect 5960 8032 5966 8044
rect 6472 8016 6500 8044
rect 7190 8032 7196 8084
rect 7248 8072 7254 8084
rect 8573 8075 8631 8081
rect 8573 8072 8585 8075
rect 7248 8044 8585 8072
rect 7248 8032 7254 8044
rect 8573 8041 8585 8044
rect 8619 8041 8631 8075
rect 8573 8035 8631 8041
rect 8941 8075 8999 8081
rect 8941 8041 8953 8075
rect 8987 8072 8999 8075
rect 9122 8072 9128 8084
rect 8987 8044 9128 8072
rect 8987 8041 8999 8044
rect 8941 8035 8999 8041
rect 9122 8032 9128 8044
rect 9180 8032 9186 8084
rect 10962 8032 10968 8084
rect 11020 8072 11026 8084
rect 11057 8075 11115 8081
rect 11057 8072 11069 8075
rect 11020 8044 11069 8072
rect 11020 8032 11026 8044
rect 11057 8041 11069 8044
rect 11103 8041 11115 8075
rect 11057 8035 11115 8041
rect 13170 8032 13176 8084
rect 13228 8072 13234 8084
rect 26973 8075 27031 8081
rect 26973 8072 26985 8075
rect 13228 8044 26985 8072
rect 13228 8032 13234 8044
rect 26973 8041 26985 8044
rect 27019 8072 27031 8075
rect 27154 8072 27160 8084
rect 27019 8044 27160 8072
rect 27019 8041 27031 8044
rect 26973 8035 27031 8041
rect 27154 8032 27160 8044
rect 27212 8032 27218 8084
rect 4724 7976 5304 8004
rect 4617 7939 4675 7945
rect 4212 7908 4384 7936
rect 4212 7896 4218 7908
rect 2225 7871 2283 7877
rect 2225 7868 2237 7871
rect 2096 7840 2237 7868
rect 2096 7828 2102 7840
rect 2225 7837 2237 7840
rect 2271 7837 2283 7871
rect 2225 7831 2283 7837
rect 2501 7871 2559 7877
rect 2501 7837 2513 7871
rect 2547 7837 2559 7871
rect 2501 7831 2559 7837
rect 2961 7871 3019 7877
rect 2961 7837 2973 7871
rect 3007 7868 3019 7871
rect 3007 7840 3372 7868
rect 3007 7837 3019 7840
rect 2961 7831 3019 7837
rect 1412 7800 1440 7828
rect 1946 7800 1952 7812
rect 1412 7772 1952 7800
rect 1946 7760 1952 7772
rect 2004 7760 2010 7812
rect 1397 7735 1455 7741
rect 1397 7732 1409 7735
rect 860 7704 1409 7732
rect 750 7556 756 7608
rect 808 7556 814 7608
rect 658 7488 664 7540
rect 716 7528 722 7540
rect 860 7528 888 7704
rect 1397 7701 1409 7704
rect 1443 7701 1455 7735
rect 1397 7695 1455 7701
rect 1578 7692 1584 7744
rect 1636 7692 1642 7744
rect 1673 7735 1731 7741
rect 1673 7701 1685 7735
rect 1719 7732 1731 7735
rect 2130 7732 2136 7744
rect 1719 7704 2136 7732
rect 1719 7701 1731 7704
rect 1673 7695 1731 7701
rect 2130 7692 2136 7704
rect 2188 7692 2194 7744
rect 2406 7692 2412 7744
rect 2464 7692 2470 7744
rect 2682 7692 2688 7744
rect 2740 7692 2746 7744
rect 3053 7735 3111 7741
rect 3053 7701 3065 7735
rect 3099 7732 3111 7735
rect 3142 7732 3148 7744
rect 3099 7704 3148 7732
rect 3099 7701 3111 7704
rect 3053 7695 3111 7701
rect 3142 7692 3148 7704
rect 3200 7692 3206 7744
rect 3344 7732 3372 7840
rect 3418 7828 3424 7880
rect 3476 7828 3482 7880
rect 3970 7828 3976 7880
rect 4028 7828 4034 7880
rect 4356 7877 4384 7908
rect 4617 7905 4629 7939
rect 4663 7905 4675 7939
rect 4617 7899 4675 7905
rect 4341 7871 4399 7877
rect 4341 7837 4353 7871
rect 4387 7837 4399 7871
rect 4341 7831 4399 7837
rect 3605 7803 3663 7809
rect 3605 7769 3617 7803
rect 3651 7800 3663 7803
rect 4724 7800 4752 7976
rect 6454 7964 6460 8016
rect 6512 7964 6518 8016
rect 7745 8007 7803 8013
rect 7392 7976 7696 8004
rect 4982 7896 4988 7948
rect 5040 7936 5046 7948
rect 7392 7945 7420 7976
rect 7668 7948 7696 7976
rect 7745 7973 7757 8007
rect 7791 8004 7803 8007
rect 7791 7976 12204 8004
rect 7791 7973 7803 7976
rect 7745 7967 7803 7973
rect 5445 7939 5503 7945
rect 5445 7936 5457 7939
rect 5040 7908 5457 7936
rect 5040 7896 5046 7908
rect 5445 7905 5457 7908
rect 5491 7905 5503 7939
rect 5445 7899 5503 7905
rect 7377 7939 7435 7945
rect 7377 7905 7389 7939
rect 7423 7905 7435 7939
rect 7377 7899 7435 7905
rect 7650 7896 7656 7948
rect 7708 7936 7714 7948
rect 8202 7936 8208 7948
rect 7708 7908 8208 7936
rect 7708 7896 7714 7908
rect 8202 7896 8208 7908
rect 8260 7896 8266 7948
rect 8294 7896 8300 7948
rect 8352 7936 8358 7948
rect 12176 7936 12204 7976
rect 12250 7964 12256 8016
rect 12308 8004 12314 8016
rect 23382 8004 23388 8016
rect 12308 7976 23388 8004
rect 12308 7964 12314 7976
rect 23382 7964 23388 7976
rect 23440 7964 23446 8016
rect 8352 7908 9904 7936
rect 12176 7908 14688 7936
rect 8352 7896 8358 7908
rect 4801 7871 4859 7877
rect 4801 7837 4813 7871
rect 4847 7837 4859 7871
rect 4801 7831 4859 7837
rect 3651 7772 4752 7800
rect 4816 7800 4844 7831
rect 5074 7828 5080 7880
rect 5132 7868 5138 7880
rect 5169 7871 5227 7877
rect 5169 7868 5181 7871
rect 5132 7840 5181 7868
rect 5132 7828 5138 7840
rect 5169 7837 5181 7840
rect 5215 7837 5227 7871
rect 5169 7831 5227 7837
rect 6730 7828 6736 7880
rect 6788 7868 6794 7880
rect 7561 7871 7619 7877
rect 7561 7868 7573 7871
rect 6788 7840 7573 7868
rect 6788 7828 6794 7840
rect 7561 7837 7573 7840
rect 7607 7837 7619 7871
rect 7561 7831 7619 7837
rect 7929 7871 7987 7877
rect 7929 7837 7941 7871
rect 7975 7837 7987 7871
rect 7929 7831 7987 7837
rect 9585 7871 9643 7877
rect 9585 7837 9597 7871
rect 9631 7868 9643 7871
rect 9674 7868 9680 7880
rect 9631 7840 9680 7868
rect 9631 7837 9643 7840
rect 9585 7831 9643 7837
rect 5534 7800 5540 7812
rect 4816 7772 5540 7800
rect 3651 7769 3663 7772
rect 3605 7763 3663 7769
rect 5534 7760 5540 7772
rect 5592 7760 5598 7812
rect 7006 7800 7012 7812
rect 6670 7772 7012 7800
rect 7006 7760 7012 7772
rect 7064 7760 7070 7812
rect 7193 7803 7251 7809
rect 7193 7769 7205 7803
rect 7239 7769 7251 7803
rect 7193 7763 7251 7769
rect 3510 7732 3516 7744
rect 3344 7704 3516 7732
rect 3510 7692 3516 7704
rect 3568 7732 3574 7744
rect 3878 7732 3884 7744
rect 3568 7704 3884 7732
rect 3568 7692 3574 7704
rect 3878 7692 3884 7704
rect 3936 7692 3942 7744
rect 4154 7692 4160 7744
rect 4212 7692 4218 7744
rect 4433 7735 4491 7741
rect 4433 7701 4445 7735
rect 4479 7732 4491 7735
rect 4798 7732 4804 7744
rect 4479 7704 4804 7732
rect 4479 7701 4491 7704
rect 4433 7695 4491 7701
rect 4798 7692 4804 7704
rect 4856 7692 4862 7744
rect 4982 7692 4988 7744
rect 5040 7692 5046 7744
rect 5718 7692 5724 7744
rect 5776 7732 5782 7744
rect 7208 7732 7236 7763
rect 7282 7760 7288 7812
rect 7340 7800 7346 7812
rect 7944 7800 7972 7831
rect 9674 7828 9680 7840
rect 9732 7828 9738 7880
rect 9876 7877 9904 7908
rect 9769 7871 9827 7877
rect 9769 7837 9781 7871
rect 9815 7837 9827 7871
rect 9769 7831 9827 7837
rect 9861 7871 9919 7877
rect 9861 7837 9873 7871
rect 9907 7837 9919 7871
rect 9861 7831 9919 7837
rect 7340 7772 7972 7800
rect 7340 7760 7346 7772
rect 8570 7760 8576 7812
rect 8628 7800 8634 7812
rect 9122 7800 9128 7812
rect 8628 7772 9128 7800
rect 8628 7760 8634 7772
rect 9122 7760 9128 7772
rect 9180 7760 9186 7812
rect 9784 7800 9812 7831
rect 10410 7828 10416 7880
rect 10468 7828 10474 7880
rect 10502 7828 10508 7880
rect 10560 7828 10566 7880
rect 10686 7828 10692 7880
rect 10744 7868 10750 7880
rect 10965 7871 11023 7877
rect 10965 7868 10977 7871
rect 10744 7840 10977 7868
rect 10744 7828 10750 7840
rect 10965 7837 10977 7840
rect 11011 7837 11023 7871
rect 10965 7831 11023 7837
rect 11701 7871 11759 7877
rect 11701 7837 11713 7871
rect 11747 7868 11759 7871
rect 12526 7868 12532 7880
rect 11747 7840 12532 7868
rect 11747 7837 11759 7840
rect 11701 7831 11759 7837
rect 12526 7828 12532 7840
rect 12584 7828 12590 7880
rect 10520 7800 10548 7828
rect 14660 7812 14688 7908
rect 27614 7896 27620 7948
rect 27672 7896 27678 7948
rect 15470 7828 15476 7880
rect 15528 7868 15534 7880
rect 27157 7871 27215 7877
rect 27157 7868 27169 7871
rect 15528 7840 27169 7868
rect 15528 7828 15534 7840
rect 27157 7837 27169 7840
rect 27203 7837 27215 7871
rect 27157 7831 27215 7837
rect 9646 7772 10548 7800
rect 9646 7732 9674 7772
rect 14642 7760 14648 7812
rect 14700 7760 14706 7812
rect 5776 7704 9674 7732
rect 5776 7692 5782 7704
rect 10042 7692 10048 7744
rect 10100 7692 10106 7744
rect 1104 7642 29048 7664
rect 1104 7590 7896 7642
rect 7948 7590 7960 7642
rect 8012 7590 8024 7642
rect 8076 7590 8088 7642
rect 8140 7590 8152 7642
rect 8204 7590 14842 7642
rect 14894 7590 14906 7642
rect 14958 7590 14970 7642
rect 15022 7590 15034 7642
rect 15086 7590 15098 7642
rect 15150 7590 21788 7642
rect 21840 7590 21852 7642
rect 21904 7590 21916 7642
rect 21968 7590 21980 7642
rect 22032 7590 22044 7642
rect 22096 7590 28734 7642
rect 28786 7590 28798 7642
rect 28850 7590 28862 7642
rect 28914 7590 28926 7642
rect 28978 7590 28990 7642
rect 29042 7590 29048 7642
rect 1104 7568 29048 7590
rect 716 7500 888 7528
rect 716 7488 722 7500
rect 1762 7488 1768 7540
rect 1820 7488 1826 7540
rect 3237 7531 3295 7537
rect 3237 7497 3249 7531
rect 3283 7528 3295 7531
rect 3970 7528 3976 7540
rect 3283 7500 3976 7528
rect 3283 7497 3295 7500
rect 3237 7491 3295 7497
rect 3970 7488 3976 7500
rect 4028 7488 4034 7540
rect 4246 7488 4252 7540
rect 4304 7488 4310 7540
rect 4982 7488 4988 7540
rect 5040 7528 5046 7540
rect 5905 7531 5963 7537
rect 5905 7528 5917 7531
rect 5040 7500 5917 7528
rect 5040 7488 5046 7500
rect 5905 7497 5917 7500
rect 5951 7497 5963 7531
rect 5905 7491 5963 7497
rect 6178 7488 6184 7540
rect 6236 7528 6242 7540
rect 6365 7531 6423 7537
rect 6365 7528 6377 7531
rect 6236 7500 6377 7528
rect 6236 7488 6242 7500
rect 6365 7497 6377 7500
rect 6411 7497 6423 7531
rect 6365 7491 6423 7497
rect 6914 7488 6920 7540
rect 6972 7488 6978 7540
rect 7006 7488 7012 7540
rect 7064 7528 7070 7540
rect 8021 7531 8079 7537
rect 8021 7528 8033 7531
rect 7064 7500 8033 7528
rect 7064 7488 7070 7500
rect 8021 7497 8033 7500
rect 8067 7497 8079 7531
rect 8021 7491 8079 7497
rect 8205 7531 8263 7537
rect 8205 7497 8217 7531
rect 8251 7528 8263 7531
rect 8386 7528 8392 7540
rect 8251 7500 8392 7528
rect 8251 7497 8263 7500
rect 8205 7491 8263 7497
rect 8386 7488 8392 7500
rect 8444 7488 8450 7540
rect 8772 7500 9720 7528
rect 1210 7420 1216 7472
rect 1268 7460 1274 7472
rect 3329 7463 3387 7469
rect 1268 7432 1716 7460
rect 1268 7420 1274 7432
rect 934 7352 940 7404
rect 992 7392 998 7404
rect 1581 7395 1639 7401
rect 1581 7392 1593 7395
rect 992 7364 1593 7392
rect 992 7352 998 7364
rect 1581 7361 1593 7364
rect 1627 7361 1639 7395
rect 1688 7392 1716 7432
rect 1872 7432 2728 7460
rect 1872 7392 1900 7432
rect 1688 7364 1900 7392
rect 1581 7355 1639 7361
rect 2498 7352 2504 7404
rect 2556 7392 2562 7404
rect 2593 7395 2651 7401
rect 2593 7392 2605 7395
rect 2556 7364 2605 7392
rect 2556 7352 2562 7364
rect 2593 7361 2605 7364
rect 2639 7361 2651 7395
rect 2700 7392 2728 7432
rect 3329 7429 3341 7463
rect 3375 7460 3387 7463
rect 3602 7460 3608 7472
rect 3375 7432 3608 7460
rect 3375 7429 3387 7432
rect 3329 7423 3387 7429
rect 3602 7420 3608 7432
rect 3660 7420 3666 7472
rect 4264 7460 4292 7488
rect 4264 7432 5028 7460
rect 5000 7401 5028 7432
rect 5718 7420 5724 7472
rect 5776 7460 5782 7472
rect 5813 7463 5871 7469
rect 5813 7460 5825 7463
rect 5776 7432 5825 7460
rect 5776 7420 5782 7432
rect 5813 7429 5825 7432
rect 5859 7429 5871 7463
rect 6822 7460 6828 7472
rect 5813 7423 5871 7429
rect 5920 7432 6828 7460
rect 4157 7395 4215 7401
rect 4157 7392 4169 7395
rect 2700 7364 4169 7392
rect 2593 7355 2651 7361
rect 4157 7361 4169 7364
rect 4203 7361 4215 7395
rect 4157 7355 4215 7361
rect 4341 7395 4399 7401
rect 4341 7361 4353 7395
rect 4387 7361 4399 7395
rect 4341 7355 4399 7361
rect 4525 7395 4583 7401
rect 4525 7361 4537 7395
rect 4571 7392 4583 7395
rect 4893 7395 4951 7401
rect 4893 7392 4905 7395
rect 4571 7364 4905 7392
rect 4571 7361 4583 7364
rect 4525 7355 4583 7361
rect 4893 7361 4905 7364
rect 4939 7361 4951 7395
rect 4893 7355 4951 7361
rect 4985 7395 5043 7401
rect 4985 7361 4997 7395
rect 5031 7392 5043 7395
rect 5920 7392 5948 7432
rect 6822 7420 6828 7432
rect 6880 7420 6886 7472
rect 6932 7460 6960 7488
rect 7101 7463 7159 7469
rect 7101 7460 7113 7463
rect 6932 7432 7113 7460
rect 7101 7429 7113 7432
rect 7147 7429 7159 7463
rect 8570 7460 8576 7472
rect 7101 7423 7159 7429
rect 7208 7432 8576 7460
rect 6270 7392 6276 7404
rect 5031 7364 5948 7392
rect 6012 7364 6276 7392
rect 5031 7361 5043 7364
rect 4985 7355 5043 7361
rect 1946 7284 1952 7336
rect 2004 7284 2010 7336
rect 3602 7284 3608 7336
rect 3660 7324 3666 7336
rect 3881 7327 3939 7333
rect 3881 7324 3893 7327
rect 3660 7296 3893 7324
rect 3660 7284 3666 7296
rect 3881 7293 3893 7296
rect 3927 7293 3939 7327
rect 3881 7287 3939 7293
rect 4062 7284 4068 7336
rect 4120 7324 4126 7336
rect 4356 7324 4384 7355
rect 4120 7296 4384 7324
rect 4120 7284 4126 7296
rect 4706 7284 4712 7336
rect 4764 7324 4770 7336
rect 6012 7333 6040 7364
rect 6270 7352 6276 7364
rect 6328 7352 6334 7404
rect 6454 7352 6460 7404
rect 6512 7392 6518 7404
rect 7208 7392 7236 7432
rect 8570 7420 8576 7432
rect 8628 7420 8634 7472
rect 8113 7395 8171 7401
rect 8113 7392 8125 7395
rect 6512 7364 7236 7392
rect 7392 7364 8125 7392
rect 6512 7352 6518 7364
rect 4801 7327 4859 7333
rect 4801 7324 4813 7327
rect 4764 7296 4813 7324
rect 4764 7284 4770 7296
rect 4801 7293 4813 7296
rect 4847 7324 4859 7327
rect 5997 7327 6055 7333
rect 5997 7324 6009 7327
rect 4847 7296 6009 7324
rect 4847 7293 4859 7296
rect 4801 7287 4859 7293
rect 1578 7216 1584 7268
rect 1636 7216 1642 7268
rect 2498 7216 2504 7268
rect 2556 7216 2562 7268
rect 1596 7188 1624 7216
rect 5000 7200 5028 7296
rect 5997 7293 6009 7296
rect 6043 7293 6055 7327
rect 5997 7287 6055 7293
rect 6086 7284 6092 7336
rect 6144 7284 6150 7336
rect 5353 7259 5411 7265
rect 5353 7225 5365 7259
rect 5399 7256 5411 7259
rect 5902 7256 5908 7268
rect 5399 7228 5908 7256
rect 5399 7225 5411 7228
rect 5353 7219 5411 7225
rect 5902 7216 5908 7228
rect 5960 7216 5966 7268
rect 3694 7188 3700 7200
rect 1596 7160 3700 7188
rect 3694 7148 3700 7160
rect 3752 7148 3758 7200
rect 4982 7148 4988 7200
rect 5040 7148 5046 7200
rect 5445 7191 5503 7197
rect 5445 7157 5457 7191
rect 5491 7188 5503 7191
rect 6104 7188 6132 7284
rect 5491 7160 6132 7188
rect 6288 7188 6316 7352
rect 7006 7284 7012 7336
rect 7064 7284 7070 7336
rect 6546 7216 6552 7268
rect 6604 7256 6610 7268
rect 7392 7256 7420 7364
rect 8113 7361 8125 7364
rect 8159 7392 8171 7395
rect 8772 7392 8800 7500
rect 9692 7460 9720 7500
rect 9766 7488 9772 7540
rect 9824 7488 9830 7540
rect 10042 7488 10048 7540
rect 10100 7528 10106 7540
rect 24394 7528 24400 7540
rect 10100 7500 24400 7528
rect 10100 7488 10106 7500
rect 24394 7488 24400 7500
rect 24452 7488 24458 7540
rect 9692 7432 10180 7460
rect 8159 7364 8800 7392
rect 8159 7361 8171 7364
rect 8113 7355 8171 7361
rect 9122 7352 9128 7404
rect 9180 7352 9186 7404
rect 9214 7352 9220 7404
rect 9272 7392 9278 7404
rect 9398 7392 9404 7404
rect 9272 7364 9404 7392
rect 9272 7352 9278 7364
rect 9398 7352 9404 7364
rect 9456 7352 9462 7404
rect 9692 7401 9720 7432
rect 9677 7395 9735 7401
rect 9677 7361 9689 7395
rect 9723 7361 9735 7395
rect 9677 7355 9735 7361
rect 9858 7352 9864 7404
rect 9916 7392 9922 7404
rect 10152 7401 10180 7432
rect 10502 7420 10508 7472
rect 10560 7460 10566 7472
rect 12250 7460 12256 7472
rect 10560 7432 12256 7460
rect 10560 7420 10566 7432
rect 12250 7420 12256 7432
rect 12308 7420 12314 7472
rect 26605 7463 26663 7469
rect 26605 7429 26617 7463
rect 26651 7460 26663 7463
rect 29178 7460 29184 7472
rect 26651 7432 29184 7460
rect 26651 7429 26663 7432
rect 26605 7423 26663 7429
rect 29178 7420 29184 7432
rect 29236 7420 29242 7472
rect 10045 7395 10103 7401
rect 10045 7392 10057 7395
rect 9916 7364 10057 7392
rect 9916 7352 9922 7364
rect 10045 7361 10057 7364
rect 10091 7361 10103 7395
rect 10045 7355 10103 7361
rect 10137 7395 10195 7401
rect 10137 7361 10149 7395
rect 10183 7392 10195 7395
rect 10318 7392 10324 7404
rect 10183 7364 10324 7392
rect 10183 7361 10195 7364
rect 10137 7355 10195 7361
rect 10318 7352 10324 7364
rect 10376 7392 10382 7404
rect 10873 7395 10931 7401
rect 10873 7392 10885 7395
rect 10376 7364 10885 7392
rect 10376 7352 10382 7364
rect 10873 7361 10885 7364
rect 10919 7392 10931 7395
rect 11790 7392 11796 7404
rect 10919 7364 11796 7392
rect 10919 7361 10931 7364
rect 10873 7355 10931 7361
rect 11790 7352 11796 7364
rect 11848 7352 11854 7404
rect 16298 7352 16304 7404
rect 16356 7392 16362 7404
rect 25409 7395 25467 7401
rect 25409 7392 25421 7395
rect 16356 7364 25421 7392
rect 16356 7352 16362 7364
rect 25409 7361 25421 7364
rect 25455 7361 25467 7395
rect 25409 7355 25467 7361
rect 27154 7352 27160 7404
rect 27212 7352 27218 7404
rect 7745 7327 7803 7333
rect 7745 7293 7757 7327
rect 7791 7293 7803 7327
rect 7745 7287 7803 7293
rect 6604 7228 7420 7256
rect 7760 7256 7788 7287
rect 8754 7284 8760 7336
rect 8812 7284 8818 7336
rect 8941 7327 8999 7333
rect 8941 7293 8953 7327
rect 8987 7324 8999 7327
rect 9030 7324 9036 7336
rect 8987 7296 9036 7324
rect 8987 7293 8999 7296
rect 8941 7287 8999 7293
rect 9030 7284 9036 7296
rect 9088 7324 9094 7336
rect 9766 7324 9772 7336
rect 9088 7296 9772 7324
rect 9088 7284 9094 7296
rect 9766 7284 9772 7296
rect 9824 7284 9830 7336
rect 28350 7284 28356 7336
rect 28408 7284 28414 7336
rect 10502 7256 10508 7268
rect 7760 7228 10508 7256
rect 6604 7216 6610 7228
rect 10502 7216 10508 7228
rect 10560 7216 10566 7268
rect 8662 7188 8668 7200
rect 6288 7160 8668 7188
rect 5491 7157 5503 7160
rect 5445 7151 5503 7157
rect 8662 7148 8668 7160
rect 8720 7148 8726 7200
rect 9306 7148 9312 7200
rect 9364 7148 9370 7200
rect 10778 7148 10784 7200
rect 10836 7188 10842 7200
rect 11146 7188 11152 7200
rect 10836 7160 11152 7188
rect 10836 7148 10842 7160
rect 11146 7148 11152 7160
rect 11204 7148 11210 7200
rect 1104 7098 28888 7120
rect 1104 7046 4423 7098
rect 4475 7046 4487 7098
rect 4539 7046 4551 7098
rect 4603 7046 4615 7098
rect 4667 7046 4679 7098
rect 4731 7046 11369 7098
rect 11421 7046 11433 7098
rect 11485 7046 11497 7098
rect 11549 7046 11561 7098
rect 11613 7046 11625 7098
rect 11677 7046 18315 7098
rect 18367 7046 18379 7098
rect 18431 7046 18443 7098
rect 18495 7046 18507 7098
rect 18559 7046 18571 7098
rect 18623 7046 25261 7098
rect 25313 7046 25325 7098
rect 25377 7046 25389 7098
rect 25441 7046 25453 7098
rect 25505 7046 25517 7098
rect 25569 7046 28888 7098
rect 1104 7024 28888 7046
rect 7834 6944 7840 6996
rect 7892 6984 7898 6996
rect 7892 6956 9260 6984
rect 7892 6944 7898 6956
rect 3234 6876 3240 6928
rect 3292 6916 3298 6928
rect 3602 6916 3608 6928
rect 3292 6888 3608 6916
rect 3292 6876 3298 6888
rect 3602 6876 3608 6888
rect 3660 6876 3666 6928
rect 9232 6916 9260 6956
rect 9306 6944 9312 6996
rect 9364 6984 9370 6996
rect 9364 6956 12434 6984
rect 9364 6944 9370 6956
rect 11974 6916 11980 6928
rect 7116 6888 9076 6916
rect 9232 6888 11980 6916
rect 1118 6808 1124 6860
rect 1176 6848 1182 6860
rect 1489 6851 1547 6857
rect 1489 6848 1501 6851
rect 1176 6820 1501 6848
rect 1176 6808 1182 6820
rect 1489 6817 1501 6820
rect 1535 6817 1547 6851
rect 3881 6851 3939 6857
rect 3881 6848 3893 6851
rect 1489 6811 1547 6817
rect 1596 6820 3893 6848
rect 290 6740 296 6792
rect 348 6780 354 6792
rect 1596 6780 1624 6820
rect 3881 6817 3893 6820
rect 3927 6817 3939 6851
rect 3881 6811 3939 6817
rect 4890 6808 4896 6860
rect 4948 6848 4954 6860
rect 4985 6851 5043 6857
rect 4985 6848 4997 6851
rect 4948 6820 4997 6848
rect 4948 6808 4954 6820
rect 4985 6817 4997 6820
rect 5031 6817 5043 6851
rect 4985 6811 5043 6817
rect 5074 6808 5080 6860
rect 5132 6848 5138 6860
rect 5132 6820 6776 6848
rect 5132 6808 5138 6820
rect 348 6752 1624 6780
rect 1673 6783 1731 6789
rect 348 6740 354 6752
rect 1673 6749 1685 6783
rect 1719 6780 1731 6783
rect 1949 6783 2007 6789
rect 1949 6780 1961 6783
rect 1719 6752 1961 6780
rect 1719 6749 1731 6752
rect 1673 6743 1731 6749
rect 1949 6749 1961 6752
rect 1995 6749 2007 6783
rect 1949 6743 2007 6749
rect 2498 6740 2504 6792
rect 2556 6740 2562 6792
rect 2685 6783 2743 6789
rect 2685 6749 2697 6783
rect 2731 6749 2743 6783
rect 2685 6743 2743 6749
rect 1302 6672 1308 6724
rect 1360 6712 1366 6724
rect 2700 6712 2728 6743
rect 2866 6740 2872 6792
rect 2924 6780 2930 6792
rect 2961 6783 3019 6789
rect 2961 6780 2973 6783
rect 2924 6752 2973 6780
rect 2924 6740 2930 6752
rect 2961 6749 2973 6752
rect 3007 6749 3019 6783
rect 2961 6743 3019 6749
rect 3605 6783 3663 6789
rect 3605 6749 3617 6783
rect 3651 6780 3663 6783
rect 3786 6780 3792 6792
rect 3651 6752 3792 6780
rect 3651 6749 3663 6752
rect 3605 6743 3663 6749
rect 3786 6740 3792 6752
rect 3844 6740 3850 6792
rect 4065 6783 4123 6789
rect 4065 6749 4077 6783
rect 4111 6749 4123 6783
rect 4341 6783 4399 6789
rect 4341 6780 4353 6783
rect 4065 6743 4123 6749
rect 4172 6752 4353 6780
rect 1360 6684 2728 6712
rect 1360 6672 1366 6684
rect 3510 6672 3516 6724
rect 3568 6712 3574 6724
rect 4080 6712 4108 6743
rect 3568 6684 4108 6712
rect 3568 6672 3574 6684
rect 1854 6604 1860 6656
rect 1912 6604 1918 6656
rect 2869 6647 2927 6653
rect 2869 6613 2881 6647
rect 2915 6644 2927 6647
rect 3878 6644 3884 6656
rect 2915 6616 3884 6644
rect 2915 6613 2927 6616
rect 2869 6607 2927 6613
rect 3878 6604 3884 6616
rect 3936 6604 3942 6656
rect 4172 6644 4200 6752
rect 4341 6749 4353 6752
rect 4387 6749 4399 6783
rect 4341 6743 4399 6749
rect 6454 6740 6460 6792
rect 6512 6740 6518 6792
rect 6748 6724 6776 6820
rect 6822 6808 6828 6860
rect 6880 6848 6886 6860
rect 7116 6857 7144 6888
rect 9048 6860 9076 6888
rect 11974 6876 11980 6888
rect 12032 6876 12038 6928
rect 12406 6916 12434 6956
rect 24946 6916 24952 6928
rect 12406 6888 24952 6916
rect 24946 6876 24952 6888
rect 25004 6876 25010 6928
rect 7101 6851 7159 6857
rect 7101 6848 7113 6851
rect 6880 6820 7113 6848
rect 6880 6808 6886 6820
rect 7101 6817 7113 6820
rect 7147 6817 7159 6851
rect 8481 6851 8539 6857
rect 8481 6848 8493 6851
rect 7101 6811 7159 6817
rect 7208 6820 8493 6848
rect 7208 6780 7236 6820
rect 8481 6817 8493 6820
rect 8527 6817 8539 6851
rect 8481 6811 8539 6817
rect 8662 6808 8668 6860
rect 8720 6808 8726 6860
rect 9030 6808 9036 6860
rect 9088 6808 9094 6860
rect 9582 6808 9588 6860
rect 9640 6808 9646 6860
rect 9677 6851 9735 6857
rect 9677 6817 9689 6851
rect 9723 6848 9735 6851
rect 9766 6848 9772 6860
rect 9723 6820 9772 6848
rect 9723 6817 9735 6820
rect 9677 6811 9735 6817
rect 7116 6752 7236 6780
rect 7377 6783 7435 6789
rect 4249 6715 4307 6721
rect 4249 6681 4261 6715
rect 4295 6712 4307 6715
rect 4295 6684 5304 6712
rect 4295 6681 4307 6684
rect 4249 6675 4307 6681
rect 4890 6644 4896 6656
rect 4172 6616 4896 6644
rect 4890 6604 4896 6616
rect 4948 6604 4954 6656
rect 5276 6644 5304 6684
rect 5350 6672 5356 6724
rect 5408 6672 5414 6724
rect 6730 6672 6736 6724
rect 6788 6672 6794 6724
rect 7116 6644 7144 6752
rect 7377 6749 7389 6783
rect 7423 6780 7435 6783
rect 8018 6780 8024 6792
rect 7423 6752 8024 6780
rect 7423 6749 7435 6752
rect 7377 6743 7435 6749
rect 8018 6740 8024 6752
rect 8076 6740 8082 6792
rect 8110 6740 8116 6792
rect 8168 6780 8174 6792
rect 8941 6783 8999 6789
rect 8941 6780 8953 6783
rect 8168 6752 8953 6780
rect 8168 6740 8174 6752
rect 8941 6749 8953 6752
rect 8987 6749 8999 6783
rect 8941 6743 8999 6749
rect 8389 6715 8447 6721
rect 8389 6681 8401 6715
rect 8435 6712 8447 6715
rect 9692 6712 9720 6811
rect 9766 6808 9772 6820
rect 9824 6848 9830 6860
rect 9824 6820 27200 6848
rect 9824 6808 9830 6820
rect 27172 6789 27200 6820
rect 9861 6783 9919 6789
rect 9861 6749 9873 6783
rect 9907 6749 9919 6783
rect 9861 6743 9919 6749
rect 10045 6783 10103 6789
rect 10045 6749 10057 6783
rect 10091 6780 10103 6783
rect 25685 6783 25743 6789
rect 25685 6780 25697 6783
rect 10091 6752 12434 6780
rect 10091 6749 10103 6752
rect 10045 6743 10103 6749
rect 8435 6684 9720 6712
rect 8435 6681 8447 6684
rect 8389 6675 8447 6681
rect 5276 6616 7144 6644
rect 7650 6604 7656 6656
rect 7708 6644 7714 6656
rect 7929 6647 7987 6653
rect 7929 6644 7941 6647
rect 7708 6616 7941 6644
rect 7708 6604 7714 6616
rect 7929 6613 7941 6616
rect 7975 6613 7987 6647
rect 7929 6607 7987 6613
rect 8018 6604 8024 6656
rect 8076 6604 8082 6656
rect 8478 6604 8484 6656
rect 8536 6644 8542 6656
rect 9876 6644 9904 6743
rect 10318 6672 10324 6724
rect 10376 6672 10382 6724
rect 8536 6616 9904 6644
rect 8536 6604 8542 6616
rect 10778 6604 10784 6656
rect 10836 6604 10842 6656
rect 12406 6644 12434 6752
rect 25516 6752 25697 6780
rect 12618 6672 12624 6724
rect 12676 6712 12682 6724
rect 25516 6721 25544 6752
rect 25685 6749 25697 6752
rect 25731 6749 25743 6783
rect 25685 6743 25743 6749
rect 27157 6783 27215 6789
rect 27157 6749 27169 6783
rect 27203 6749 27215 6783
rect 27157 6743 27215 6749
rect 25501 6715 25559 6721
rect 25501 6712 25513 6715
rect 12676 6684 25513 6712
rect 12676 6672 12682 6684
rect 25501 6681 25513 6684
rect 25547 6681 25559 6715
rect 25501 6675 25559 6681
rect 26878 6672 26884 6724
rect 26936 6672 26942 6724
rect 28350 6672 28356 6724
rect 28408 6672 28414 6724
rect 22370 6644 22376 6656
rect 12406 6616 22376 6644
rect 22370 6604 22376 6616
rect 22428 6604 22434 6656
rect 1104 6554 29048 6576
rect 1104 6502 7896 6554
rect 7948 6502 7960 6554
rect 8012 6502 8024 6554
rect 8076 6502 8088 6554
rect 8140 6502 8152 6554
rect 8204 6502 14842 6554
rect 14894 6502 14906 6554
rect 14958 6502 14970 6554
rect 15022 6502 15034 6554
rect 15086 6502 15098 6554
rect 15150 6502 21788 6554
rect 21840 6502 21852 6554
rect 21904 6502 21916 6554
rect 21968 6502 21980 6554
rect 22032 6502 22044 6554
rect 22096 6502 28734 6554
rect 28786 6502 28798 6554
rect 28850 6502 28862 6554
rect 28914 6502 28926 6554
rect 28978 6502 28990 6554
rect 29042 6502 29048 6554
rect 1104 6480 29048 6502
rect 2041 6443 2099 6449
rect 2041 6409 2053 6443
rect 2087 6440 2099 6443
rect 2222 6440 2228 6452
rect 2087 6412 2228 6440
rect 2087 6409 2099 6412
rect 2041 6403 2099 6409
rect 2222 6400 2228 6412
rect 2280 6400 2286 6452
rect 3878 6400 3884 6452
rect 3936 6400 3942 6452
rect 4338 6400 4344 6452
rect 4396 6440 4402 6452
rect 4617 6443 4675 6449
rect 4617 6440 4629 6443
rect 4396 6412 4629 6440
rect 4396 6400 4402 6412
rect 4617 6409 4629 6412
rect 4663 6409 4675 6443
rect 4617 6403 4675 6409
rect 5350 6400 5356 6452
rect 5408 6400 5414 6452
rect 6362 6400 6368 6452
rect 6420 6400 6426 6452
rect 7374 6400 7380 6452
rect 7432 6400 7438 6452
rect 7650 6400 7656 6452
rect 7708 6400 7714 6452
rect 8294 6440 8300 6452
rect 7852 6412 8300 6440
rect 3896 6372 3924 6400
rect 7190 6372 7196 6384
rect 3896 6344 7196 6372
rect 7190 6332 7196 6344
rect 7248 6332 7254 6384
rect 3602 6304 3608 6316
rect 2746 6276 3608 6304
rect 1489 6239 1547 6245
rect 1489 6205 1501 6239
rect 1535 6205 1547 6239
rect 1489 6199 1547 6205
rect 1504 6168 1532 6199
rect 2222 6196 2228 6248
rect 2280 6196 2286 6248
rect 2746 6168 2774 6276
rect 3602 6264 3608 6276
rect 3660 6264 3666 6316
rect 4172 6276 5120 6304
rect 3053 6239 3111 6245
rect 3053 6205 3065 6239
rect 3099 6236 3111 6239
rect 3694 6236 3700 6248
rect 3099 6208 3700 6236
rect 3099 6205 3111 6208
rect 3053 6199 3111 6205
rect 3694 6196 3700 6208
rect 3752 6236 3758 6248
rect 4172 6236 4200 6276
rect 5092 6248 5120 6276
rect 5902 6264 5908 6316
rect 5960 6264 5966 6316
rect 7101 6307 7159 6313
rect 7101 6304 7113 6307
rect 6932 6276 7113 6304
rect 3752 6208 4200 6236
rect 3752 6196 3758 6208
rect 4246 6196 4252 6248
rect 4304 6236 4310 6248
rect 4433 6239 4491 6245
rect 4433 6236 4445 6239
rect 4304 6208 4445 6236
rect 4304 6196 4310 6208
rect 4433 6205 4445 6208
rect 4479 6205 4491 6239
rect 4433 6199 4491 6205
rect 5074 6196 5080 6248
rect 5132 6196 5138 6248
rect 5261 6239 5319 6245
rect 5261 6205 5273 6239
rect 5307 6236 5319 6239
rect 6638 6236 6644 6248
rect 5307 6208 6644 6236
rect 5307 6205 5319 6208
rect 5261 6199 5319 6205
rect 6638 6196 6644 6208
rect 6696 6196 6702 6248
rect 1504 6140 2774 6168
rect 3605 6171 3663 6177
rect 3605 6137 3617 6171
rect 3651 6168 3663 6171
rect 4338 6168 4344 6180
rect 3651 6140 4344 6168
rect 3651 6137 3663 6140
rect 3605 6131 3663 6137
rect 4338 6128 4344 6140
rect 4396 6128 4402 6180
rect 2774 6060 2780 6112
rect 2832 6060 2838 6112
rect 3878 6060 3884 6112
rect 3936 6060 3942 6112
rect 5902 6060 5908 6112
rect 5960 6100 5966 6112
rect 6932 6100 6960 6276
rect 7101 6273 7113 6276
rect 7147 6273 7159 6307
rect 7101 6267 7159 6273
rect 7285 6307 7343 6313
rect 7285 6273 7297 6307
rect 7331 6304 7343 6307
rect 7392 6304 7420 6400
rect 7331 6276 7420 6304
rect 7331 6273 7343 6276
rect 7285 6267 7343 6273
rect 7009 6239 7067 6245
rect 7009 6205 7021 6239
rect 7055 6205 7067 6239
rect 7668 6236 7696 6400
rect 7852 6372 7880 6412
rect 8294 6400 8300 6412
rect 8352 6440 8358 6452
rect 8938 6440 8944 6452
rect 8352 6412 8944 6440
rect 8352 6400 8358 6412
rect 8938 6400 8944 6412
rect 8996 6400 9002 6452
rect 9766 6400 9772 6452
rect 9824 6400 9830 6452
rect 9858 6400 9864 6452
rect 9916 6440 9922 6452
rect 10137 6443 10195 6449
rect 10137 6440 10149 6443
rect 9916 6412 10149 6440
rect 9916 6400 9922 6412
rect 10137 6409 10149 6412
rect 10183 6440 10195 6443
rect 10318 6440 10324 6452
rect 10183 6412 10324 6440
rect 10183 6409 10195 6412
rect 10137 6403 10195 6409
rect 10318 6400 10324 6412
rect 10376 6400 10382 6452
rect 10888 6412 25452 6440
rect 7760 6344 7880 6372
rect 7760 6313 7788 6344
rect 9030 6332 9036 6384
rect 9088 6332 9094 6384
rect 9784 6313 9812 6400
rect 7745 6307 7803 6313
rect 7745 6273 7757 6307
rect 7791 6273 7803 6307
rect 7745 6267 7803 6273
rect 9769 6307 9827 6313
rect 9769 6273 9781 6307
rect 9815 6273 9827 6307
rect 9769 6267 9827 6273
rect 8021 6239 8079 6245
rect 8021 6236 8033 6239
rect 7668 6208 8033 6236
rect 7009 6199 7067 6205
rect 8021 6205 8033 6208
rect 8067 6205 8079 6239
rect 8021 6199 8079 6205
rect 7024 6168 7052 6199
rect 9214 6196 9220 6248
rect 9272 6236 9278 6248
rect 10888 6236 10916 6412
rect 23750 6264 23756 6316
rect 23808 6304 23814 6316
rect 23937 6307 23995 6313
rect 23937 6304 23949 6307
rect 23808 6276 23949 6304
rect 23808 6264 23814 6276
rect 23937 6273 23949 6276
rect 23983 6273 23995 6307
rect 23937 6267 23995 6273
rect 24578 6264 24584 6316
rect 24636 6304 24642 6316
rect 25424 6313 25452 6412
rect 25409 6307 25467 6313
rect 24636 6276 24854 6304
rect 24636 6264 24642 6276
rect 9272 6208 10916 6236
rect 9272 6196 9278 6208
rect 24670 6196 24676 6248
rect 24728 6196 24734 6248
rect 24826 6236 24854 6276
rect 25409 6273 25421 6307
rect 25455 6273 25467 6307
rect 27157 6307 27215 6313
rect 27157 6304 27169 6307
rect 25409 6267 25467 6273
rect 25516 6276 27169 6304
rect 25516 6236 25544 6276
rect 27157 6273 27169 6276
rect 27203 6273 27215 6307
rect 27157 6267 27215 6273
rect 24826 6208 25544 6236
rect 26142 6196 26148 6248
rect 26200 6196 26206 6248
rect 28353 6239 28411 6245
rect 28353 6205 28365 6239
rect 28399 6236 28411 6239
rect 28626 6236 28632 6248
rect 28399 6208 28632 6236
rect 28399 6205 28411 6208
rect 28353 6199 28411 6205
rect 28626 6196 28632 6208
rect 28684 6196 28690 6248
rect 7024 6140 7880 6168
rect 5960 6072 6960 6100
rect 5960 6060 5966 6072
rect 7466 6060 7472 6112
rect 7524 6060 7530 6112
rect 7852 6100 7880 6140
rect 9490 6128 9496 6180
rect 9548 6168 9554 6180
rect 24854 6168 24860 6180
rect 9548 6140 24860 6168
rect 9548 6128 9554 6140
rect 24854 6128 24860 6140
rect 24912 6128 24918 6180
rect 8570 6100 8576 6112
rect 7852 6072 8576 6100
rect 8570 6060 8576 6072
rect 8628 6060 8634 6112
rect 10226 6060 10232 6112
rect 10284 6100 10290 6112
rect 10505 6103 10563 6109
rect 10505 6100 10517 6103
rect 10284 6072 10517 6100
rect 10284 6060 10290 6072
rect 10505 6069 10517 6072
rect 10551 6100 10563 6103
rect 17218 6100 17224 6112
rect 10551 6072 17224 6100
rect 10551 6069 10563 6072
rect 10505 6063 10563 6069
rect 17218 6060 17224 6072
rect 17276 6060 17282 6112
rect 23750 6060 23756 6112
rect 23808 6060 23814 6112
rect 1104 6010 28888 6032
rect 1104 5958 4423 6010
rect 4475 5958 4487 6010
rect 4539 5958 4551 6010
rect 4603 5958 4615 6010
rect 4667 5958 4679 6010
rect 4731 5958 11369 6010
rect 11421 5958 11433 6010
rect 11485 5958 11497 6010
rect 11549 5958 11561 6010
rect 11613 5958 11625 6010
rect 11677 5958 18315 6010
rect 18367 5958 18379 6010
rect 18431 5958 18443 6010
rect 18495 5958 18507 6010
rect 18559 5958 18571 6010
rect 18623 5958 25261 6010
rect 25313 5958 25325 6010
rect 25377 5958 25389 6010
rect 25441 5958 25453 6010
rect 25505 5958 25517 6010
rect 25569 5958 28888 6010
rect 1104 5936 28888 5958
rect 2777 5899 2835 5905
rect 2777 5865 2789 5899
rect 2823 5896 2835 5899
rect 2958 5896 2964 5908
rect 2823 5868 2964 5896
rect 2823 5865 2835 5868
rect 2777 5859 2835 5865
rect 2958 5856 2964 5868
rect 3016 5856 3022 5908
rect 3418 5856 3424 5908
rect 3476 5896 3482 5908
rect 3513 5899 3571 5905
rect 3513 5896 3525 5899
rect 3476 5868 3525 5896
rect 3476 5856 3482 5868
rect 3513 5865 3525 5868
rect 3559 5865 3571 5899
rect 3513 5859 3571 5865
rect 3878 5856 3884 5908
rect 3936 5896 3942 5908
rect 4230 5899 4288 5905
rect 4230 5896 4242 5899
rect 3936 5868 4242 5896
rect 3936 5856 3942 5868
rect 4230 5865 4242 5868
rect 4276 5865 4288 5899
rect 4230 5859 4288 5865
rect 6730 5856 6736 5908
rect 6788 5896 6794 5908
rect 7561 5899 7619 5905
rect 7561 5896 7573 5899
rect 6788 5868 7573 5896
rect 6788 5856 6794 5868
rect 7561 5865 7573 5868
rect 7607 5896 7619 5899
rect 8294 5896 8300 5908
rect 7607 5868 8300 5896
rect 7607 5865 7619 5868
rect 7561 5859 7619 5865
rect 8294 5856 8300 5868
rect 8352 5856 8358 5908
rect 8386 5856 8392 5908
rect 8444 5896 8450 5908
rect 8665 5899 8723 5905
rect 8665 5896 8677 5899
rect 8444 5868 8677 5896
rect 8444 5856 8450 5868
rect 8665 5865 8677 5868
rect 8711 5865 8723 5899
rect 8665 5859 8723 5865
rect 9030 5856 9036 5908
rect 9088 5856 9094 5908
rect 9122 5856 9128 5908
rect 9180 5896 9186 5908
rect 9401 5899 9459 5905
rect 9401 5896 9413 5899
rect 9180 5868 9413 5896
rect 9180 5856 9186 5868
rect 9401 5865 9413 5868
rect 9447 5865 9459 5899
rect 9401 5859 9459 5865
rect 9858 5856 9864 5908
rect 9916 5856 9922 5908
rect 10226 5856 10232 5908
rect 10284 5856 10290 5908
rect 17218 5856 17224 5908
rect 17276 5896 17282 5908
rect 26694 5896 26700 5908
rect 17276 5868 26700 5896
rect 17276 5856 17282 5868
rect 26694 5856 26700 5868
rect 26752 5856 26758 5908
rect 2041 5831 2099 5837
rect 2041 5797 2053 5831
rect 2087 5828 2099 5831
rect 3326 5828 3332 5840
rect 2087 5800 3332 5828
rect 2087 5797 2099 5800
rect 2041 5791 2099 5797
rect 3326 5788 3332 5800
rect 3384 5788 3390 5840
rect 6638 5788 6644 5840
rect 6696 5828 6702 5840
rect 7834 5828 7840 5840
rect 6696 5800 7840 5828
rect 6696 5788 6702 5800
rect 7834 5788 7840 5800
rect 7892 5788 7898 5840
rect 7926 5788 7932 5840
rect 7984 5788 7990 5840
rect 8018 5788 8024 5840
rect 8076 5828 8082 5840
rect 11698 5828 11704 5840
rect 8076 5800 11704 5828
rect 8076 5788 8082 5800
rect 11698 5788 11704 5800
rect 11756 5788 11762 5840
rect 2590 5720 2596 5772
rect 2648 5760 2654 5772
rect 2869 5763 2927 5769
rect 2869 5760 2881 5763
rect 2648 5732 2881 5760
rect 2648 5720 2654 5732
rect 2869 5729 2881 5732
rect 2915 5729 2927 5763
rect 2869 5723 2927 5729
rect 3694 5720 3700 5772
rect 3752 5760 3758 5772
rect 3973 5763 4031 5769
rect 3973 5760 3985 5763
rect 3752 5732 3985 5760
rect 3752 5720 3758 5732
rect 3973 5729 3985 5732
rect 4019 5760 4031 5763
rect 5994 5760 6000 5772
rect 4019 5732 6000 5760
rect 4019 5729 4031 5732
rect 3973 5723 4031 5729
rect 5994 5720 6000 5732
rect 6052 5720 6058 5772
rect 10226 5760 10232 5772
rect 6564 5732 10232 5760
rect 1489 5695 1547 5701
rect 1489 5661 1501 5695
rect 1535 5692 1547 5695
rect 1762 5692 1768 5704
rect 1535 5664 1768 5692
rect 1535 5661 1547 5664
rect 1489 5655 1547 5661
rect 1762 5652 1768 5664
rect 1820 5652 1826 5704
rect 2225 5695 2283 5701
rect 2225 5661 2237 5695
rect 2271 5692 2283 5695
rect 6564 5692 6592 5732
rect 10226 5720 10232 5732
rect 10284 5720 10290 5772
rect 13998 5720 14004 5772
rect 14056 5760 14062 5772
rect 14056 5732 24854 5760
rect 14056 5720 14062 5732
rect 2271 5664 2774 5692
rect 2271 5661 2283 5664
rect 2225 5655 2283 5661
rect 2746 5556 2774 5664
rect 6012 5664 6592 5692
rect 6012 5636 6040 5664
rect 7466 5652 7472 5704
rect 7524 5652 7530 5704
rect 7558 5652 7564 5704
rect 7616 5692 7622 5704
rect 8113 5695 8171 5701
rect 8113 5692 8125 5695
rect 7616 5664 8125 5692
rect 7616 5652 7622 5664
rect 8113 5661 8125 5664
rect 8159 5661 8171 5695
rect 8113 5655 8171 5661
rect 8389 5695 8447 5701
rect 8389 5661 8401 5695
rect 8435 5692 8447 5695
rect 8662 5692 8668 5704
rect 8435 5664 8668 5692
rect 8435 5661 8447 5664
rect 8389 5655 8447 5661
rect 8662 5652 8668 5664
rect 8720 5652 8726 5704
rect 9125 5695 9183 5701
rect 9125 5661 9137 5695
rect 9171 5692 9183 5695
rect 9858 5692 9864 5704
rect 9171 5664 9864 5692
rect 9171 5661 9183 5664
rect 9125 5655 9183 5661
rect 9858 5652 9864 5664
rect 9916 5652 9922 5704
rect 22830 5652 22836 5704
rect 22888 5652 22894 5704
rect 24826 5692 24854 5732
rect 26418 5720 26424 5772
rect 26476 5720 26482 5772
rect 25685 5695 25743 5701
rect 25685 5692 25697 5695
rect 24826 5664 25697 5692
rect 25685 5661 25697 5664
rect 25731 5661 25743 5695
rect 26712 5692 26740 5856
rect 28353 5763 28411 5769
rect 28353 5729 28365 5763
rect 28399 5760 28411 5763
rect 28810 5760 28816 5772
rect 28399 5732 28816 5760
rect 28399 5729 28411 5732
rect 28353 5723 28411 5729
rect 28810 5720 28816 5732
rect 28868 5720 28874 5772
rect 27157 5695 27215 5701
rect 27157 5692 27169 5695
rect 26712 5664 27169 5692
rect 25685 5655 25743 5661
rect 27157 5661 27169 5664
rect 27203 5661 27215 5695
rect 27157 5655 27215 5661
rect 4798 5584 4804 5636
rect 4856 5584 4862 5636
rect 5994 5584 6000 5636
rect 6052 5584 6058 5636
rect 6086 5584 6092 5636
rect 6144 5624 6150 5636
rect 7098 5624 7104 5636
rect 6144 5596 7104 5624
rect 6144 5584 6150 5596
rect 7098 5584 7104 5596
rect 7156 5584 7162 5636
rect 7484 5624 7512 5652
rect 24029 5627 24087 5633
rect 7484 5596 12434 5624
rect 4430 5556 4436 5568
rect 2746 5528 4436 5556
rect 4430 5516 4436 5528
rect 4488 5516 4494 5568
rect 5810 5516 5816 5568
rect 5868 5556 5874 5568
rect 8205 5559 8263 5565
rect 8205 5556 8217 5559
rect 5868 5528 8217 5556
rect 5868 5516 5874 5528
rect 8205 5525 8217 5528
rect 8251 5525 8263 5559
rect 8205 5519 8263 5525
rect 9674 5516 9680 5568
rect 9732 5556 9738 5568
rect 11790 5556 11796 5568
rect 9732 5528 11796 5556
rect 9732 5516 9738 5528
rect 11790 5516 11796 5528
rect 11848 5516 11854 5568
rect 12406 5556 12434 5596
rect 24029 5593 24041 5627
rect 24075 5624 24087 5627
rect 27246 5624 27252 5636
rect 24075 5596 27252 5624
rect 24075 5593 24087 5596
rect 24029 5587 24087 5593
rect 27246 5584 27252 5596
rect 27304 5584 27310 5636
rect 13078 5556 13084 5568
rect 12406 5528 13084 5556
rect 13078 5516 13084 5528
rect 13136 5516 13142 5568
rect 1104 5466 29048 5488
rect 1104 5414 7896 5466
rect 7948 5414 7960 5466
rect 8012 5414 8024 5466
rect 8076 5414 8088 5466
rect 8140 5414 8152 5466
rect 8204 5414 14842 5466
rect 14894 5414 14906 5466
rect 14958 5414 14970 5466
rect 15022 5414 15034 5466
rect 15086 5414 15098 5466
rect 15150 5414 21788 5466
rect 21840 5414 21852 5466
rect 21904 5414 21916 5466
rect 21968 5414 21980 5466
rect 22032 5414 22044 5466
rect 22096 5414 28734 5466
rect 28786 5414 28798 5466
rect 28850 5414 28862 5466
rect 28914 5414 28926 5466
rect 28978 5414 28990 5466
rect 29042 5414 29048 5466
rect 1104 5392 29048 5414
rect 658 5312 664 5364
rect 716 5312 722 5364
rect 3050 5312 3056 5364
rect 3108 5352 3114 5364
rect 3694 5352 3700 5364
rect 3108 5324 3700 5352
rect 3108 5312 3114 5324
rect 3694 5312 3700 5324
rect 3752 5312 3758 5364
rect 4246 5312 4252 5364
rect 4304 5352 4310 5364
rect 4433 5355 4491 5361
rect 4433 5352 4445 5355
rect 4304 5324 4445 5352
rect 4304 5312 4310 5324
rect 4433 5321 4445 5324
rect 4479 5321 4491 5355
rect 4433 5315 4491 5321
rect 5442 5312 5448 5364
rect 5500 5312 5506 5364
rect 6086 5352 6092 5364
rect 5552 5324 6092 5352
rect 676 5284 704 5312
rect 3326 5284 3332 5296
rect 676 5256 3332 5284
rect 3326 5244 3332 5256
rect 3384 5244 3390 5296
rect 4341 5287 4399 5293
rect 4341 5253 4353 5287
rect 4387 5284 4399 5287
rect 5552 5284 5580 5324
rect 6086 5312 6092 5324
rect 6144 5312 6150 5364
rect 6454 5312 6460 5364
rect 6512 5312 6518 5364
rect 8478 5352 8484 5364
rect 8266 5324 8484 5352
rect 5994 5284 6000 5296
rect 4387 5256 5580 5284
rect 5644 5256 6000 5284
rect 4387 5253 4399 5256
rect 4341 5247 4399 5253
rect 382 5176 388 5228
rect 440 5216 446 5228
rect 1397 5219 1455 5225
rect 1397 5216 1409 5219
rect 440 5188 1409 5216
rect 440 5176 446 5188
rect 1397 5185 1409 5188
rect 1443 5185 1455 5219
rect 1397 5179 1455 5185
rect 1578 5176 1584 5228
rect 1636 5176 1642 5228
rect 2130 5176 2136 5228
rect 2188 5216 2194 5228
rect 3970 5216 3976 5228
rect 2188 5188 3976 5216
rect 2188 5176 2194 5188
rect 3970 5176 3976 5188
rect 4028 5176 4034 5228
rect 4801 5219 4859 5225
rect 4801 5185 4813 5219
rect 4847 5216 4859 5219
rect 5644 5216 5672 5256
rect 5994 5244 6000 5256
rect 6052 5244 6058 5296
rect 7742 5244 7748 5296
rect 7800 5244 7806 5296
rect 8266 5284 8294 5324
rect 8478 5312 8484 5324
rect 8536 5312 8542 5364
rect 8665 5355 8723 5361
rect 8665 5321 8677 5355
rect 8711 5352 8723 5355
rect 8754 5352 8760 5364
rect 8711 5324 8760 5352
rect 8711 5321 8723 5324
rect 8665 5315 8723 5321
rect 8754 5312 8760 5324
rect 8812 5312 8818 5364
rect 9030 5312 9036 5364
rect 9088 5352 9094 5364
rect 24578 5352 24584 5364
rect 9088 5324 24584 5352
rect 9088 5312 9094 5324
rect 24578 5312 24584 5324
rect 24636 5312 24642 5364
rect 26694 5312 26700 5364
rect 26752 5312 26758 5364
rect 9858 5284 9864 5296
rect 8128 5256 8294 5284
rect 9508 5256 9864 5284
rect 6546 5216 6552 5228
rect 4847 5188 5672 5216
rect 5828 5188 6552 5216
rect 4847 5185 4859 5188
rect 4801 5179 4859 5185
rect 1946 5108 1952 5160
rect 2004 5108 2010 5160
rect 4893 5151 4951 5157
rect 4893 5148 4905 5151
rect 2746 5120 4905 5148
rect 1765 5083 1823 5089
rect 1765 5049 1777 5083
rect 1811 5080 1823 5083
rect 2746 5080 2774 5120
rect 4893 5117 4905 5120
rect 4939 5117 4951 5151
rect 4893 5111 4951 5117
rect 4982 5108 4988 5160
rect 5040 5108 5046 5160
rect 5350 5108 5356 5160
rect 5408 5148 5414 5160
rect 5828 5148 5856 5188
rect 6546 5176 6552 5188
rect 6604 5176 6610 5228
rect 8128 5216 8156 5256
rect 8036 5188 8156 5216
rect 5408 5120 5856 5148
rect 5408 5108 5414 5120
rect 6086 5108 6092 5160
rect 6144 5108 6150 5160
rect 7285 5151 7343 5157
rect 7285 5117 7297 5151
rect 7331 5148 7343 5151
rect 7331 5120 7420 5148
rect 7331 5117 7343 5120
rect 7285 5111 7343 5117
rect 7392 5089 7420 5120
rect 7834 5108 7840 5160
rect 7892 5108 7898 5160
rect 8036 5157 8064 5188
rect 8248 5176 8254 5228
rect 8306 5216 8312 5228
rect 8306 5176 8340 5216
rect 8386 5176 8392 5228
rect 8444 5176 8450 5228
rect 8478 5176 8484 5228
rect 8536 5176 8542 5228
rect 8938 5176 8944 5228
rect 8996 5176 9002 5228
rect 9214 5176 9220 5228
rect 9272 5176 9278 5228
rect 9508 5225 9536 5256
rect 9858 5244 9864 5256
rect 9916 5284 9922 5296
rect 10505 5287 10563 5293
rect 10505 5284 10517 5287
rect 9916 5256 10517 5284
rect 9916 5244 9922 5256
rect 10505 5253 10517 5256
rect 10551 5253 10563 5287
rect 10505 5247 10563 5253
rect 14458 5244 14464 5296
rect 14516 5284 14522 5296
rect 14516 5256 27016 5284
rect 14516 5244 14522 5256
rect 9493 5219 9551 5225
rect 9493 5185 9505 5219
rect 9539 5185 9551 5219
rect 9493 5179 9551 5185
rect 17402 5176 17408 5228
rect 17460 5216 17466 5228
rect 21913 5219 21971 5225
rect 21913 5216 21925 5219
rect 17460 5188 21925 5216
rect 17460 5176 17466 5188
rect 21913 5185 21925 5188
rect 21959 5185 21971 5219
rect 21913 5179 21971 5185
rect 23474 5176 23480 5228
rect 23532 5176 23538 5228
rect 24854 5176 24860 5228
rect 24912 5176 24918 5228
rect 26988 5225 27016 5256
rect 26973 5219 27031 5225
rect 26973 5185 26985 5219
rect 27019 5185 27031 5219
rect 26973 5179 27031 5185
rect 8021 5151 8079 5157
rect 8021 5117 8033 5151
rect 8067 5117 8079 5151
rect 8312 5148 8340 5176
rect 10962 5148 10968 5160
rect 8312 5120 10968 5148
rect 8021 5111 8079 5117
rect 10962 5108 10968 5120
rect 11020 5108 11026 5160
rect 23109 5151 23167 5157
rect 23109 5117 23121 5151
rect 23155 5117 23167 5151
rect 23109 5111 23167 5117
rect 24581 5151 24639 5157
rect 24581 5117 24593 5151
rect 24627 5117 24639 5151
rect 24581 5111 24639 5117
rect 1811 5052 2774 5080
rect 7377 5083 7435 5089
rect 1811 5049 1823 5052
rect 1765 5043 1823 5049
rect 7377 5049 7389 5083
rect 7423 5049 7435 5083
rect 7377 5043 7435 5049
rect 8110 5040 8116 5092
rect 8168 5080 8174 5092
rect 9033 5083 9091 5089
rect 9033 5080 9045 5083
rect 8168 5052 9045 5080
rect 8168 5040 8174 5052
rect 9033 5049 9045 5052
rect 9079 5049 9091 5083
rect 9033 5043 9091 5049
rect 2498 4972 2504 5024
rect 2556 4972 2562 5024
rect 2682 4972 2688 5024
rect 2740 5012 2746 5024
rect 4890 5012 4896 5024
rect 2740 4984 4896 5012
rect 2740 4972 2746 4984
rect 4890 4972 4896 4984
rect 4948 4972 4954 5024
rect 6638 4972 6644 5024
rect 6696 4972 6702 5024
rect 8202 4972 8208 5024
rect 8260 4972 8266 5024
rect 8570 4972 8576 5024
rect 8628 5012 8634 5024
rect 8757 5015 8815 5021
rect 8757 5012 8769 5015
rect 8628 4984 8769 5012
rect 8628 4972 8634 4984
rect 8757 4981 8769 4984
rect 8803 4981 8815 5015
rect 8757 4975 8815 4981
rect 8846 4972 8852 5024
rect 8904 5012 8910 5024
rect 9401 5015 9459 5021
rect 9401 5012 9413 5015
rect 8904 4984 9413 5012
rect 8904 4972 8910 4984
rect 9401 4981 9413 4984
rect 9447 4981 9459 5015
rect 9401 4975 9459 4981
rect 10229 5015 10287 5021
rect 10229 4981 10241 5015
rect 10275 5012 10287 5015
rect 10778 5012 10784 5024
rect 10275 4984 10784 5012
rect 10275 4981 10287 4984
rect 10229 4975 10287 4981
rect 10778 4972 10784 4984
rect 10836 5012 10842 5024
rect 10965 5015 11023 5021
rect 10965 5012 10977 5015
rect 10836 4984 10977 5012
rect 10836 4972 10842 4984
rect 10965 4981 10977 4984
rect 11011 5012 11023 5015
rect 11146 5012 11152 5024
rect 11011 4984 11152 5012
rect 11011 4981 11023 4984
rect 10965 4975 11023 4981
rect 11146 4972 11152 4984
rect 11204 4972 11210 5024
rect 23124 5012 23152 5111
rect 24596 5080 24624 5111
rect 24762 5108 24768 5160
rect 24820 5148 24826 5160
rect 25317 5151 25375 5157
rect 25317 5148 25329 5151
rect 24820 5120 25329 5148
rect 24820 5108 24826 5120
rect 25317 5117 25329 5120
rect 25363 5117 25375 5151
rect 25317 5111 25375 5117
rect 25958 5108 25964 5160
rect 26016 5148 26022 5160
rect 27433 5151 27491 5157
rect 27433 5148 27445 5151
rect 26016 5120 27445 5148
rect 26016 5108 26022 5120
rect 27433 5117 27445 5120
rect 27479 5117 27491 5151
rect 27433 5111 27491 5117
rect 26510 5080 26516 5092
rect 24596 5052 26516 5080
rect 26510 5040 26516 5052
rect 26568 5040 26574 5092
rect 28074 5012 28080 5024
rect 23124 4984 28080 5012
rect 28074 4972 28080 4984
rect 28132 4972 28138 5024
rect 1104 4922 28888 4944
rect 1104 4870 4423 4922
rect 4475 4870 4487 4922
rect 4539 4870 4551 4922
rect 4603 4870 4615 4922
rect 4667 4870 4679 4922
rect 4731 4870 11369 4922
rect 11421 4870 11433 4922
rect 11485 4870 11497 4922
rect 11549 4870 11561 4922
rect 11613 4870 11625 4922
rect 11677 4870 18315 4922
rect 18367 4870 18379 4922
rect 18431 4870 18443 4922
rect 18495 4870 18507 4922
rect 18559 4870 18571 4922
rect 18623 4870 25261 4922
rect 25313 4870 25325 4922
rect 25377 4870 25389 4922
rect 25441 4870 25453 4922
rect 25505 4870 25517 4922
rect 25569 4870 28888 4922
rect 1104 4848 28888 4870
rect 2222 4768 2228 4820
rect 2280 4808 2286 4820
rect 3789 4811 3847 4817
rect 3789 4808 3801 4811
rect 2280 4780 3801 4808
rect 2280 4768 2286 4780
rect 3789 4777 3801 4780
rect 3835 4777 3847 4811
rect 3789 4771 3847 4777
rect 3970 4768 3976 4820
rect 4028 4768 4034 4820
rect 4062 4768 4068 4820
rect 4120 4768 4126 4820
rect 5077 4811 5135 4817
rect 5077 4777 5089 4811
rect 5123 4808 5135 4811
rect 5166 4808 5172 4820
rect 5123 4780 5172 4808
rect 5123 4777 5135 4780
rect 5077 4771 5135 4777
rect 5166 4768 5172 4780
rect 5224 4768 5230 4820
rect 5534 4768 5540 4820
rect 5592 4808 5598 4820
rect 5905 4811 5963 4817
rect 5905 4808 5917 4811
rect 5592 4780 5917 4808
rect 5592 4768 5598 4780
rect 5905 4777 5917 4780
rect 5951 4777 5963 4811
rect 5905 4771 5963 4777
rect 6840 4780 8984 4808
rect 2869 4743 2927 4749
rect 2869 4709 2881 4743
rect 2915 4740 2927 4743
rect 3510 4740 3516 4752
rect 2915 4712 3516 4740
rect 2915 4709 2927 4712
rect 2869 4703 2927 4709
rect 3510 4700 3516 4712
rect 3568 4700 3574 4752
rect 3605 4743 3663 4749
rect 3605 4709 3617 4743
rect 3651 4740 3663 4743
rect 4080 4740 4108 4768
rect 3651 4712 4108 4740
rect 3651 4709 3663 4712
rect 3605 4703 3663 4709
rect 4338 4700 4344 4752
rect 4396 4700 4402 4752
rect 6840 4740 6868 4780
rect 6564 4712 6868 4740
rect 1210 4632 1216 4684
rect 1268 4672 1274 4684
rect 1489 4675 1547 4681
rect 1489 4672 1501 4675
rect 1268 4644 1501 4672
rect 1268 4632 1274 4644
rect 1489 4641 1501 4644
rect 1535 4641 1547 4675
rect 1489 4635 1547 4641
rect 2746 4644 3924 4672
rect 1302 4564 1308 4616
rect 1360 4604 1366 4616
rect 2225 4607 2283 4613
rect 2225 4604 2237 4607
rect 1360 4576 2237 4604
rect 1360 4564 1366 4576
rect 2225 4573 2237 4576
rect 2271 4573 2283 4607
rect 2225 4567 2283 4573
rect 2133 4539 2191 4545
rect 2133 4505 2145 4539
rect 2179 4536 2191 4539
rect 2746 4536 2774 4644
rect 3896 4616 3924 4644
rect 3970 4632 3976 4684
rect 4028 4672 4034 4684
rect 5350 4672 5356 4684
rect 4028 4644 5356 4672
rect 4028 4632 4034 4644
rect 5350 4632 5356 4644
rect 5408 4632 5414 4684
rect 5810 4632 5816 4684
rect 5868 4632 5874 4684
rect 6564 4681 6592 4712
rect 8018 4700 8024 4752
rect 8076 4740 8082 4752
rect 8956 4740 8984 4780
rect 9398 4768 9404 4820
rect 9456 4768 9462 4820
rect 9858 4768 9864 4820
rect 9916 4808 9922 4820
rect 10137 4811 10195 4817
rect 10137 4808 10149 4811
rect 9916 4780 10149 4808
rect 9916 4768 9922 4780
rect 10137 4777 10149 4780
rect 10183 4777 10195 4811
rect 10137 4771 10195 4777
rect 12434 4768 12440 4820
rect 12492 4808 12498 4820
rect 22922 4808 22928 4820
rect 12492 4780 22928 4808
rect 12492 4768 12498 4780
rect 22922 4768 22928 4780
rect 22980 4768 22986 4820
rect 12342 4740 12348 4752
rect 8076 4712 8800 4740
rect 8956 4712 12348 4740
rect 8076 4700 8082 4712
rect 6549 4675 6607 4681
rect 6549 4641 6561 4675
rect 6595 4641 6607 4675
rect 6549 4635 6607 4641
rect 6638 4632 6644 4684
rect 6696 4672 6702 4684
rect 7009 4675 7067 4681
rect 7009 4672 7021 4675
rect 6696 4644 7021 4672
rect 6696 4632 6702 4644
rect 7009 4641 7021 4644
rect 7055 4641 7067 4675
rect 7009 4635 7067 4641
rect 7098 4632 7104 4684
rect 7156 4672 7162 4684
rect 8772 4681 8800 4712
rect 12342 4700 12348 4712
rect 12400 4700 12406 4752
rect 12618 4700 12624 4752
rect 12676 4700 12682 4752
rect 19242 4700 19248 4752
rect 19300 4740 19306 4752
rect 19300 4712 21588 4740
rect 19300 4700 19306 4712
rect 8757 4675 8815 4681
rect 7156 4644 8294 4672
rect 7156 4632 7162 4644
rect 3053 4607 3111 4613
rect 3053 4573 3065 4607
rect 3099 4573 3111 4607
rect 3053 4567 3111 4573
rect 2179 4508 2774 4536
rect 3068 4536 3096 4567
rect 3878 4564 3884 4616
rect 3936 4564 3942 4616
rect 4062 4564 4068 4616
rect 4120 4564 4126 4616
rect 4525 4607 4583 4613
rect 4525 4573 4537 4607
rect 4571 4573 4583 4607
rect 4525 4567 4583 4573
rect 5169 4607 5227 4613
rect 5169 4573 5181 4607
rect 5215 4604 5227 4607
rect 5258 4604 5264 4616
rect 5215 4576 5264 4604
rect 5215 4573 5227 4576
rect 5169 4567 5227 4573
rect 4080 4536 4108 4564
rect 3068 4508 4108 4536
rect 4540 4536 4568 4567
rect 5258 4564 5264 4576
rect 5316 4564 5322 4616
rect 5902 4564 5908 4616
rect 5960 4604 5966 4616
rect 5960 4576 6132 4604
rect 5960 4564 5966 4576
rect 6104 4536 6132 4576
rect 6730 4564 6736 4616
rect 6788 4564 6794 4616
rect 8266 4604 8294 4644
rect 8757 4641 8769 4675
rect 8803 4672 8815 4675
rect 8941 4675 8999 4681
rect 8941 4672 8953 4675
rect 8803 4644 8953 4672
rect 8803 4641 8815 4644
rect 8757 4635 8815 4641
rect 8941 4641 8953 4644
rect 8987 4672 8999 4675
rect 9030 4672 9036 4684
rect 8987 4644 9036 4672
rect 8987 4641 8999 4644
rect 8941 4635 8999 4641
rect 9030 4632 9036 4644
rect 9088 4632 9094 4684
rect 10597 4675 10655 4681
rect 10597 4641 10609 4675
rect 10643 4672 10655 4675
rect 10778 4672 10784 4684
rect 10643 4644 10784 4672
rect 10643 4641 10655 4644
rect 10597 4635 10655 4641
rect 10778 4632 10784 4644
rect 10836 4672 10842 4684
rect 12636 4672 12664 4700
rect 10836 4644 12664 4672
rect 10836 4632 10842 4644
rect 16114 4632 16120 4684
rect 16172 4672 16178 4684
rect 20898 4672 20904 4684
rect 16172 4644 20904 4672
rect 16172 4632 16178 4644
rect 20898 4632 20904 4644
rect 20956 4632 20962 4684
rect 9125 4607 9183 4613
rect 9125 4604 9137 4607
rect 8266 4576 9137 4604
rect 9125 4573 9137 4576
rect 9171 4573 9183 4607
rect 9125 4567 9183 4573
rect 9398 4564 9404 4616
rect 9456 4604 9462 4616
rect 9585 4607 9643 4613
rect 9585 4604 9597 4607
rect 9456 4576 9597 4604
rect 9456 4564 9462 4576
rect 9585 4573 9597 4576
rect 9631 4573 9643 4607
rect 9585 4567 9643 4573
rect 9674 4564 9680 4616
rect 9732 4604 9738 4616
rect 9861 4607 9919 4613
rect 9861 4604 9873 4607
rect 9732 4576 9873 4604
rect 9732 4564 9738 4576
rect 9861 4573 9873 4576
rect 9907 4573 9919 4607
rect 9861 4567 9919 4573
rect 16482 4564 16488 4616
rect 16540 4604 16546 4616
rect 21361 4607 21419 4613
rect 21361 4604 21373 4607
rect 16540 4576 21373 4604
rect 16540 4564 16546 4576
rect 21361 4573 21373 4576
rect 21407 4573 21419 4607
rect 21560 4604 21588 4712
rect 25041 4675 25099 4681
rect 25041 4641 25053 4675
rect 25087 4641 25099 4675
rect 25041 4635 25099 4641
rect 22833 4607 22891 4613
rect 22833 4604 22845 4607
rect 21560 4576 22845 4604
rect 21361 4567 21419 4573
rect 22833 4573 22845 4576
rect 22879 4573 22891 4607
rect 22833 4567 22891 4573
rect 22922 4564 22928 4616
rect 22980 4604 22986 4616
rect 24397 4607 24455 4613
rect 24397 4604 24409 4607
rect 22980 4576 24409 4604
rect 22980 4564 22986 4576
rect 24397 4573 24409 4576
rect 24443 4573 24455 4607
rect 24397 4567 24455 4573
rect 7098 4536 7104 4548
rect 4540 4508 6040 4536
rect 6104 4508 7104 4536
rect 2179 4505 2191 4508
rect 2133 4499 2191 4505
rect 1486 4428 1492 4480
rect 1544 4468 1550 4480
rect 3973 4471 4031 4477
rect 3973 4468 3985 4471
rect 1544 4440 3985 4468
rect 1544 4428 1550 4440
rect 3973 4437 3985 4440
rect 4019 4437 4031 4471
rect 6012 4468 6040 4508
rect 7098 4496 7104 4508
rect 7156 4496 7162 4548
rect 8754 4536 8760 4548
rect 8234 4508 8760 4536
rect 8754 4496 8760 4508
rect 8812 4496 8818 4548
rect 8864 4508 9720 4536
rect 8864 4468 8892 4508
rect 6012 4440 8892 4468
rect 3973 4431 4031 4437
rect 9306 4428 9312 4480
rect 9364 4428 9370 4480
rect 9692 4477 9720 4508
rect 22554 4496 22560 4548
rect 22612 4496 22618 4548
rect 24029 4539 24087 4545
rect 24029 4505 24041 4539
rect 24075 4536 24087 4539
rect 24854 4536 24860 4548
rect 24075 4508 24860 4536
rect 24075 4505 24087 4508
rect 24029 4499 24087 4505
rect 24854 4496 24860 4508
rect 24912 4496 24918 4548
rect 9677 4471 9735 4477
rect 9677 4437 9689 4471
rect 9723 4437 9735 4471
rect 9677 4431 9735 4437
rect 10965 4471 11023 4477
rect 10965 4437 10977 4471
rect 11011 4468 11023 4471
rect 11146 4468 11152 4480
rect 11011 4440 11152 4468
rect 11011 4437 11023 4440
rect 10965 4431 11023 4437
rect 11146 4428 11152 4440
rect 11204 4468 11210 4480
rect 12066 4468 12072 4480
rect 11204 4440 12072 4468
rect 11204 4428 11210 4440
rect 12066 4428 12072 4440
rect 12124 4428 12130 4480
rect 23658 4428 23664 4480
rect 23716 4468 23722 4480
rect 25056 4468 25084 4635
rect 25130 4632 25136 4684
rect 25188 4672 25194 4684
rect 26329 4675 26387 4681
rect 26329 4672 26341 4675
rect 25188 4644 26341 4672
rect 25188 4632 25194 4644
rect 26329 4641 26341 4644
rect 26375 4641 26387 4675
rect 26329 4635 26387 4641
rect 25866 4564 25872 4616
rect 25924 4564 25930 4616
rect 23716 4440 25084 4468
rect 23716 4428 23722 4440
rect 1104 4378 29048 4400
rect 1104 4326 7896 4378
rect 7948 4326 7960 4378
rect 8012 4326 8024 4378
rect 8076 4326 8088 4378
rect 8140 4326 8152 4378
rect 8204 4326 14842 4378
rect 14894 4326 14906 4378
rect 14958 4326 14970 4378
rect 15022 4326 15034 4378
rect 15086 4326 15098 4378
rect 15150 4326 21788 4378
rect 21840 4326 21852 4378
rect 21904 4326 21916 4378
rect 21968 4326 21980 4378
rect 22032 4326 22044 4378
rect 22096 4326 28734 4378
rect 28786 4326 28798 4378
rect 28850 4326 28862 4378
rect 28914 4326 28926 4378
rect 28978 4326 28990 4378
rect 29042 4326 29048 4378
rect 1104 4304 29048 4326
rect 1578 4224 1584 4276
rect 1636 4264 1642 4276
rect 1673 4267 1731 4273
rect 1673 4264 1685 4267
rect 1636 4236 1685 4264
rect 1636 4224 1642 4236
rect 1673 4233 1685 4236
rect 1719 4233 1731 4267
rect 1673 4227 1731 4233
rect 2498 4224 2504 4276
rect 2556 4224 2562 4276
rect 4157 4267 4215 4273
rect 4157 4233 4169 4267
rect 4203 4264 4215 4267
rect 8481 4267 8539 4273
rect 4203 4236 4292 4264
rect 4203 4233 4215 4236
rect 4157 4227 4215 4233
rect 842 4156 848 4208
rect 900 4196 906 4208
rect 1302 4196 1308 4208
rect 900 4168 1308 4196
rect 900 4156 906 4168
rect 1302 4156 1308 4168
rect 1360 4156 1366 4208
rect 2516 4196 2544 4224
rect 2685 4199 2743 4205
rect 2685 4196 2697 4199
rect 2516 4168 2697 4196
rect 2685 4165 2697 4168
rect 2731 4165 2743 4199
rect 2685 4159 2743 4165
rect 3142 4156 3148 4208
rect 3200 4156 3206 4208
rect 4264 4196 4292 4236
rect 8481 4233 8493 4267
rect 8527 4264 8539 4267
rect 8527 4236 9168 4264
rect 8527 4233 8539 4236
rect 8481 4227 8539 4233
rect 4080 4168 4292 4196
rect 1578 4088 1584 4140
rect 1636 4088 1642 4140
rect 2314 4088 2320 4140
rect 2372 4088 2378 4140
rect 2409 4063 2467 4069
rect 2409 4029 2421 4063
rect 2455 4029 2467 4063
rect 2409 4023 2467 4029
rect 1489 3927 1547 3933
rect 1489 3893 1501 3927
rect 1535 3924 1547 3927
rect 2314 3924 2320 3936
rect 1535 3896 2320 3924
rect 1535 3893 1547 3896
rect 1489 3887 1547 3893
rect 2314 3884 2320 3896
rect 2372 3884 2378 3936
rect 2424 3924 2452 4023
rect 3694 4020 3700 4072
rect 3752 4060 3758 4072
rect 4080 4060 4108 4168
rect 4154 4088 4160 4140
rect 4212 4088 4218 4140
rect 4264 4128 4292 4168
rect 4893 4199 4951 4205
rect 4893 4165 4905 4199
rect 4939 4196 4951 4199
rect 6178 4196 6184 4208
rect 4939 4168 6184 4196
rect 4939 4165 4951 4168
rect 4893 4159 4951 4165
rect 6178 4156 6184 4168
rect 6236 4196 6242 4208
rect 8570 4196 8576 4208
rect 6236 4168 7972 4196
rect 6236 4156 6242 4168
rect 5442 4128 5448 4140
rect 4264 4100 5448 4128
rect 5442 4088 5448 4100
rect 5500 4088 5506 4140
rect 5626 4088 5632 4140
rect 5684 4128 5690 4140
rect 5721 4131 5779 4137
rect 5721 4128 5733 4131
rect 5684 4100 5733 4128
rect 5684 4088 5690 4100
rect 5721 4097 5733 4100
rect 5767 4097 5779 4131
rect 5721 4091 5779 4097
rect 5810 4088 5816 4140
rect 5868 4088 5874 4140
rect 7944 4128 7972 4168
rect 8266 4168 8576 4196
rect 8266 4128 8294 4168
rect 8570 4156 8576 4168
rect 8628 4156 8634 4208
rect 9140 4196 9168 4236
rect 9214 4224 9220 4276
rect 9272 4224 9278 4276
rect 9306 4224 9312 4276
rect 9364 4264 9370 4276
rect 9364 4236 19334 4264
rect 9364 4224 9370 4236
rect 9674 4196 9680 4208
rect 9140 4168 9680 4196
rect 9674 4156 9680 4168
rect 9732 4156 9738 4208
rect 9766 4156 9772 4208
rect 9824 4156 9830 4208
rect 9858 4156 9864 4208
rect 9916 4156 9922 4208
rect 10778 4156 10784 4208
rect 10836 4156 10842 4208
rect 19306 4196 19334 4236
rect 22554 4224 22560 4276
rect 22612 4264 22618 4276
rect 28350 4264 28356 4276
rect 22612 4236 28356 4264
rect 22612 4224 22618 4236
rect 28350 4224 28356 4236
rect 28408 4224 28414 4276
rect 23290 4196 23296 4208
rect 19306 4168 23296 4196
rect 23290 4156 23296 4168
rect 23348 4156 23354 4208
rect 5920 4100 7880 4128
rect 7944 4100 8294 4128
rect 3752 4032 4108 4060
rect 4172 4060 4200 4088
rect 4985 4063 5043 4069
rect 4985 4060 4997 4063
rect 4172 4032 4997 4060
rect 3752 4020 3758 4032
rect 4985 4029 4997 4032
rect 5031 4029 5043 4063
rect 4985 4023 5043 4029
rect 5077 4063 5135 4069
rect 5077 4029 5089 4063
rect 5123 4060 5135 4063
rect 5537 4063 5595 4069
rect 5537 4060 5549 4063
rect 5123 4032 5549 4060
rect 5123 4029 5135 4032
rect 5077 4023 5135 4029
rect 5537 4029 5549 4032
rect 5583 4029 5595 4063
rect 5537 4023 5595 4029
rect 5092 3992 5120 4023
rect 5000 3964 5120 3992
rect 5000 3936 5028 3964
rect 5166 3952 5172 4004
rect 5224 3992 5230 4004
rect 5920 3992 5948 4100
rect 7852 4069 7880 4100
rect 9306 4088 9312 4140
rect 9364 4088 9370 4140
rect 9493 4131 9551 4137
rect 9493 4126 9505 4131
rect 9416 4098 9505 4126
rect 6917 4063 6975 4069
rect 6917 4060 6929 4063
rect 6196 4032 6929 4060
rect 6196 4001 6224 4032
rect 6917 4029 6929 4032
rect 6963 4029 6975 4063
rect 6917 4023 6975 4029
rect 7101 4063 7159 4069
rect 7101 4029 7113 4063
rect 7147 4029 7159 4063
rect 7101 4023 7159 4029
rect 7837 4063 7895 4069
rect 7837 4029 7849 4063
rect 7883 4029 7895 4063
rect 7837 4023 7895 4029
rect 8573 4063 8631 4069
rect 8573 4029 8585 4063
rect 8619 4029 8631 4063
rect 8573 4023 8631 4029
rect 5224 3964 5948 3992
rect 6181 3995 6239 4001
rect 5224 3952 5230 3964
rect 6181 3961 6193 3995
rect 6227 3961 6239 3995
rect 6181 3955 6239 3961
rect 6822 3952 6828 4004
rect 6880 3992 6886 4004
rect 7116 3992 7144 4023
rect 6880 3964 7144 3992
rect 6880 3952 6886 3964
rect 8294 3952 8300 4004
rect 8352 3992 8358 4004
rect 8588 3992 8616 4023
rect 8352 3964 8616 3992
rect 8352 3952 8358 3964
rect 8754 3952 8760 4004
rect 8812 3992 8818 4004
rect 9416 3992 9444 4098
rect 9493 4097 9505 4098
rect 9539 4097 9551 4131
rect 9784 4128 9812 4156
rect 9953 4131 10011 4137
rect 9953 4128 9965 4131
rect 9784 4100 9965 4128
rect 9493 4091 9551 4097
rect 9953 4097 9965 4100
rect 9999 4097 10011 4131
rect 9953 4091 10011 4097
rect 10226 4088 10232 4140
rect 10284 4088 10290 4140
rect 10505 4131 10563 4137
rect 10505 4097 10517 4131
rect 10551 4128 10563 4131
rect 10551 4100 10640 4128
rect 10551 4097 10563 4100
rect 10505 4091 10563 4097
rect 9677 4063 9735 4069
rect 9677 4029 9689 4063
rect 9723 4060 9735 4063
rect 10042 4060 10048 4072
rect 9723 4032 10048 4060
rect 9723 4029 9735 4032
rect 9677 4023 9735 4029
rect 10042 4020 10048 4032
rect 10100 4020 10106 4072
rect 10612 4060 10640 4100
rect 11330 4088 11336 4140
rect 11388 4128 11394 4140
rect 20257 4131 20315 4137
rect 20257 4128 20269 4131
rect 11388 4100 20269 4128
rect 11388 4088 11394 4100
rect 20257 4097 20269 4100
rect 20303 4097 20315 4131
rect 20257 4091 20315 4097
rect 22370 4088 22376 4140
rect 22428 4088 22434 4140
rect 23842 4088 23848 4140
rect 23900 4088 23906 4140
rect 24118 4088 24124 4140
rect 24176 4128 24182 4140
rect 25317 4131 25375 4137
rect 25317 4128 25329 4131
rect 24176 4100 25329 4128
rect 24176 4088 24182 4100
rect 25317 4097 25329 4100
rect 25363 4097 25375 4131
rect 25317 4091 25375 4097
rect 26602 4088 26608 4140
rect 26660 4128 26666 4140
rect 27154 4128 27160 4140
rect 26660 4100 27160 4128
rect 26660 4088 26666 4100
rect 27154 4088 27160 4100
rect 27212 4088 27218 4140
rect 10686 4060 10692 4072
rect 10612 4032 10692 4060
rect 10686 4020 10692 4032
rect 10744 4020 10750 4072
rect 21453 4063 21511 4069
rect 21453 4029 21465 4063
rect 21499 4029 21511 4063
rect 21453 4023 21511 4029
rect 10502 3992 10508 4004
rect 8812 3964 9444 3992
rect 10336 3964 10508 3992
rect 8812 3952 8818 3964
rect 3050 3924 3056 3936
rect 2424 3896 3056 3924
rect 3050 3884 3056 3896
rect 3108 3884 3114 3936
rect 4246 3884 4252 3936
rect 4304 3924 4310 3936
rect 4525 3927 4583 3933
rect 4525 3924 4537 3927
rect 4304 3896 4537 3924
rect 4304 3884 4310 3896
rect 4525 3893 4537 3896
rect 4571 3893 4583 3927
rect 4525 3887 4583 3893
rect 4982 3884 4988 3936
rect 5040 3884 5046 3936
rect 5902 3884 5908 3936
rect 5960 3924 5966 3936
rect 6365 3927 6423 3933
rect 6365 3924 6377 3927
rect 5960 3896 6377 3924
rect 5960 3884 5966 3896
rect 6365 3893 6377 3896
rect 6411 3893 6423 3927
rect 6365 3887 6423 3893
rect 7745 3927 7803 3933
rect 7745 3893 7757 3927
rect 7791 3924 7803 3927
rect 9582 3924 9588 3936
rect 7791 3896 9588 3924
rect 7791 3893 7803 3896
rect 7745 3887 7803 3893
rect 9582 3884 9588 3896
rect 9640 3884 9646 3936
rect 10045 3927 10103 3933
rect 10045 3893 10057 3927
rect 10091 3924 10103 3927
rect 10134 3924 10140 3936
rect 10091 3896 10140 3924
rect 10091 3893 10103 3896
rect 10045 3887 10103 3893
rect 10134 3884 10140 3896
rect 10192 3884 10198 3936
rect 10336 3933 10364 3964
rect 10502 3952 10508 3964
rect 10560 3952 10566 4004
rect 11793 3995 11851 4001
rect 11793 3961 11805 3995
rect 11839 3992 11851 3995
rect 12066 3992 12072 4004
rect 11839 3964 12072 3992
rect 11839 3961 11851 3964
rect 11793 3955 11851 3961
rect 12066 3952 12072 3964
rect 12124 3952 12130 4004
rect 21468 3992 21496 4023
rect 22278 4020 22284 4072
rect 22336 4060 22342 4072
rect 22833 4063 22891 4069
rect 22833 4060 22845 4063
rect 22336 4032 22845 4060
rect 22336 4020 22342 4032
rect 22833 4029 22845 4032
rect 22879 4029 22891 4063
rect 22833 4023 22891 4029
rect 23106 4020 23112 4072
rect 23164 4060 23170 4072
rect 24305 4063 24363 4069
rect 24305 4060 24317 4063
rect 23164 4032 24317 4060
rect 23164 4020 23170 4032
rect 24305 4029 24317 4032
rect 24351 4029 24363 4063
rect 25777 4063 25835 4069
rect 25777 4060 25789 4063
rect 24305 4023 24363 4029
rect 24826 4032 25789 4060
rect 21468 3964 23888 3992
rect 10321 3927 10379 3933
rect 10321 3893 10333 3927
rect 10367 3893 10379 3927
rect 10321 3887 10379 3893
rect 10594 3884 10600 3936
rect 10652 3924 10658 3936
rect 11241 3927 11299 3933
rect 11241 3924 11253 3927
rect 10652 3896 11253 3924
rect 10652 3884 10658 3896
rect 11241 3893 11253 3896
rect 11287 3924 11299 3927
rect 11882 3924 11888 3936
rect 11287 3896 11888 3924
rect 11287 3893 11299 3896
rect 11241 3887 11299 3893
rect 11882 3884 11888 3896
rect 11940 3924 11946 3936
rect 23750 3924 23756 3936
rect 11940 3896 23756 3924
rect 11940 3884 11946 3896
rect 23750 3884 23756 3896
rect 23808 3884 23814 3936
rect 23860 3924 23888 3964
rect 23934 3952 23940 4004
rect 23992 3992 23998 4004
rect 24826 3992 24854 4032
rect 25777 4029 25789 4032
rect 25823 4029 25835 4063
rect 25777 4023 25835 4029
rect 27433 4063 27491 4069
rect 27433 4029 27445 4063
rect 27479 4029 27491 4063
rect 27433 4023 27491 4029
rect 23992 3964 24854 3992
rect 23992 3952 23998 3964
rect 25130 3952 25136 4004
rect 25188 3992 25194 4004
rect 27448 3992 27476 4023
rect 25188 3964 27476 3992
rect 25188 3952 25194 3964
rect 25590 3924 25596 3936
rect 23860 3896 25596 3924
rect 25590 3884 25596 3896
rect 25648 3884 25654 3936
rect 1104 3834 28888 3856
rect 1104 3782 4423 3834
rect 4475 3782 4487 3834
rect 4539 3782 4551 3834
rect 4603 3782 4615 3834
rect 4667 3782 4679 3834
rect 4731 3782 11369 3834
rect 11421 3782 11433 3834
rect 11485 3782 11497 3834
rect 11549 3782 11561 3834
rect 11613 3782 11625 3834
rect 11677 3782 18315 3834
rect 18367 3782 18379 3834
rect 18431 3782 18443 3834
rect 18495 3782 18507 3834
rect 18559 3782 18571 3834
rect 18623 3782 25261 3834
rect 25313 3782 25325 3834
rect 25377 3782 25389 3834
rect 25441 3782 25453 3834
rect 25505 3782 25517 3834
rect 25569 3782 28888 3834
rect 1104 3760 28888 3782
rect 1673 3723 1731 3729
rect 1673 3689 1685 3723
rect 1719 3720 1731 3723
rect 2682 3720 2688 3732
rect 1719 3692 2688 3720
rect 1719 3689 1731 3692
rect 1673 3683 1731 3689
rect 2682 3680 2688 3692
rect 2740 3680 2746 3732
rect 3050 3680 3056 3732
rect 3108 3720 3114 3732
rect 3108 3692 3464 3720
rect 3108 3680 3114 3692
rect 3436 3593 3464 3692
rect 4522 3680 4528 3732
rect 4580 3720 4586 3732
rect 4982 3720 4988 3732
rect 4580 3692 4988 3720
rect 4580 3680 4586 3692
rect 4982 3680 4988 3692
rect 5040 3680 5046 3732
rect 5169 3723 5227 3729
rect 5169 3689 5181 3723
rect 5215 3720 5227 3723
rect 7742 3720 7748 3732
rect 5215 3692 7748 3720
rect 5215 3689 5227 3692
rect 5169 3683 5227 3689
rect 7742 3680 7748 3692
rect 7800 3680 7806 3732
rect 8478 3680 8484 3732
rect 8536 3720 8542 3732
rect 8573 3723 8631 3729
rect 8573 3720 8585 3723
rect 8536 3692 8585 3720
rect 8536 3680 8542 3692
rect 8573 3689 8585 3692
rect 8619 3689 8631 3723
rect 8573 3683 8631 3689
rect 8846 3680 8852 3732
rect 8904 3680 8910 3732
rect 10226 3680 10232 3732
rect 10284 3720 10290 3732
rect 10413 3723 10471 3729
rect 10413 3720 10425 3723
rect 10284 3692 10425 3720
rect 10284 3680 10290 3692
rect 10413 3689 10425 3692
rect 10459 3689 10471 3723
rect 10413 3683 10471 3689
rect 10689 3723 10747 3729
rect 10689 3689 10701 3723
rect 10735 3720 10747 3723
rect 10870 3720 10876 3732
rect 10735 3692 10876 3720
rect 10735 3689 10747 3692
rect 10689 3683 10747 3689
rect 10870 3680 10876 3692
rect 10928 3680 10934 3732
rect 10962 3680 10968 3732
rect 11020 3720 11026 3732
rect 11333 3723 11391 3729
rect 11333 3720 11345 3723
rect 11020 3692 11345 3720
rect 11020 3680 11026 3692
rect 11333 3689 11345 3692
rect 11379 3689 11391 3723
rect 11333 3683 11391 3689
rect 11882 3680 11888 3732
rect 11940 3680 11946 3732
rect 12066 3680 12072 3732
rect 12124 3720 12130 3732
rect 12161 3723 12219 3729
rect 12161 3720 12173 3723
rect 12124 3692 12173 3720
rect 12124 3680 12130 3692
rect 12161 3689 12173 3692
rect 12207 3689 12219 3723
rect 12161 3683 12219 3689
rect 24118 3680 24124 3732
rect 24176 3680 24182 3732
rect 27154 3680 27160 3732
rect 27212 3720 27218 3732
rect 27525 3723 27583 3729
rect 27525 3720 27537 3723
rect 27212 3692 27537 3720
rect 27212 3680 27218 3692
rect 27525 3689 27537 3692
rect 27571 3689 27583 3723
rect 27525 3683 27583 3689
rect 8864 3652 8892 3680
rect 6656 3624 8892 3652
rect 3421 3587 3479 3593
rect 3421 3553 3433 3587
rect 3467 3584 3479 3587
rect 4062 3584 4068 3596
rect 3467 3556 4068 3584
rect 3467 3553 3479 3556
rect 3421 3547 3479 3553
rect 4062 3544 4068 3556
rect 4120 3584 4126 3596
rect 5261 3587 5319 3593
rect 5261 3584 5273 3587
rect 4120 3556 5273 3584
rect 4120 3544 4126 3556
rect 5261 3553 5273 3556
rect 5307 3553 5319 3587
rect 5261 3547 5319 3553
rect 5537 3587 5595 3593
rect 5537 3553 5549 3587
rect 5583 3584 5595 3587
rect 5902 3584 5908 3596
rect 5583 3556 5908 3584
rect 5583 3553 5595 3556
rect 5537 3547 5595 3553
rect 5902 3544 5908 3556
rect 5960 3544 5966 3596
rect 1489 3519 1547 3525
rect 1489 3485 1501 3519
rect 1535 3516 1547 3519
rect 2590 3516 2596 3528
rect 1535 3488 2596 3516
rect 1535 3485 1547 3488
rect 1489 3479 1547 3485
rect 2590 3476 2596 3488
rect 2648 3476 2654 3528
rect 2774 3476 2780 3528
rect 2832 3516 2838 3528
rect 3154 3519 3212 3525
rect 3154 3516 3166 3519
rect 2832 3488 3166 3516
rect 2832 3476 2838 3488
rect 3154 3485 3166 3488
rect 3200 3485 3212 3519
rect 3154 3479 3212 3485
rect 3326 3476 3332 3528
rect 3384 3516 3390 3528
rect 3789 3519 3847 3525
rect 3789 3516 3801 3519
rect 3384 3488 3801 3516
rect 3384 3476 3390 3488
rect 3789 3485 3801 3488
rect 3835 3485 3847 3519
rect 3789 3479 3847 3485
rect 3878 3476 3884 3528
rect 3936 3516 3942 3528
rect 3936 3488 4660 3516
rect 3936 3476 3942 3488
rect 1578 3408 1584 3460
rect 1636 3448 1642 3460
rect 1636 3420 2820 3448
rect 1636 3408 1642 3420
rect 2038 3340 2044 3392
rect 2096 3340 2102 3392
rect 2792 3380 2820 3420
rect 2866 3408 2872 3460
rect 2924 3448 2930 3460
rect 3050 3448 3056 3460
rect 2924 3420 3056 3448
rect 2924 3408 2930 3420
rect 3050 3408 3056 3420
rect 3108 3408 3114 3460
rect 4522 3408 4528 3460
rect 4580 3408 4586 3460
rect 4632 3448 4660 3488
rect 4798 3476 4804 3528
rect 4856 3476 4862 3528
rect 4985 3519 5043 3525
rect 4985 3485 4997 3519
rect 5031 3485 5043 3519
rect 6656 3502 6684 3624
rect 10042 3612 10048 3664
rect 10100 3652 10106 3664
rect 20346 3652 20352 3664
rect 10100 3624 20352 3652
rect 10100 3612 10106 3624
rect 20346 3612 20352 3624
rect 20404 3612 20410 3664
rect 21450 3612 21456 3664
rect 21508 3652 21514 3664
rect 21508 3624 22048 3652
rect 21508 3612 21514 3624
rect 22020 3593 22048 3624
rect 22005 3587 22063 3593
rect 6840 3556 8984 3584
rect 4985 3479 5043 3485
rect 5000 3448 5028 3479
rect 4632 3420 5028 3448
rect 3878 3380 3884 3392
rect 2792 3352 3884 3380
rect 3878 3340 3884 3352
rect 3936 3340 3942 3392
rect 4890 3340 4896 3392
rect 4948 3380 4954 3392
rect 6840 3380 6868 3556
rect 7098 3476 7104 3528
rect 7156 3516 7162 3528
rect 7285 3519 7343 3525
rect 7285 3516 7297 3519
rect 7156 3488 7297 3516
rect 7156 3476 7162 3488
rect 7285 3485 7297 3488
rect 7331 3516 7343 3519
rect 7466 3516 7472 3528
rect 7331 3488 7472 3516
rect 7331 3485 7343 3488
rect 7285 3479 7343 3485
rect 7466 3476 7472 3488
rect 7524 3476 7530 3528
rect 7561 3519 7619 3525
rect 7561 3485 7573 3519
rect 7607 3516 7619 3519
rect 7650 3516 7656 3528
rect 7607 3488 7656 3516
rect 7607 3485 7619 3488
rect 7561 3479 7619 3485
rect 7650 3476 7656 3488
rect 7708 3476 7714 3528
rect 7926 3476 7932 3528
rect 7984 3476 7990 3528
rect 8956 3525 8984 3556
rect 10428 3556 21588 3584
rect 8941 3519 8999 3525
rect 8941 3485 8953 3519
rect 8987 3485 8999 3519
rect 8941 3479 8999 3485
rect 9582 3476 9588 3528
rect 9640 3516 9646 3528
rect 9769 3519 9827 3525
rect 9769 3516 9781 3519
rect 9640 3488 9781 3516
rect 9640 3476 9646 3488
rect 9769 3485 9781 3488
rect 9815 3485 9827 3519
rect 9769 3479 9827 3485
rect 7190 3408 7196 3460
rect 7248 3408 7254 3460
rect 7745 3451 7803 3457
rect 7745 3417 7757 3451
rect 7791 3448 7803 3451
rect 10428 3448 10456 3556
rect 10505 3519 10563 3525
rect 10505 3485 10517 3519
rect 10551 3485 10563 3519
rect 10505 3479 10563 3485
rect 7791 3420 10456 3448
rect 7791 3417 7803 3420
rect 7745 3411 7803 3417
rect 4948 3352 6868 3380
rect 7208 3380 7236 3408
rect 10520 3392 10548 3479
rect 10962 3476 10968 3528
rect 11020 3476 11026 3528
rect 11241 3519 11299 3525
rect 11241 3485 11253 3519
rect 11287 3516 11299 3519
rect 11330 3516 11336 3528
rect 11287 3488 11336 3516
rect 11287 3485 11299 3488
rect 11241 3479 11299 3485
rect 11330 3476 11336 3488
rect 11388 3476 11394 3528
rect 11517 3519 11575 3525
rect 11517 3485 11529 3519
rect 11563 3485 11575 3519
rect 11517 3479 11575 3485
rect 11146 3408 11152 3460
rect 11204 3448 11210 3460
rect 11532 3448 11560 3479
rect 20070 3476 20076 3528
rect 20128 3476 20134 3528
rect 21560 3525 21588 3556
rect 22005 3553 22017 3587
rect 22051 3553 22063 3587
rect 22005 3547 22063 3553
rect 22830 3544 22836 3596
rect 22888 3584 22894 3596
rect 24857 3587 24915 3593
rect 24857 3584 24869 3587
rect 22888 3556 24869 3584
rect 22888 3544 22894 3556
rect 24857 3553 24869 3556
rect 24903 3553 24915 3587
rect 26329 3587 26387 3593
rect 26329 3584 26341 3587
rect 24857 3547 24915 3553
rect 25240 3556 26341 3584
rect 21545 3519 21603 3525
rect 21545 3485 21557 3519
rect 21591 3485 21603 3519
rect 21545 3479 21603 3485
rect 24394 3476 24400 3528
rect 24452 3476 24458 3528
rect 11204 3420 11560 3448
rect 21269 3451 21327 3457
rect 11204 3408 11210 3420
rect 21269 3417 21281 3451
rect 21315 3448 21327 3451
rect 21315 3420 22094 3448
rect 21315 3417 21327 3420
rect 21269 3411 21327 3417
rect 8754 3380 8760 3392
rect 7208 3352 8760 3380
rect 4948 3340 4954 3352
rect 8754 3340 8760 3352
rect 8812 3340 8818 3392
rect 9585 3383 9643 3389
rect 9585 3349 9597 3383
rect 9631 3380 9643 3383
rect 10410 3380 10416 3392
rect 9631 3352 10416 3380
rect 9631 3349 9643 3352
rect 9585 3343 9643 3349
rect 10410 3340 10416 3352
rect 10468 3340 10474 3392
rect 10502 3340 10508 3392
rect 10560 3340 10566 3392
rect 10778 3340 10784 3392
rect 10836 3340 10842 3392
rect 11054 3340 11060 3392
rect 11112 3340 11118 3392
rect 22066 3380 22094 3420
rect 24210 3408 24216 3460
rect 24268 3448 24274 3460
rect 25240 3448 25268 3556
rect 26329 3553 26341 3556
rect 26375 3553 26387 3587
rect 26329 3547 26387 3553
rect 25866 3476 25872 3528
rect 25924 3476 25930 3528
rect 28537 3519 28595 3525
rect 28537 3485 28549 3519
rect 28583 3516 28595 3519
rect 29454 3516 29460 3528
rect 28583 3488 29460 3516
rect 28583 3485 28595 3488
rect 28537 3479 28595 3485
rect 29454 3476 29460 3488
rect 29512 3476 29518 3528
rect 24268 3420 25268 3448
rect 24268 3408 24274 3420
rect 27062 3380 27068 3392
rect 22066 3352 27068 3380
rect 27062 3340 27068 3352
rect 27120 3340 27126 3392
rect 1104 3290 29048 3312
rect 1104 3238 7896 3290
rect 7948 3238 7960 3290
rect 8012 3238 8024 3290
rect 8076 3238 8088 3290
rect 8140 3238 8152 3290
rect 8204 3238 14842 3290
rect 14894 3238 14906 3290
rect 14958 3238 14970 3290
rect 15022 3238 15034 3290
rect 15086 3238 15098 3290
rect 15150 3238 21788 3290
rect 21840 3238 21852 3290
rect 21904 3238 21916 3290
rect 21968 3238 21980 3290
rect 22032 3238 22044 3290
rect 22096 3238 28734 3290
rect 28786 3238 28798 3290
rect 28850 3238 28862 3290
rect 28914 3238 28926 3290
rect 28978 3238 28990 3290
rect 29042 3238 29048 3290
rect 1104 3216 29048 3238
rect 1946 3136 1952 3188
rect 2004 3176 2010 3188
rect 2225 3179 2283 3185
rect 2225 3176 2237 3179
rect 2004 3148 2237 3176
rect 2004 3136 2010 3148
rect 2225 3145 2237 3148
rect 2271 3145 2283 3179
rect 2225 3139 2283 3145
rect 2314 3136 2320 3188
rect 2372 3176 2378 3188
rect 2372 3148 4200 3176
rect 2372 3136 2378 3148
rect 2133 3111 2191 3117
rect 2133 3077 2145 3111
rect 2179 3108 2191 3111
rect 4172 3108 4200 3148
rect 5442 3136 5448 3188
rect 5500 3176 5506 3188
rect 5500 3148 6316 3176
rect 5500 3136 5506 3148
rect 2179 3080 4016 3108
rect 4172 3080 4922 3108
rect 2179 3077 2191 3080
rect 2133 3071 2191 3077
rect 2593 3043 2651 3049
rect 2593 3009 2605 3043
rect 2639 3040 2651 3043
rect 2639 3012 3004 3040
rect 2639 3009 2651 3012
rect 2593 3003 2651 3009
rect 1581 2975 1639 2981
rect 1581 2941 1593 2975
rect 1627 2941 1639 2975
rect 1581 2935 1639 2941
rect 1596 2904 1624 2935
rect 1854 2932 1860 2984
rect 1912 2972 1918 2984
rect 2685 2975 2743 2981
rect 2685 2972 2697 2975
rect 1912 2944 2697 2972
rect 1912 2932 1918 2944
rect 2685 2941 2697 2944
rect 2731 2941 2743 2975
rect 2685 2935 2743 2941
rect 2866 2932 2872 2984
rect 2924 2932 2930 2984
rect 2976 2972 3004 3012
rect 3050 3000 3056 3052
rect 3108 3000 3114 3052
rect 3694 3000 3700 3052
rect 3752 3000 3758 3052
rect 3878 3000 3884 3052
rect 3936 3000 3942 3052
rect 3712 2972 3740 3000
rect 2976 2944 3740 2972
rect 3988 2972 4016 3080
rect 6178 3068 6184 3120
rect 6236 3068 6242 3120
rect 6288 3108 6316 3148
rect 7558 3136 7564 3188
rect 7616 3136 7622 3188
rect 8297 3179 8355 3185
rect 8297 3145 8309 3179
rect 8343 3176 8355 3179
rect 8386 3176 8392 3188
rect 8343 3148 8392 3176
rect 8343 3145 8355 3148
rect 8297 3139 8355 3145
rect 8386 3136 8392 3148
rect 8444 3136 8450 3188
rect 9033 3179 9091 3185
rect 9033 3145 9045 3179
rect 9079 3176 9091 3179
rect 9398 3176 9404 3188
rect 9079 3148 9404 3176
rect 9079 3145 9091 3148
rect 9033 3139 9091 3145
rect 9398 3136 9404 3148
rect 9456 3136 9462 3188
rect 10134 3176 10140 3188
rect 9646 3148 10140 3176
rect 9306 3108 9312 3120
rect 6288 3080 9312 3108
rect 9306 3068 9312 3080
rect 9364 3068 9370 3120
rect 4062 3000 4068 3052
rect 4120 3040 4126 3052
rect 4157 3043 4215 3049
rect 4157 3040 4169 3043
rect 4120 3012 4169 3040
rect 4120 3000 4126 3012
rect 4157 3009 4169 3012
rect 4203 3009 4215 3043
rect 6196 3040 6224 3068
rect 6365 3043 6423 3049
rect 6365 3040 6377 3043
rect 6196 3012 6377 3040
rect 4157 3003 4215 3009
rect 6365 3009 6377 3012
rect 6411 3009 6423 3043
rect 6365 3003 6423 3009
rect 6546 3000 6552 3052
rect 6604 3000 6610 3052
rect 7466 3000 7472 3052
rect 7524 3040 7530 3052
rect 9646 3040 9674 3148
rect 10134 3136 10140 3148
rect 10192 3136 10198 3188
rect 10410 3136 10416 3188
rect 10468 3136 10474 3188
rect 10502 3136 10508 3188
rect 10560 3176 10566 3188
rect 10597 3179 10655 3185
rect 10597 3176 10609 3179
rect 10560 3148 10609 3176
rect 10560 3136 10566 3148
rect 10597 3145 10609 3148
rect 10643 3145 10655 3179
rect 10597 3139 10655 3145
rect 11238 3136 11244 3188
rect 11296 3176 11302 3188
rect 11517 3179 11575 3185
rect 11517 3176 11529 3179
rect 11296 3148 11529 3176
rect 11296 3136 11302 3148
rect 11517 3145 11529 3148
rect 11563 3145 11575 3179
rect 11517 3139 11575 3145
rect 11793 3179 11851 3185
rect 11793 3145 11805 3179
rect 11839 3176 11851 3179
rect 11882 3176 11888 3188
rect 11839 3148 11888 3176
rect 11839 3145 11851 3148
rect 11793 3139 11851 3145
rect 11882 3136 11888 3148
rect 11940 3136 11946 3188
rect 11974 3136 11980 3188
rect 12032 3176 12038 3188
rect 12069 3179 12127 3185
rect 12069 3176 12081 3179
rect 12032 3148 12081 3176
rect 12032 3136 12038 3148
rect 12069 3145 12081 3148
rect 12115 3145 12127 3179
rect 12069 3139 12127 3145
rect 12342 3136 12348 3188
rect 12400 3136 12406 3188
rect 23382 3176 23388 3188
rect 22066 3148 23388 3176
rect 9950 3068 9956 3120
rect 10008 3068 10014 3120
rect 10428 3108 10456 3136
rect 19981 3111 20039 3117
rect 10428 3080 12434 3108
rect 7524 3012 9674 3040
rect 9968 3040 9996 3068
rect 10778 3040 10784 3052
rect 9968 3012 10784 3040
rect 7524 3000 7530 3012
rect 10778 3000 10784 3012
rect 10836 3000 10842 3052
rect 11698 3000 11704 3052
rect 11756 3000 11762 3052
rect 11977 3043 12035 3049
rect 11977 3009 11989 3043
rect 12023 3009 12035 3043
rect 11977 3003 12035 3009
rect 4433 2975 4491 2981
rect 4433 2972 4445 2975
rect 3988 2944 4445 2972
rect 4433 2941 4445 2944
rect 4479 2941 4491 2975
rect 4433 2935 4491 2941
rect 7009 2975 7067 2981
rect 7009 2941 7021 2975
rect 7055 2972 7067 2975
rect 7374 2972 7380 2984
rect 7055 2944 7380 2972
rect 7055 2941 7067 2944
rect 7009 2935 7067 2941
rect 7374 2932 7380 2944
rect 7432 2932 7438 2984
rect 7745 2975 7803 2981
rect 7745 2941 7757 2975
rect 7791 2972 7803 2975
rect 8202 2972 8208 2984
rect 7791 2944 8208 2972
rect 7791 2941 7803 2944
rect 7745 2935 7803 2941
rect 8202 2932 8208 2944
rect 8260 2932 8266 2984
rect 8481 2975 8539 2981
rect 8481 2941 8493 2975
rect 8527 2972 8539 2975
rect 8754 2972 8760 2984
rect 8527 2944 8760 2972
rect 8527 2941 8539 2944
rect 8481 2935 8539 2941
rect 8754 2932 8760 2944
rect 8812 2932 8818 2984
rect 9214 2932 9220 2984
rect 9272 2932 9278 2984
rect 9490 2932 9496 2984
rect 9548 2972 9554 2984
rect 9861 2975 9919 2981
rect 9861 2972 9873 2975
rect 9548 2944 9873 2972
rect 9548 2932 9554 2944
rect 9861 2941 9873 2944
rect 9907 2941 9919 2975
rect 9861 2935 9919 2941
rect 10134 2932 10140 2984
rect 10192 2972 10198 2984
rect 10413 2975 10471 2981
rect 10413 2972 10425 2975
rect 10192 2944 10425 2972
rect 10192 2932 10198 2944
rect 10413 2941 10425 2944
rect 10459 2941 10471 2975
rect 10413 2935 10471 2941
rect 10594 2932 10600 2984
rect 10652 2972 10658 2984
rect 11149 2975 11207 2981
rect 11149 2972 11161 2975
rect 10652 2944 11161 2972
rect 10652 2932 10658 2944
rect 11149 2941 11161 2944
rect 11195 2941 11207 2975
rect 11149 2935 11207 2941
rect 1596 2876 4292 2904
rect 4264 2848 4292 2876
rect 6730 2864 6736 2916
rect 6788 2864 6794 2916
rect 9674 2864 9680 2916
rect 9732 2904 9738 2916
rect 11992 2904 12020 3003
rect 12250 3000 12256 3052
rect 12308 3000 12314 3052
rect 12406 3040 12434 3080
rect 19981 3077 19993 3111
rect 20027 3108 20039 3111
rect 22066 3108 22094 3148
rect 23382 3136 23388 3148
rect 23440 3136 23446 3188
rect 26786 3108 26792 3120
rect 20027 3080 22094 3108
rect 22204 3080 26792 3108
rect 20027 3077 20039 3080
rect 19981 3071 20039 3077
rect 12529 3043 12587 3049
rect 12529 3040 12541 3043
rect 12406 3012 12541 3040
rect 12529 3009 12541 3012
rect 12575 3009 12587 3043
rect 12529 3003 12587 3009
rect 15838 3000 15844 3052
rect 15896 3040 15902 3052
rect 18785 3043 18843 3049
rect 18785 3040 18797 3043
rect 15896 3012 18797 3040
rect 15896 3000 15902 3012
rect 18785 3009 18797 3012
rect 18831 3009 18843 3043
rect 18785 3003 18843 3009
rect 18874 3000 18880 3052
rect 18932 3040 18938 3052
rect 20257 3043 20315 3049
rect 20257 3040 20269 3043
rect 18932 3012 20269 3040
rect 18932 3000 18938 3012
rect 20257 3009 20269 3012
rect 20303 3009 20315 3043
rect 20257 3003 20315 3009
rect 21818 3000 21824 3052
rect 21876 3000 21882 3052
rect 21453 2975 21511 2981
rect 21453 2941 21465 2975
rect 21499 2972 21511 2975
rect 22204 2972 22232 3080
rect 26786 3068 26792 3080
rect 26844 3068 26850 3120
rect 23290 3000 23296 3052
rect 23348 3000 23354 3052
rect 23400 3012 23888 3040
rect 21499 2944 22232 2972
rect 22281 2975 22339 2981
rect 21499 2941 21511 2944
rect 21453 2935 21511 2941
rect 22281 2941 22293 2975
rect 22327 2941 22339 2975
rect 22281 2935 22339 2941
rect 9732 2876 12020 2904
rect 9732 2864 9738 2876
rect 21358 2864 21364 2916
rect 21416 2904 21422 2916
rect 22296 2904 22324 2935
rect 22554 2932 22560 2984
rect 22612 2972 22618 2984
rect 23400 2972 23428 3012
rect 22612 2944 23428 2972
rect 23753 2975 23811 2981
rect 22612 2932 22618 2944
rect 23753 2941 23765 2975
rect 23799 2941 23811 2975
rect 23860 2972 23888 3012
rect 24946 3000 24952 3052
rect 25004 3000 25010 3052
rect 26970 3000 26976 3052
rect 27028 3000 27034 3052
rect 25225 2975 25283 2981
rect 25225 2972 25237 2975
rect 23860 2944 25237 2972
rect 23753 2935 23811 2941
rect 25225 2941 25237 2944
rect 25271 2941 25283 2975
rect 25225 2935 25283 2941
rect 27433 2975 27491 2981
rect 27433 2941 27445 2975
rect 27479 2941 27491 2975
rect 27433 2935 27491 2941
rect 21416 2876 22324 2904
rect 21416 2864 21422 2876
rect 1762 2796 1768 2848
rect 1820 2836 1826 2848
rect 3786 2836 3792 2848
rect 1820 2808 3792 2836
rect 1820 2796 1826 2808
rect 3786 2796 3792 2808
rect 3844 2796 3850 2848
rect 4246 2796 4252 2848
rect 4304 2796 4310 2848
rect 4798 2796 4804 2848
rect 4856 2836 4862 2848
rect 8294 2836 8300 2848
rect 4856 2808 8300 2836
rect 4856 2796 4862 2808
rect 8294 2796 8300 2808
rect 8352 2796 8358 2848
rect 9769 2839 9827 2845
rect 9769 2805 9781 2839
rect 9815 2836 9827 2839
rect 11330 2836 11336 2848
rect 9815 2808 11336 2836
rect 9815 2805 9827 2808
rect 9769 2799 9827 2805
rect 11330 2796 11336 2808
rect 11388 2796 11394 2848
rect 21542 2796 21548 2848
rect 21600 2836 21606 2848
rect 23768 2836 23796 2935
rect 24670 2864 24676 2916
rect 24728 2904 24734 2916
rect 27448 2904 27476 2935
rect 24728 2876 27476 2904
rect 24728 2864 24734 2876
rect 21600 2808 23796 2836
rect 21600 2796 21606 2808
rect 1104 2746 28888 2768
rect 1104 2694 4423 2746
rect 4475 2694 4487 2746
rect 4539 2694 4551 2746
rect 4603 2694 4615 2746
rect 4667 2694 4679 2746
rect 4731 2694 11369 2746
rect 11421 2694 11433 2746
rect 11485 2694 11497 2746
rect 11549 2694 11561 2746
rect 11613 2694 11625 2746
rect 11677 2694 18315 2746
rect 18367 2694 18379 2746
rect 18431 2694 18443 2746
rect 18495 2694 18507 2746
rect 18559 2694 18571 2746
rect 18623 2694 25261 2746
rect 25313 2694 25325 2746
rect 25377 2694 25389 2746
rect 25441 2694 25453 2746
rect 25505 2694 25517 2746
rect 25569 2694 28888 2746
rect 1104 2672 28888 2694
rect 3973 2635 4031 2641
rect 3973 2601 3985 2635
rect 4019 2632 4031 2635
rect 6270 2632 6276 2644
rect 4019 2604 6276 2632
rect 4019 2601 4031 2604
rect 3973 2595 4031 2601
rect 6270 2592 6276 2604
rect 6328 2592 6334 2644
rect 6549 2635 6607 2641
rect 6549 2601 6561 2635
rect 6595 2632 6607 2635
rect 7006 2632 7012 2644
rect 6595 2604 7012 2632
rect 6595 2601 6607 2604
rect 6549 2595 6607 2601
rect 7006 2592 7012 2604
rect 7064 2592 7070 2644
rect 8021 2635 8079 2641
rect 8021 2601 8033 2635
rect 8067 2632 8079 2635
rect 9674 2632 9680 2644
rect 8067 2604 9680 2632
rect 8067 2601 8079 2604
rect 8021 2595 8079 2601
rect 9674 2592 9680 2604
rect 9732 2592 9738 2644
rect 10502 2592 10508 2644
rect 10560 2592 10566 2644
rect 11333 2635 11391 2641
rect 11333 2601 11345 2635
rect 11379 2632 11391 2635
rect 11698 2632 11704 2644
rect 11379 2604 11704 2632
rect 11379 2601 11391 2604
rect 11333 2595 11391 2601
rect 11698 2592 11704 2604
rect 11756 2592 11762 2644
rect 12158 2592 12164 2644
rect 12216 2632 12222 2644
rect 12253 2635 12311 2641
rect 12253 2632 12265 2635
rect 12216 2604 12265 2632
rect 12216 2592 12222 2604
rect 12253 2601 12265 2604
rect 12299 2601 12311 2635
rect 12253 2595 12311 2601
rect 12526 2592 12532 2644
rect 12584 2592 12590 2644
rect 7098 2564 7104 2576
rect 5552 2536 7104 2564
rect 2314 2456 2320 2508
rect 2372 2456 2378 2508
rect 2590 2456 2596 2508
rect 2648 2496 2654 2508
rect 5552 2505 5580 2536
rect 7098 2524 7104 2536
rect 7156 2524 7162 2576
rect 9125 2567 9183 2573
rect 9125 2533 9137 2567
rect 9171 2564 9183 2567
rect 10520 2564 10548 2592
rect 9171 2536 10548 2564
rect 9171 2533 9183 2536
rect 9125 2527 9183 2533
rect 10962 2524 10968 2576
rect 11020 2564 11026 2576
rect 11020 2536 13032 2564
rect 11020 2524 11026 2536
rect 4065 2499 4123 2505
rect 4065 2496 4077 2499
rect 2648 2468 4077 2496
rect 2648 2456 2654 2468
rect 4065 2465 4077 2468
rect 4111 2465 4123 2499
rect 5537 2499 5595 2505
rect 4065 2459 4123 2465
rect 4724 2468 5488 2496
rect 1581 2431 1639 2437
rect 1581 2397 1593 2431
rect 1627 2428 1639 2431
rect 1627 2400 2774 2428
rect 1627 2397 1639 2400
rect 1581 2391 1639 2397
rect 2746 2360 2774 2400
rect 3050 2388 3056 2440
rect 3108 2388 3114 2440
rect 4724 2437 4752 2468
rect 3789 2431 3847 2437
rect 3789 2397 3801 2431
rect 3835 2397 3847 2431
rect 3789 2391 3847 2397
rect 4709 2431 4767 2437
rect 4709 2397 4721 2431
rect 4755 2397 4767 2431
rect 4709 2391 4767 2397
rect 4893 2431 4951 2437
rect 4893 2397 4905 2431
rect 4939 2428 4951 2431
rect 5350 2428 5356 2440
rect 4939 2400 5356 2428
rect 4939 2397 4951 2400
rect 4893 2391 4951 2397
rect 3804 2360 3832 2391
rect 5350 2388 5356 2400
rect 5408 2388 5414 2440
rect 5460 2428 5488 2468
rect 5537 2465 5549 2499
rect 5583 2465 5595 2499
rect 5537 2459 5595 2465
rect 6178 2456 6184 2508
rect 6236 2456 6242 2508
rect 8113 2499 8171 2505
rect 8113 2496 8125 2499
rect 6380 2468 8125 2496
rect 6270 2428 6276 2440
rect 5460 2400 6276 2428
rect 6270 2388 6276 2400
rect 6328 2388 6334 2440
rect 6380 2437 6408 2468
rect 8113 2465 8125 2468
rect 8159 2465 8171 2499
rect 9490 2496 9496 2508
rect 8113 2459 8171 2465
rect 8956 2468 9496 2496
rect 6365 2431 6423 2437
rect 6365 2397 6377 2431
rect 6411 2397 6423 2431
rect 6365 2391 6423 2397
rect 7285 2431 7343 2437
rect 7285 2397 7297 2431
rect 7331 2397 7343 2431
rect 7285 2391 7343 2397
rect 7469 2431 7527 2437
rect 7469 2397 7481 2431
rect 7515 2428 7527 2431
rect 8478 2428 8484 2440
rect 7515 2400 8484 2428
rect 7515 2397 7527 2400
rect 7469 2391 7527 2397
rect 6641 2363 6699 2369
rect 6641 2360 6653 2363
rect 2746 2332 3740 2360
rect 3804 2332 6653 2360
rect 2130 2252 2136 2304
rect 2188 2252 2194 2304
rect 2866 2252 2872 2304
rect 2924 2252 2930 2304
rect 3602 2252 3608 2304
rect 3660 2252 3666 2304
rect 3712 2292 3740 2332
rect 6641 2329 6653 2332
rect 6687 2329 6699 2363
rect 7300 2360 7328 2391
rect 8478 2388 8484 2400
rect 8536 2388 8542 2440
rect 8757 2431 8815 2437
rect 8757 2397 8769 2431
rect 8803 2428 8815 2431
rect 8846 2428 8852 2440
rect 8803 2400 8852 2428
rect 8803 2397 8815 2400
rect 8757 2391 8815 2397
rect 8846 2388 8852 2400
rect 8904 2388 8910 2440
rect 8956 2437 8984 2468
rect 9490 2456 9496 2468
rect 9548 2456 9554 2508
rect 10597 2499 10655 2505
rect 10597 2465 10609 2499
rect 10643 2496 10655 2499
rect 10643 2468 12756 2496
rect 10643 2465 10655 2468
rect 10597 2459 10655 2465
rect 8941 2431 8999 2437
rect 8941 2397 8953 2431
rect 8987 2397 8999 2431
rect 8941 2391 8999 2397
rect 9309 2431 9367 2437
rect 9309 2397 9321 2431
rect 9355 2428 9367 2431
rect 9858 2428 9864 2440
rect 9355 2400 9864 2428
rect 9355 2397 9367 2400
rect 9309 2391 9367 2397
rect 9858 2388 9864 2400
rect 9916 2388 9922 2440
rect 10045 2431 10103 2437
rect 10045 2397 10057 2431
rect 10091 2428 10103 2431
rect 10686 2428 10692 2440
rect 10091 2400 10692 2428
rect 10091 2397 10103 2400
rect 10045 2391 10103 2397
rect 10686 2388 10692 2400
rect 10744 2388 10750 2440
rect 10778 2388 10784 2440
rect 10836 2388 10842 2440
rect 11054 2388 11060 2440
rect 11112 2388 11118 2440
rect 11238 2388 11244 2440
rect 11296 2428 11302 2440
rect 12728 2437 12756 2468
rect 13004 2437 13032 2536
rect 13078 2524 13084 2576
rect 13136 2564 13142 2576
rect 13136 2536 24440 2564
rect 13136 2524 13142 2536
rect 20714 2456 20720 2508
rect 20772 2456 20778 2508
rect 21174 2456 21180 2508
rect 21232 2496 21238 2508
rect 22281 2499 22339 2505
rect 22281 2496 22293 2499
rect 21232 2468 22293 2496
rect 21232 2456 21238 2468
rect 22281 2465 22293 2468
rect 22327 2465 22339 2499
rect 22281 2459 22339 2465
rect 11517 2431 11575 2437
rect 11517 2428 11529 2431
rect 11296 2400 11529 2428
rect 11296 2388 11302 2400
rect 11517 2397 11529 2400
rect 11563 2397 11575 2431
rect 11517 2391 11575 2397
rect 12161 2431 12219 2437
rect 12161 2397 12173 2431
rect 12207 2428 12219 2431
rect 12437 2431 12495 2437
rect 12437 2428 12449 2431
rect 12207 2400 12449 2428
rect 12207 2397 12219 2400
rect 12161 2391 12219 2397
rect 12437 2397 12449 2400
rect 12483 2397 12495 2431
rect 12437 2391 12495 2397
rect 12713 2431 12771 2437
rect 12713 2397 12725 2431
rect 12759 2397 12771 2431
rect 12713 2391 12771 2397
rect 12989 2431 13047 2437
rect 12989 2397 13001 2431
rect 13035 2397 13047 2431
rect 12989 2391 13047 2397
rect 13262 2388 13268 2440
rect 13320 2388 13326 2440
rect 17678 2388 17684 2440
rect 17736 2388 17742 2440
rect 20257 2431 20315 2437
rect 20257 2428 20269 2431
rect 20088 2400 20269 2428
rect 7650 2360 7656 2372
rect 7300 2332 7656 2360
rect 6641 2323 6699 2329
rect 7650 2320 7656 2332
rect 7708 2320 7714 2372
rect 5258 2292 5264 2304
rect 3712 2264 5264 2292
rect 5258 2252 5264 2264
rect 5316 2252 5322 2304
rect 5445 2295 5503 2301
rect 5445 2261 5457 2295
rect 5491 2292 5503 2295
rect 8938 2292 8944 2304
rect 5491 2264 8944 2292
rect 5491 2261 5503 2264
rect 5445 2255 5503 2261
rect 8938 2252 8944 2264
rect 8996 2252 9002 2304
rect 9861 2295 9919 2301
rect 9861 2261 9873 2295
rect 9907 2292 9919 2295
rect 11072 2292 11100 2388
rect 18874 2320 18880 2372
rect 18932 2320 18938 2372
rect 9907 2264 11100 2292
rect 9907 2261 9919 2264
rect 9861 2255 9919 2261
rect 11974 2252 11980 2304
rect 12032 2292 12038 2304
rect 12805 2295 12863 2301
rect 12805 2292 12817 2295
rect 12032 2264 12817 2292
rect 12032 2252 12038 2264
rect 12805 2261 12817 2264
rect 12851 2261 12863 2295
rect 12805 2255 12863 2261
rect 13078 2252 13084 2304
rect 13136 2252 13142 2304
rect 15194 2252 15200 2304
rect 15252 2292 15258 2304
rect 20088 2301 20116 2400
rect 20257 2397 20269 2400
rect 20303 2397 20315 2431
rect 20257 2391 20315 2397
rect 20346 2388 20352 2440
rect 20404 2428 20410 2440
rect 24412 2437 24440 2536
rect 24578 2456 24584 2508
rect 24636 2496 24642 2508
rect 24857 2499 24915 2505
rect 24857 2496 24869 2499
rect 24636 2468 24869 2496
rect 24636 2456 24642 2468
rect 24857 2465 24869 2468
rect 24903 2465 24915 2499
rect 27433 2499 27491 2505
rect 27433 2496 27445 2499
rect 24857 2459 24915 2465
rect 25240 2468 27445 2496
rect 21821 2431 21879 2437
rect 21821 2428 21833 2431
rect 20404 2400 21833 2428
rect 20404 2388 20410 2400
rect 21821 2397 21833 2400
rect 21867 2397 21879 2431
rect 21821 2391 21879 2397
rect 24397 2431 24455 2437
rect 24397 2397 24409 2431
rect 24443 2397 24455 2431
rect 24397 2391 24455 2397
rect 23382 2320 23388 2372
rect 23440 2360 23446 2372
rect 25240 2360 25268 2468
rect 27433 2465 27445 2468
rect 27479 2465 27491 2499
rect 27433 2459 27491 2465
rect 26973 2431 27031 2437
rect 26973 2397 26985 2431
rect 27019 2397 27031 2431
rect 26973 2391 27031 2397
rect 23440 2332 25268 2360
rect 23440 2320 23446 2332
rect 20073 2295 20131 2301
rect 20073 2292 20085 2295
rect 15252 2264 20085 2292
rect 15252 2252 15258 2264
rect 20073 2261 20085 2264
rect 20119 2261 20131 2295
rect 20073 2255 20131 2261
rect 26234 2252 26240 2304
rect 26292 2292 26298 2304
rect 26697 2295 26755 2301
rect 26697 2292 26709 2295
rect 26292 2264 26709 2292
rect 26292 2252 26298 2264
rect 26697 2261 26709 2264
rect 26743 2292 26755 2295
rect 26988 2292 27016 2391
rect 26743 2264 27016 2292
rect 26743 2261 26755 2264
rect 26697 2255 26755 2261
rect 1104 2202 29048 2224
rect 1104 2150 7896 2202
rect 7948 2150 7960 2202
rect 8012 2150 8024 2202
rect 8076 2150 8088 2202
rect 8140 2150 8152 2202
rect 8204 2150 14842 2202
rect 14894 2150 14906 2202
rect 14958 2150 14970 2202
rect 15022 2150 15034 2202
rect 15086 2150 15098 2202
rect 15150 2150 21788 2202
rect 21840 2150 21852 2202
rect 21904 2150 21916 2202
rect 21968 2150 21980 2202
rect 22032 2150 22044 2202
rect 22096 2150 28734 2202
rect 28786 2150 28798 2202
rect 28850 2150 28862 2202
rect 28914 2150 28926 2202
rect 28978 2150 28990 2202
rect 29042 2150 29048 2202
rect 1104 2128 29048 2150
rect 5350 2048 5356 2100
rect 5408 2088 5414 2100
rect 6546 2088 6552 2100
rect 5408 2060 6552 2088
rect 5408 2048 5414 2060
rect 6546 2048 6552 2060
rect 6604 2048 6610 2100
rect 13078 2048 13084 2100
rect 13136 2048 13142 2100
rect 18874 2048 18880 2100
rect 18932 2088 18938 2100
rect 18932 2060 24854 2088
rect 18932 2048 18938 2060
rect 3050 1980 3056 2032
rect 3108 2020 3114 2032
rect 5994 2020 6000 2032
rect 3108 1992 6000 2020
rect 3108 1980 3114 1992
rect 5994 1980 6000 1992
rect 6052 1980 6058 2032
rect 6178 1980 6184 2032
rect 6236 2020 6242 2032
rect 10870 2020 10876 2032
rect 6236 1992 10876 2020
rect 6236 1980 6242 1992
rect 10870 1980 10876 1992
rect 10928 1980 10934 2032
rect 2314 1912 2320 1964
rect 2372 1952 2378 1964
rect 5718 1952 5724 1964
rect 2372 1924 5724 1952
rect 2372 1912 2378 1924
rect 5718 1912 5724 1924
rect 5776 1912 5782 1964
rect 2406 1844 2412 1896
rect 2464 1884 2470 1896
rect 13096 1884 13124 2048
rect 24826 2020 24854 2060
rect 25590 2048 25596 2100
rect 25648 2088 25654 2100
rect 26418 2088 26424 2100
rect 25648 2060 26424 2088
rect 25648 2048 25654 2060
rect 26418 2048 26424 2060
rect 26476 2048 26482 2100
rect 27246 2048 27252 2100
rect 27304 2088 27310 2100
rect 27798 2088 27804 2100
rect 27304 2060 27804 2088
rect 27304 2048 27310 2060
rect 27798 2048 27804 2060
rect 27856 2048 27862 2100
rect 28902 2020 28908 2032
rect 24826 1992 28908 2020
rect 28902 1980 28908 1992
rect 28960 1980 28966 2032
rect 14642 1912 14648 1964
rect 14700 1952 14706 1964
rect 26234 1952 26240 1964
rect 14700 1924 26240 1952
rect 14700 1912 14706 1924
rect 26234 1912 26240 1924
rect 26292 1912 26298 1964
rect 2464 1856 13124 1884
rect 2464 1844 2470 1856
rect 24854 1844 24860 1896
rect 24912 1884 24918 1896
rect 26418 1884 26424 1896
rect 24912 1856 26424 1884
rect 24912 1844 24918 1856
rect 26418 1844 26424 1856
rect 26476 1844 26482 1896
rect 3602 1776 3608 1828
rect 3660 1776 3666 1828
rect 3620 1748 3648 1776
rect 10962 1748 10968 1760
rect 3620 1720 10968 1748
rect 10962 1708 10968 1720
rect 11020 1708 11026 1760
rect 2130 1640 2136 1692
rect 2188 1680 2194 1692
rect 8662 1680 8668 1692
rect 2188 1652 8668 1680
rect 2188 1640 2194 1652
rect 8662 1640 8668 1652
rect 8720 1640 8726 1692
rect 2866 1504 2872 1556
rect 2924 1544 2930 1556
rect 11146 1544 11152 1556
rect 2924 1516 11152 1544
rect 2924 1504 2930 1516
rect 11146 1504 11152 1516
rect 11204 1504 11210 1556
rect 24578 1504 24584 1556
rect 24636 1504 24642 1556
rect 22002 1368 22008 1420
rect 22060 1408 22066 1420
rect 24596 1408 24624 1504
rect 22060 1380 24624 1408
rect 22060 1368 22066 1380
<< via1 >>
rect 4423 27718 4475 27770
rect 4487 27718 4539 27770
rect 4551 27718 4603 27770
rect 4615 27718 4667 27770
rect 4679 27718 4731 27770
rect 11369 27718 11421 27770
rect 11433 27718 11485 27770
rect 11497 27718 11549 27770
rect 11561 27718 11613 27770
rect 11625 27718 11677 27770
rect 18315 27718 18367 27770
rect 18379 27718 18431 27770
rect 18443 27718 18495 27770
rect 18507 27718 18559 27770
rect 18571 27718 18623 27770
rect 25261 27718 25313 27770
rect 25325 27718 25377 27770
rect 25389 27718 25441 27770
rect 25453 27718 25505 27770
rect 25517 27718 25569 27770
rect 28540 27523 28592 27532
rect 28540 27489 28549 27523
rect 28549 27489 28583 27523
rect 28583 27489 28592 27523
rect 28540 27480 28592 27489
rect 7896 27174 7948 27226
rect 7960 27174 8012 27226
rect 8024 27174 8076 27226
rect 8088 27174 8140 27226
rect 8152 27174 8204 27226
rect 14842 27174 14894 27226
rect 14906 27174 14958 27226
rect 14970 27174 15022 27226
rect 15034 27174 15086 27226
rect 15098 27174 15150 27226
rect 21788 27174 21840 27226
rect 21852 27174 21904 27226
rect 21916 27174 21968 27226
rect 21980 27174 22032 27226
rect 22044 27174 22096 27226
rect 28734 27174 28786 27226
rect 28798 27174 28850 27226
rect 28862 27174 28914 27226
rect 28926 27174 28978 27226
rect 28990 27174 29042 27226
rect 22744 26732 22796 26784
rect 28356 26911 28408 26920
rect 28356 26877 28365 26911
rect 28365 26877 28399 26911
rect 28399 26877 28408 26911
rect 28356 26868 28408 26877
rect 4423 26630 4475 26682
rect 4487 26630 4539 26682
rect 4551 26630 4603 26682
rect 4615 26630 4667 26682
rect 4679 26630 4731 26682
rect 11369 26630 11421 26682
rect 11433 26630 11485 26682
rect 11497 26630 11549 26682
rect 11561 26630 11613 26682
rect 11625 26630 11677 26682
rect 18315 26630 18367 26682
rect 18379 26630 18431 26682
rect 18443 26630 18495 26682
rect 18507 26630 18559 26682
rect 18571 26630 18623 26682
rect 25261 26630 25313 26682
rect 25325 26630 25377 26682
rect 25389 26630 25441 26682
rect 25453 26630 25505 26682
rect 25517 26630 25569 26682
rect 14280 26256 14332 26308
rect 28356 26299 28408 26308
rect 28356 26265 28365 26299
rect 28365 26265 28399 26299
rect 28399 26265 28408 26299
rect 28356 26256 28408 26265
rect 7896 26086 7948 26138
rect 7960 26086 8012 26138
rect 8024 26086 8076 26138
rect 8088 26086 8140 26138
rect 8152 26086 8204 26138
rect 14842 26086 14894 26138
rect 14906 26086 14958 26138
rect 14970 26086 15022 26138
rect 15034 26086 15086 26138
rect 15098 26086 15150 26138
rect 21788 26086 21840 26138
rect 21852 26086 21904 26138
rect 21916 26086 21968 26138
rect 21980 26086 22032 26138
rect 22044 26086 22096 26138
rect 28734 26086 28786 26138
rect 28798 26086 28850 26138
rect 28862 26086 28914 26138
rect 28926 26086 28978 26138
rect 28990 26086 29042 26138
rect 4423 25542 4475 25594
rect 4487 25542 4539 25594
rect 4551 25542 4603 25594
rect 4615 25542 4667 25594
rect 4679 25542 4731 25594
rect 11369 25542 11421 25594
rect 11433 25542 11485 25594
rect 11497 25542 11549 25594
rect 11561 25542 11613 25594
rect 11625 25542 11677 25594
rect 18315 25542 18367 25594
rect 18379 25542 18431 25594
rect 18443 25542 18495 25594
rect 18507 25542 18559 25594
rect 18571 25542 18623 25594
rect 25261 25542 25313 25594
rect 25325 25542 25377 25594
rect 25389 25542 25441 25594
rect 25453 25542 25505 25594
rect 25517 25542 25569 25594
rect 25688 25100 25740 25152
rect 28356 25211 28408 25220
rect 28356 25177 28365 25211
rect 28365 25177 28399 25211
rect 28399 25177 28408 25211
rect 28356 25168 28408 25177
rect 7896 24998 7948 25050
rect 7960 24998 8012 25050
rect 8024 24998 8076 25050
rect 8088 24998 8140 25050
rect 8152 24998 8204 25050
rect 14842 24998 14894 25050
rect 14906 24998 14958 25050
rect 14970 24998 15022 25050
rect 15034 24998 15086 25050
rect 15098 24998 15150 25050
rect 21788 24998 21840 25050
rect 21852 24998 21904 25050
rect 21916 24998 21968 25050
rect 21980 24998 22032 25050
rect 22044 24998 22096 25050
rect 28734 24998 28786 25050
rect 28798 24998 28850 25050
rect 28862 24998 28914 25050
rect 28926 24998 28978 25050
rect 28990 24998 29042 25050
rect 12808 24556 12860 24608
rect 28356 24735 28408 24744
rect 28356 24701 28365 24735
rect 28365 24701 28399 24735
rect 28399 24701 28408 24735
rect 28356 24692 28408 24701
rect 4423 24454 4475 24506
rect 4487 24454 4539 24506
rect 4551 24454 4603 24506
rect 4615 24454 4667 24506
rect 4679 24454 4731 24506
rect 11369 24454 11421 24506
rect 11433 24454 11485 24506
rect 11497 24454 11549 24506
rect 11561 24454 11613 24506
rect 11625 24454 11677 24506
rect 18315 24454 18367 24506
rect 18379 24454 18431 24506
rect 18443 24454 18495 24506
rect 18507 24454 18559 24506
rect 18571 24454 18623 24506
rect 25261 24454 25313 24506
rect 25325 24454 25377 24506
rect 25389 24454 25441 24506
rect 25453 24454 25505 24506
rect 25517 24454 25569 24506
rect 7896 23910 7948 23962
rect 7960 23910 8012 23962
rect 8024 23910 8076 23962
rect 8088 23910 8140 23962
rect 8152 23910 8204 23962
rect 14842 23910 14894 23962
rect 14906 23910 14958 23962
rect 14970 23910 15022 23962
rect 15034 23910 15086 23962
rect 15098 23910 15150 23962
rect 21788 23910 21840 23962
rect 21852 23910 21904 23962
rect 21916 23910 21968 23962
rect 21980 23910 22032 23962
rect 22044 23910 22096 23962
rect 28734 23910 28786 23962
rect 28798 23910 28850 23962
rect 28862 23910 28914 23962
rect 28926 23910 28978 23962
rect 28990 23910 29042 23962
rect 1400 23715 1452 23724
rect 1400 23681 1409 23715
rect 1409 23681 1443 23715
rect 1443 23681 1452 23715
rect 1400 23672 1452 23681
rect 1584 23511 1636 23520
rect 1584 23477 1593 23511
rect 1593 23477 1627 23511
rect 1627 23477 1636 23511
rect 1584 23468 1636 23477
rect 25780 23468 25832 23520
rect 28724 23604 28776 23656
rect 4423 23366 4475 23418
rect 4487 23366 4539 23418
rect 4551 23366 4603 23418
rect 4615 23366 4667 23418
rect 4679 23366 4731 23418
rect 11369 23366 11421 23418
rect 11433 23366 11485 23418
rect 11497 23366 11549 23418
rect 11561 23366 11613 23418
rect 11625 23366 11677 23418
rect 18315 23366 18367 23418
rect 18379 23366 18431 23418
rect 18443 23366 18495 23418
rect 18507 23366 18559 23418
rect 18571 23366 18623 23418
rect 25261 23366 25313 23418
rect 25325 23366 25377 23418
rect 25389 23366 25441 23418
rect 25453 23366 25505 23418
rect 25517 23366 25569 23418
rect 4252 23196 4304 23248
rect 940 23060 992 23112
rect 1032 22992 1084 23044
rect 1860 22967 1912 22976
rect 1860 22933 1869 22967
rect 1869 22933 1903 22967
rect 1903 22933 1912 22967
rect 1860 22924 1912 22933
rect 16028 22924 16080 22976
rect 28356 23035 28408 23044
rect 28356 23001 28365 23035
rect 28365 23001 28399 23035
rect 28399 23001 28408 23035
rect 28356 22992 28408 23001
rect 7896 22822 7948 22874
rect 7960 22822 8012 22874
rect 8024 22822 8076 22874
rect 8088 22822 8140 22874
rect 8152 22822 8204 22874
rect 14842 22822 14894 22874
rect 14906 22822 14958 22874
rect 14970 22822 15022 22874
rect 15034 22822 15086 22874
rect 15098 22822 15150 22874
rect 21788 22822 21840 22874
rect 21852 22822 21904 22874
rect 21916 22822 21968 22874
rect 21980 22822 22032 22874
rect 22044 22822 22096 22874
rect 28734 22822 28786 22874
rect 28798 22822 28850 22874
rect 28862 22822 28914 22874
rect 28926 22822 28978 22874
rect 28990 22822 29042 22874
rect 1032 22584 1084 22636
rect 940 22516 992 22568
rect 2044 22448 2096 22500
rect 10232 22380 10284 22432
rect 4423 22278 4475 22330
rect 4487 22278 4539 22330
rect 4551 22278 4603 22330
rect 4615 22278 4667 22330
rect 4679 22278 4731 22330
rect 11369 22278 11421 22330
rect 11433 22278 11485 22330
rect 11497 22278 11549 22330
rect 11561 22278 11613 22330
rect 11625 22278 11677 22330
rect 18315 22278 18367 22330
rect 18379 22278 18431 22330
rect 18443 22278 18495 22330
rect 18507 22278 18559 22330
rect 18571 22278 18623 22330
rect 25261 22278 25313 22330
rect 25325 22278 25377 22330
rect 25389 22278 25441 22330
rect 25453 22278 25505 22330
rect 25517 22278 25569 22330
rect 28816 22040 28868 22092
rect 940 21972 992 22024
rect 1032 21904 1084 21956
rect 9220 21904 9272 21956
rect 9680 21836 9732 21888
rect 14648 21836 14700 21888
rect 7896 21734 7948 21786
rect 7960 21734 8012 21786
rect 8024 21734 8076 21786
rect 8088 21734 8140 21786
rect 8152 21734 8204 21786
rect 14842 21734 14894 21786
rect 14906 21734 14958 21786
rect 14970 21734 15022 21786
rect 15034 21734 15086 21786
rect 15098 21734 15150 21786
rect 21788 21734 21840 21786
rect 21852 21734 21904 21786
rect 21916 21734 21968 21786
rect 21980 21734 22032 21786
rect 22044 21734 22096 21786
rect 28734 21734 28786 21786
rect 28798 21734 28850 21786
rect 28862 21734 28914 21786
rect 28926 21734 28978 21786
rect 28990 21734 29042 21786
rect 1032 21496 1084 21548
rect 940 21428 992 21480
rect 15752 21496 15804 21548
rect 28356 21471 28408 21480
rect 28356 21437 28365 21471
rect 28365 21437 28399 21471
rect 28399 21437 28408 21471
rect 28356 21428 28408 21437
rect 7472 21360 7524 21412
rect 8392 21292 8444 21344
rect 4423 21190 4475 21242
rect 4487 21190 4539 21242
rect 4551 21190 4603 21242
rect 4615 21190 4667 21242
rect 4679 21190 4731 21242
rect 11369 21190 11421 21242
rect 11433 21190 11485 21242
rect 11497 21190 11549 21242
rect 11561 21190 11613 21242
rect 11625 21190 11677 21242
rect 18315 21190 18367 21242
rect 18379 21190 18431 21242
rect 18443 21190 18495 21242
rect 18507 21190 18559 21242
rect 18571 21190 18623 21242
rect 25261 21190 25313 21242
rect 25325 21190 25377 21242
rect 25389 21190 25441 21242
rect 25453 21190 25505 21242
rect 25517 21190 25569 21242
rect 4068 21020 4120 21072
rect 1400 20927 1452 20936
rect 1400 20893 1409 20927
rect 1409 20893 1443 20927
rect 1443 20893 1452 20927
rect 1400 20884 1452 20893
rect 940 20816 992 20868
rect 7656 20748 7708 20800
rect 7896 20646 7948 20698
rect 7960 20646 8012 20698
rect 8024 20646 8076 20698
rect 8088 20646 8140 20698
rect 8152 20646 8204 20698
rect 14842 20646 14894 20698
rect 14906 20646 14958 20698
rect 14970 20646 15022 20698
rect 15034 20646 15086 20698
rect 15098 20646 15150 20698
rect 21788 20646 21840 20698
rect 21852 20646 21904 20698
rect 21916 20646 21968 20698
rect 21980 20646 22032 20698
rect 22044 20646 22096 20698
rect 28734 20646 28786 20698
rect 28798 20646 28850 20698
rect 28862 20646 28914 20698
rect 28926 20646 28978 20698
rect 28990 20646 29042 20698
rect 940 20408 992 20460
rect 1032 20340 1084 20392
rect 1584 20247 1636 20256
rect 1584 20213 1593 20247
rect 1593 20213 1627 20247
rect 1627 20213 1636 20247
rect 1584 20204 1636 20213
rect 5540 20204 5592 20256
rect 16212 20204 16264 20256
rect 28356 20383 28408 20392
rect 28356 20349 28365 20383
rect 28365 20349 28399 20383
rect 28399 20349 28408 20383
rect 28356 20340 28408 20349
rect 4423 20102 4475 20154
rect 4487 20102 4539 20154
rect 4551 20102 4603 20154
rect 4615 20102 4667 20154
rect 4679 20102 4731 20154
rect 11369 20102 11421 20154
rect 11433 20102 11485 20154
rect 11497 20102 11549 20154
rect 11561 20102 11613 20154
rect 11625 20102 11677 20154
rect 18315 20102 18367 20154
rect 18379 20102 18431 20154
rect 18443 20102 18495 20154
rect 18507 20102 18559 20154
rect 18571 20102 18623 20154
rect 25261 20102 25313 20154
rect 25325 20102 25377 20154
rect 25389 20102 25441 20154
rect 25453 20102 25505 20154
rect 25517 20102 25569 20154
rect 5632 19932 5684 19984
rect 940 19796 992 19848
rect 1032 19728 1084 19780
rect 1860 19703 1912 19712
rect 1860 19669 1869 19703
rect 1869 19669 1903 19703
rect 1903 19669 1912 19703
rect 1860 19660 1912 19669
rect 10784 19660 10836 19712
rect 28356 19771 28408 19780
rect 28356 19737 28365 19771
rect 28365 19737 28399 19771
rect 28399 19737 28408 19771
rect 28356 19728 28408 19737
rect 7896 19558 7948 19610
rect 7960 19558 8012 19610
rect 8024 19558 8076 19610
rect 8088 19558 8140 19610
rect 8152 19558 8204 19610
rect 14842 19558 14894 19610
rect 14906 19558 14958 19610
rect 14970 19558 15022 19610
rect 15034 19558 15086 19610
rect 15098 19558 15150 19610
rect 21788 19558 21840 19610
rect 21852 19558 21904 19610
rect 21916 19558 21968 19610
rect 21980 19558 22032 19610
rect 22044 19558 22096 19610
rect 28734 19558 28786 19610
rect 28798 19558 28850 19610
rect 28862 19558 28914 19610
rect 28926 19558 28978 19610
rect 28990 19558 29042 19610
rect 3608 19456 3660 19508
rect 3976 19388 4028 19440
rect 1400 19363 1452 19372
rect 1400 19329 1409 19363
rect 1409 19329 1443 19363
rect 1443 19329 1452 19363
rect 1400 19320 1452 19329
rect 1676 19363 1728 19372
rect 1676 19329 1685 19363
rect 1685 19329 1719 19363
rect 1719 19329 1728 19363
rect 1676 19320 1728 19329
rect 4423 19014 4475 19066
rect 4487 19014 4539 19066
rect 4551 19014 4603 19066
rect 4615 19014 4667 19066
rect 4679 19014 4731 19066
rect 11369 19014 11421 19066
rect 11433 19014 11485 19066
rect 11497 19014 11549 19066
rect 11561 19014 11613 19066
rect 11625 19014 11677 19066
rect 18315 19014 18367 19066
rect 18379 19014 18431 19066
rect 18443 19014 18495 19066
rect 18507 19014 18559 19066
rect 18571 19014 18623 19066
rect 25261 19014 25313 19066
rect 25325 19014 25377 19066
rect 25389 19014 25441 19066
rect 25453 19014 25505 19066
rect 25517 19014 25569 19066
rect 12808 18955 12860 18964
rect 12808 18921 12817 18955
rect 12817 18921 12851 18955
rect 12851 18921 12860 18955
rect 12808 18912 12860 18921
rect 3332 18844 3384 18896
rect 28816 18776 28868 18828
rect 940 18708 992 18760
rect 1032 18640 1084 18692
rect 3792 18572 3844 18624
rect 17776 18572 17828 18624
rect 7896 18470 7948 18522
rect 7960 18470 8012 18522
rect 8024 18470 8076 18522
rect 8088 18470 8140 18522
rect 8152 18470 8204 18522
rect 14842 18470 14894 18522
rect 14906 18470 14958 18522
rect 14970 18470 15022 18522
rect 15034 18470 15086 18522
rect 15098 18470 15150 18522
rect 21788 18470 21840 18522
rect 21852 18470 21904 18522
rect 21916 18470 21968 18522
rect 21980 18470 22032 18522
rect 22044 18470 22096 18522
rect 28734 18470 28786 18522
rect 28798 18470 28850 18522
rect 28862 18470 28914 18522
rect 28926 18470 28978 18522
rect 28990 18470 29042 18522
rect 12808 18368 12860 18420
rect 13728 18368 13780 18420
rect 8300 18300 8352 18352
rect 1400 18275 1452 18284
rect 1400 18241 1409 18275
rect 1409 18241 1443 18275
rect 1443 18241 1452 18275
rect 1400 18232 1452 18241
rect 940 18164 992 18216
rect 9220 18275 9272 18284
rect 9220 18241 9229 18275
rect 9229 18241 9263 18275
rect 9263 18241 9272 18275
rect 9220 18232 9272 18241
rect 9404 18275 9456 18284
rect 9404 18241 9413 18275
rect 9413 18241 9447 18275
rect 9447 18241 9456 18275
rect 9404 18232 9456 18241
rect 9680 18275 9732 18284
rect 9680 18241 9689 18275
rect 9689 18241 9723 18275
rect 9723 18241 9732 18275
rect 9680 18232 9732 18241
rect 9864 18275 9916 18284
rect 9864 18241 9873 18275
rect 9873 18241 9907 18275
rect 9907 18241 9916 18275
rect 9864 18232 9916 18241
rect 10600 18232 10652 18284
rect 4252 18164 4304 18216
rect 10140 18164 10192 18216
rect 10508 18164 10560 18216
rect 3424 18096 3476 18148
rect 10876 18096 10928 18148
rect 28356 18207 28408 18216
rect 28356 18173 28365 18207
rect 28365 18173 28399 18207
rect 28399 18173 28408 18207
rect 28356 18164 28408 18173
rect 4160 18028 4212 18080
rect 10048 18071 10100 18080
rect 10048 18037 10057 18071
rect 10057 18037 10091 18071
rect 10091 18037 10100 18071
rect 10048 18028 10100 18037
rect 12716 18071 12768 18080
rect 12716 18037 12725 18071
rect 12725 18037 12759 18071
rect 12759 18037 12768 18071
rect 12716 18028 12768 18037
rect 4423 17926 4475 17978
rect 4487 17926 4539 17978
rect 4551 17926 4603 17978
rect 4615 17926 4667 17978
rect 4679 17926 4731 17978
rect 11369 17926 11421 17978
rect 11433 17926 11485 17978
rect 11497 17926 11549 17978
rect 11561 17926 11613 17978
rect 11625 17926 11677 17978
rect 18315 17926 18367 17978
rect 18379 17926 18431 17978
rect 18443 17926 18495 17978
rect 18507 17926 18559 17978
rect 18571 17926 18623 17978
rect 25261 17926 25313 17978
rect 25325 17926 25377 17978
rect 25389 17926 25441 17978
rect 25453 17926 25505 17978
rect 25517 17926 25569 17978
rect 10600 17867 10652 17876
rect 10600 17833 10609 17867
rect 10609 17833 10643 17867
rect 10643 17833 10652 17867
rect 10600 17824 10652 17833
rect 3700 17756 3752 17808
rect 9772 17756 9824 17808
rect 10784 17756 10836 17808
rect 10232 17731 10284 17740
rect 10232 17697 10241 17731
rect 10241 17697 10275 17731
rect 10275 17697 10284 17731
rect 10232 17688 10284 17697
rect 11704 17688 11756 17740
rect 11796 17688 11848 17740
rect 16028 17688 16080 17740
rect 1032 17620 1084 17672
rect 940 17552 992 17604
rect 9864 17663 9916 17672
rect 9864 17629 9873 17663
rect 9873 17629 9907 17663
rect 9907 17629 9916 17663
rect 9864 17620 9916 17629
rect 10416 17663 10468 17672
rect 10416 17629 10425 17663
rect 10425 17629 10459 17663
rect 10459 17629 10468 17663
rect 10416 17620 10468 17629
rect 10692 17663 10744 17672
rect 10692 17629 10701 17663
rect 10701 17629 10735 17663
rect 10735 17629 10744 17663
rect 10692 17620 10744 17629
rect 13176 17552 13228 17604
rect 3516 17484 3568 17536
rect 8760 17484 8812 17536
rect 9312 17527 9364 17536
rect 9312 17493 9321 17527
rect 9321 17493 9355 17527
rect 9355 17493 9364 17527
rect 9312 17484 9364 17493
rect 7896 17382 7948 17434
rect 7960 17382 8012 17434
rect 8024 17382 8076 17434
rect 8088 17382 8140 17434
rect 8152 17382 8204 17434
rect 14842 17382 14894 17434
rect 14906 17382 14958 17434
rect 14970 17382 15022 17434
rect 15034 17382 15086 17434
rect 15098 17382 15150 17434
rect 21788 17382 21840 17434
rect 21852 17382 21904 17434
rect 21916 17382 21968 17434
rect 21980 17382 22032 17434
rect 22044 17382 22096 17434
rect 28734 17382 28786 17434
rect 28798 17382 28850 17434
rect 28862 17382 28914 17434
rect 28926 17382 28978 17434
rect 28990 17382 29042 17434
rect 5264 17280 5316 17332
rect 8852 17280 8904 17332
rect 9864 17280 9916 17332
rect 10048 17323 10100 17332
rect 10048 17289 10057 17323
rect 10057 17289 10091 17323
rect 10091 17289 10100 17323
rect 10048 17280 10100 17289
rect 10692 17280 10744 17332
rect 10876 17323 10928 17332
rect 10876 17289 10885 17323
rect 10885 17289 10919 17323
rect 10919 17289 10928 17323
rect 10876 17280 10928 17289
rect 11796 17280 11848 17332
rect 1860 17212 1912 17264
rect 12716 17280 12768 17332
rect 940 17144 992 17196
rect 1032 17076 1084 17128
rect 5540 17144 5592 17196
rect 7196 17119 7248 17128
rect 7196 17085 7205 17119
rect 7205 17085 7239 17119
rect 7239 17085 7248 17119
rect 7196 17076 7248 17085
rect 7380 17144 7432 17196
rect 7656 17144 7708 17196
rect 1308 17008 1360 17060
rect 7564 17008 7616 17060
rect 9772 17144 9824 17196
rect 10968 17187 11020 17196
rect 10968 17153 10977 17187
rect 10977 17153 11011 17187
rect 11011 17153 11020 17187
rect 10968 17144 11020 17153
rect 13728 17187 13780 17196
rect 13728 17153 13737 17187
rect 13737 17153 13771 17187
rect 13771 17153 13780 17187
rect 13728 17144 13780 17153
rect 14740 17187 14792 17196
rect 14740 17153 14749 17187
rect 14749 17153 14783 17187
rect 14783 17153 14792 17187
rect 14740 17144 14792 17153
rect 16580 17144 16632 17196
rect 8760 17119 8812 17128
rect 8760 17085 8769 17119
rect 8769 17085 8803 17119
rect 8803 17085 8812 17119
rect 8760 17076 8812 17085
rect 6460 16940 6512 16992
rect 7380 16983 7432 16992
rect 7380 16949 7389 16983
rect 7389 16949 7423 16983
rect 7423 16949 7432 16983
rect 7380 16940 7432 16949
rect 7748 16940 7800 16992
rect 10508 17076 10560 17128
rect 11152 17076 11204 17128
rect 11704 17119 11756 17128
rect 11704 17085 11713 17119
rect 11713 17085 11747 17119
rect 11747 17085 11756 17119
rect 11704 17076 11756 17085
rect 28356 17119 28408 17128
rect 28356 17085 28365 17119
rect 28365 17085 28399 17119
rect 28399 17085 28408 17119
rect 28356 17076 28408 17085
rect 13820 16983 13872 16992
rect 13820 16949 13829 16983
rect 13829 16949 13863 16983
rect 13863 16949 13872 16983
rect 13820 16940 13872 16949
rect 4423 16838 4475 16890
rect 4487 16838 4539 16890
rect 4551 16838 4603 16890
rect 4615 16838 4667 16890
rect 4679 16838 4731 16890
rect 11369 16838 11421 16890
rect 11433 16838 11485 16890
rect 11497 16838 11549 16890
rect 11561 16838 11613 16890
rect 11625 16838 11677 16890
rect 18315 16838 18367 16890
rect 18379 16838 18431 16890
rect 18443 16838 18495 16890
rect 18507 16838 18559 16890
rect 18571 16838 18623 16890
rect 25261 16838 25313 16890
rect 25325 16838 25377 16890
rect 25389 16838 25441 16890
rect 25453 16838 25505 16890
rect 25517 16838 25569 16890
rect 10968 16736 11020 16788
rect 13636 16736 13688 16788
rect 13820 16736 13872 16788
rect 11060 16668 11112 16720
rect 6460 16600 6512 16652
rect 8300 16600 8352 16652
rect 8392 16643 8444 16652
rect 8392 16609 8401 16643
rect 8401 16609 8435 16643
rect 8435 16609 8444 16643
rect 8392 16600 8444 16609
rect 9312 16600 9364 16652
rect 10784 16600 10836 16652
rect 940 16532 992 16584
rect 1032 16464 1084 16516
rect 5724 16532 5776 16584
rect 664 16396 716 16448
rect 1676 16439 1728 16448
rect 1676 16405 1685 16439
rect 1685 16405 1719 16439
rect 1719 16405 1728 16439
rect 1676 16396 1728 16405
rect 8576 16575 8628 16584
rect 8576 16541 8585 16575
rect 8585 16541 8619 16575
rect 8619 16541 8628 16575
rect 8576 16532 8628 16541
rect 6644 16464 6696 16516
rect 9864 16464 9916 16516
rect 11704 16575 11756 16584
rect 11704 16541 11713 16575
rect 11713 16541 11747 16575
rect 11747 16541 11756 16575
rect 11704 16532 11756 16541
rect 13636 16532 13688 16584
rect 14648 16532 14700 16584
rect 23480 16532 23532 16584
rect 13268 16464 13320 16516
rect 28356 16507 28408 16516
rect 28356 16473 28365 16507
rect 28365 16473 28399 16507
rect 28399 16473 28408 16507
rect 28356 16464 28408 16473
rect 8300 16396 8352 16448
rect 11336 16396 11388 16448
rect 11520 16439 11572 16448
rect 11520 16405 11529 16439
rect 11529 16405 11563 16439
rect 11563 16405 11572 16439
rect 11520 16396 11572 16405
rect 7896 16294 7948 16346
rect 7960 16294 8012 16346
rect 8024 16294 8076 16346
rect 8088 16294 8140 16346
rect 8152 16294 8204 16346
rect 14842 16294 14894 16346
rect 14906 16294 14958 16346
rect 14970 16294 15022 16346
rect 15034 16294 15086 16346
rect 15098 16294 15150 16346
rect 21788 16294 21840 16346
rect 21852 16294 21904 16346
rect 21916 16294 21968 16346
rect 21980 16294 22032 16346
rect 22044 16294 22096 16346
rect 28734 16294 28786 16346
rect 28798 16294 28850 16346
rect 28862 16294 28914 16346
rect 28926 16294 28978 16346
rect 28990 16294 29042 16346
rect 388 16192 440 16244
rect 1676 16192 1728 16244
rect 6644 16235 6696 16244
rect 6644 16201 6653 16235
rect 6653 16201 6687 16235
rect 6687 16201 6696 16235
rect 6644 16192 6696 16201
rect 7196 16192 7248 16244
rect 7380 16192 7432 16244
rect 8392 16192 8444 16244
rect 11520 16192 11572 16244
rect 940 16056 992 16108
rect 1032 15988 1084 16040
rect 7012 15988 7064 16040
rect 8300 16099 8352 16108
rect 8300 16065 8309 16099
rect 8309 16065 8343 16099
rect 8343 16065 8352 16099
rect 8300 16056 8352 16065
rect 11336 16099 11388 16108
rect 11336 16065 11345 16099
rect 11345 16065 11379 16099
rect 11379 16065 11388 16099
rect 11336 16056 11388 16065
rect 11704 16124 11756 16176
rect 13268 16192 13320 16244
rect 13084 16124 13136 16176
rect 15200 16124 15252 16176
rect 15752 16124 15804 16176
rect 7380 16031 7432 16040
rect 7380 15997 7389 16031
rect 7389 15997 7423 16031
rect 7423 15997 7432 16031
rect 7380 15988 7432 15997
rect 7472 15988 7524 16040
rect 7656 15920 7708 15972
rect 7748 15920 7800 15972
rect 10324 16031 10376 16040
rect 10324 15997 10333 16031
rect 10333 15997 10367 16031
rect 10367 15997 10376 16031
rect 10324 15988 10376 15997
rect 10968 16031 11020 16040
rect 10968 15997 10977 16031
rect 10977 15997 11011 16031
rect 11011 15997 11020 16031
rect 10968 15988 11020 15997
rect 1676 15852 1728 15904
rect 3240 15852 3292 15904
rect 7380 15852 7432 15904
rect 8208 15895 8260 15904
rect 8208 15861 8217 15895
rect 8217 15861 8251 15895
rect 8251 15861 8260 15895
rect 8208 15852 8260 15861
rect 9680 15852 9732 15904
rect 11796 16031 11848 16040
rect 11796 15997 11805 16031
rect 11805 15997 11839 16031
rect 11839 15997 11848 16031
rect 11796 15988 11848 15997
rect 13268 15852 13320 15904
rect 4423 15750 4475 15802
rect 4487 15750 4539 15802
rect 4551 15750 4603 15802
rect 4615 15750 4667 15802
rect 4679 15750 4731 15802
rect 11369 15750 11421 15802
rect 11433 15750 11485 15802
rect 11497 15750 11549 15802
rect 11561 15750 11613 15802
rect 11625 15750 11677 15802
rect 18315 15750 18367 15802
rect 18379 15750 18431 15802
rect 18443 15750 18495 15802
rect 18507 15750 18559 15802
rect 18571 15750 18623 15802
rect 25261 15750 25313 15802
rect 25325 15750 25377 15802
rect 25389 15750 25441 15802
rect 25453 15750 25505 15802
rect 25517 15750 25569 15802
rect 8208 15648 8260 15700
rect 9864 15691 9916 15700
rect 9864 15657 9873 15691
rect 9873 15657 9907 15691
rect 9907 15657 9916 15691
rect 9864 15648 9916 15657
rect 10968 15648 11020 15700
rect 11152 15648 11204 15700
rect 11796 15648 11848 15700
rect 13084 15648 13136 15700
rect 13176 15648 13228 15700
rect 14280 15691 14332 15700
rect 14280 15657 14289 15691
rect 14289 15657 14323 15691
rect 14323 15657 14332 15691
rect 14280 15648 14332 15657
rect 940 15580 992 15632
rect 8392 15512 8444 15564
rect 940 15444 992 15496
rect 1584 15444 1636 15496
rect 1860 15487 1912 15496
rect 1860 15453 1869 15487
rect 1869 15453 1903 15487
rect 1903 15453 1912 15487
rect 1860 15444 1912 15453
rect 7748 15376 7800 15428
rect 11060 15512 11112 15564
rect 12256 15512 12308 15564
rect 13268 15580 13320 15632
rect 9680 15376 9732 15428
rect 13268 15487 13320 15496
rect 13268 15453 13277 15487
rect 13277 15453 13311 15487
rect 13311 15453 13320 15487
rect 13268 15444 13320 15453
rect 480 15308 532 15360
rect 8760 15351 8812 15360
rect 8760 15317 8769 15351
rect 8769 15317 8803 15351
rect 8803 15317 8812 15351
rect 8760 15308 8812 15317
rect 10324 15351 10376 15360
rect 10324 15317 10333 15351
rect 10333 15317 10367 15351
rect 10367 15317 10376 15351
rect 16212 15376 16264 15428
rect 10324 15308 10376 15317
rect 12348 15308 12400 15360
rect 26976 15351 27028 15360
rect 26976 15317 26985 15351
rect 26985 15317 27019 15351
rect 27019 15317 27028 15351
rect 28356 15419 28408 15428
rect 28356 15385 28365 15419
rect 28365 15385 28399 15419
rect 28399 15385 28408 15419
rect 28356 15376 28408 15385
rect 26976 15308 27028 15317
rect 7896 15206 7948 15258
rect 7960 15206 8012 15258
rect 8024 15206 8076 15258
rect 8088 15206 8140 15258
rect 8152 15206 8204 15258
rect 14842 15206 14894 15258
rect 14906 15206 14958 15258
rect 14970 15206 15022 15258
rect 15034 15206 15086 15258
rect 15098 15206 15150 15258
rect 21788 15206 21840 15258
rect 21852 15206 21904 15258
rect 21916 15206 21968 15258
rect 21980 15206 22032 15258
rect 22044 15206 22096 15258
rect 28734 15206 28786 15258
rect 28798 15206 28850 15258
rect 28862 15206 28914 15258
rect 28926 15206 28978 15258
rect 28990 15206 29042 15258
rect 1768 15036 1820 15088
rect 940 14968 992 15020
rect 5632 14968 5684 15020
rect 6920 14943 6972 14952
rect 6920 14909 6929 14943
rect 6929 14909 6963 14943
rect 6963 14909 6972 14943
rect 6920 14900 6972 14909
rect 7288 15011 7340 15020
rect 7288 14977 7297 15011
rect 7297 14977 7331 15011
rect 7331 14977 7340 15011
rect 7288 14968 7340 14977
rect 7656 14968 7708 15020
rect 9680 14968 9732 15020
rect 11888 15036 11940 15088
rect 13268 15104 13320 15156
rect 14280 15104 14332 15156
rect 14740 15104 14792 15156
rect 12256 14943 12308 14952
rect 12256 14909 12265 14943
rect 12265 14909 12299 14943
rect 12299 14909 12308 14943
rect 12256 14900 12308 14909
rect 1584 14832 1636 14884
rect 6276 14764 6328 14816
rect 7104 14807 7156 14816
rect 7104 14773 7113 14807
rect 7113 14773 7147 14807
rect 7147 14773 7156 14807
rect 7104 14764 7156 14773
rect 7656 14807 7708 14816
rect 7656 14773 7665 14807
rect 7665 14773 7699 14807
rect 7699 14773 7708 14807
rect 7656 14764 7708 14773
rect 9772 14832 9824 14884
rect 10968 14832 11020 14884
rect 13728 14968 13780 15020
rect 14740 14968 14792 15020
rect 15292 14900 15344 14952
rect 13544 14832 13596 14884
rect 13728 14807 13780 14816
rect 13728 14773 13737 14807
rect 13737 14773 13771 14807
rect 13771 14773 13780 14807
rect 13728 14764 13780 14773
rect 14188 14807 14240 14816
rect 14188 14773 14197 14807
rect 14197 14773 14231 14807
rect 14231 14773 14240 14807
rect 14188 14764 14240 14773
rect 15476 14764 15528 14816
rect 15752 14764 15804 14816
rect 15936 14764 15988 14816
rect 28356 14943 28408 14952
rect 28356 14909 28365 14943
rect 28365 14909 28399 14943
rect 28399 14909 28408 14943
rect 28356 14900 28408 14909
rect 4423 14662 4475 14714
rect 4487 14662 4539 14714
rect 4551 14662 4603 14714
rect 4615 14662 4667 14714
rect 4679 14662 4731 14714
rect 11369 14662 11421 14714
rect 11433 14662 11485 14714
rect 11497 14662 11549 14714
rect 11561 14662 11613 14714
rect 11625 14662 11677 14714
rect 18315 14662 18367 14714
rect 18379 14662 18431 14714
rect 18443 14662 18495 14714
rect 18507 14662 18559 14714
rect 18571 14662 18623 14714
rect 25261 14662 25313 14714
rect 25325 14662 25377 14714
rect 25389 14662 25441 14714
rect 25453 14662 25505 14714
rect 25517 14662 25569 14714
rect 8300 14560 8352 14612
rect 6276 14424 6328 14476
rect 9772 14424 9824 14476
rect 940 14356 992 14408
rect 1032 14288 1084 14340
rect 5724 14356 5776 14408
rect 7656 14356 7708 14408
rect 9680 14356 9732 14408
rect 10324 14356 10376 14408
rect 10416 14399 10468 14408
rect 10416 14365 10425 14399
rect 10425 14365 10459 14399
rect 10459 14365 10468 14399
rect 10416 14356 10468 14365
rect 7472 14288 7524 14340
rect 10784 14399 10836 14408
rect 10784 14365 10793 14399
rect 10793 14365 10827 14399
rect 10827 14365 10836 14399
rect 10784 14356 10836 14365
rect 10968 14399 11020 14408
rect 10968 14365 10977 14399
rect 10977 14365 11011 14399
rect 11011 14365 11020 14399
rect 10968 14356 11020 14365
rect 11888 14560 11940 14612
rect 12348 14560 12400 14612
rect 13728 14560 13780 14612
rect 14188 14492 14240 14544
rect 11244 14399 11296 14408
rect 11244 14365 11253 14399
rect 11253 14365 11287 14399
rect 11287 14365 11296 14399
rect 11244 14356 11296 14365
rect 11888 14399 11940 14408
rect 11888 14365 11897 14399
rect 11897 14365 11931 14399
rect 11931 14365 11940 14399
rect 11888 14356 11940 14365
rect 13176 14356 13228 14408
rect 14740 14424 14792 14476
rect 1860 14263 1912 14272
rect 1860 14229 1869 14263
rect 1869 14229 1903 14263
rect 1903 14229 1912 14263
rect 1860 14220 1912 14229
rect 1952 14220 2004 14272
rect 13544 14288 13596 14340
rect 22744 14424 22796 14476
rect 15752 14399 15804 14408
rect 15752 14365 15761 14399
rect 15761 14365 15795 14399
rect 15795 14365 15804 14399
rect 15752 14356 15804 14365
rect 9772 14220 9824 14272
rect 12348 14220 12400 14272
rect 12440 14220 12492 14272
rect 14188 14220 14240 14272
rect 16304 14220 16356 14272
rect 7896 14118 7948 14170
rect 7960 14118 8012 14170
rect 8024 14118 8076 14170
rect 8088 14118 8140 14170
rect 8152 14118 8204 14170
rect 14842 14118 14894 14170
rect 14906 14118 14958 14170
rect 14970 14118 15022 14170
rect 15034 14118 15086 14170
rect 15098 14118 15150 14170
rect 21788 14118 21840 14170
rect 21852 14118 21904 14170
rect 21916 14118 21968 14170
rect 21980 14118 22032 14170
rect 22044 14118 22096 14170
rect 28734 14118 28786 14170
rect 28798 14118 28850 14170
rect 28862 14118 28914 14170
rect 28926 14118 28978 14170
rect 28990 14118 29042 14170
rect 1584 14059 1636 14068
rect 1584 14025 1593 14059
rect 1593 14025 1627 14059
rect 1627 14025 1636 14059
rect 1584 14016 1636 14025
rect 1860 14059 1912 14068
rect 1860 14025 1869 14059
rect 1869 14025 1903 14059
rect 1903 14025 1912 14059
rect 1860 14016 1912 14025
rect 6920 14016 6972 14068
rect 7104 14016 7156 14068
rect 9680 14016 9732 14068
rect 10416 14016 10468 14068
rect 12532 14016 12584 14068
rect 13176 14016 13228 14068
rect 1400 13923 1452 13932
rect 1400 13889 1409 13923
rect 1409 13889 1443 13923
rect 1443 13889 1452 13923
rect 1400 13880 1452 13889
rect 1676 13923 1728 13932
rect 1676 13889 1685 13923
rect 1685 13889 1719 13923
rect 1719 13889 1728 13923
rect 1676 13880 1728 13889
rect 7472 13948 7524 14000
rect 10048 13948 10100 14000
rect 11060 13948 11112 14000
rect 12440 13948 12492 14000
rect 14188 13948 14240 14000
rect 14740 13991 14792 14000
rect 14740 13957 14749 13991
rect 14749 13957 14783 13991
rect 14783 13957 14792 13991
rect 14740 13948 14792 13957
rect 17684 13948 17736 14000
rect 8392 13880 8444 13932
rect 9496 13880 9548 13932
rect 9588 13880 9640 13932
rect 7104 13812 7156 13864
rect 7380 13812 7432 13864
rect 9128 13855 9180 13864
rect 9128 13821 9137 13855
rect 9137 13821 9171 13855
rect 9171 13821 9180 13855
rect 9128 13812 9180 13821
rect 9312 13855 9364 13864
rect 9312 13821 9321 13855
rect 9321 13821 9355 13855
rect 9355 13821 9364 13855
rect 9312 13812 9364 13821
rect 2044 13744 2096 13796
rect 6736 13744 6788 13796
rect 8760 13744 8812 13796
rect 10140 13880 10192 13932
rect 10968 13923 11020 13932
rect 10968 13889 10977 13923
rect 10977 13889 11011 13923
rect 11011 13889 11020 13923
rect 10968 13880 11020 13889
rect 10416 13855 10468 13864
rect 10416 13821 10425 13855
rect 10425 13821 10459 13855
rect 10459 13821 10468 13855
rect 10416 13812 10468 13821
rect 11888 13812 11940 13864
rect 12348 13812 12400 13864
rect 15476 13880 15528 13932
rect 14280 13812 14332 13864
rect 15292 13812 15344 13864
rect 16488 13812 16540 13864
rect 28356 13855 28408 13864
rect 28356 13821 28365 13855
rect 28365 13821 28399 13855
rect 28399 13821 28408 13855
rect 28356 13812 28408 13821
rect 8116 13719 8168 13728
rect 8116 13685 8125 13719
rect 8125 13685 8159 13719
rect 8159 13685 8168 13719
rect 8116 13676 8168 13685
rect 8668 13719 8720 13728
rect 8668 13685 8677 13719
rect 8677 13685 8711 13719
rect 8711 13685 8720 13719
rect 8668 13676 8720 13685
rect 9680 13676 9732 13728
rect 11152 13676 11204 13728
rect 12164 13676 12216 13728
rect 12440 13676 12492 13728
rect 4423 13574 4475 13626
rect 4487 13574 4539 13626
rect 4551 13574 4603 13626
rect 4615 13574 4667 13626
rect 4679 13574 4731 13626
rect 11369 13574 11421 13626
rect 11433 13574 11485 13626
rect 11497 13574 11549 13626
rect 11561 13574 11613 13626
rect 11625 13574 11677 13626
rect 18315 13574 18367 13626
rect 18379 13574 18431 13626
rect 18443 13574 18495 13626
rect 18507 13574 18559 13626
rect 18571 13574 18623 13626
rect 25261 13574 25313 13626
rect 25325 13574 25377 13626
rect 25389 13574 25441 13626
rect 25453 13574 25505 13626
rect 25517 13574 25569 13626
rect 6736 13472 6788 13524
rect 8760 13472 8812 13524
rect 9128 13472 9180 13524
rect 1860 13447 1912 13456
rect 1860 13413 1869 13447
rect 1869 13413 1903 13447
rect 1903 13413 1912 13447
rect 1860 13404 1912 13413
rect 7656 13404 7708 13456
rect 8116 13404 8168 13456
rect 3976 13336 4028 13388
rect 6736 13336 6788 13388
rect 8300 13336 8352 13388
rect 8668 13379 8720 13388
rect 8668 13345 8677 13379
rect 8677 13345 8711 13379
rect 8711 13345 8720 13379
rect 8668 13336 8720 13345
rect 9036 13336 9088 13388
rect 9772 13336 9824 13388
rect 11060 13336 11112 13388
rect 11428 13379 11480 13388
rect 11428 13345 11437 13379
rect 11437 13345 11471 13379
rect 11471 13345 11480 13379
rect 11428 13336 11480 13345
rect 13728 13336 13780 13388
rect 940 13268 992 13320
rect 1032 13200 1084 13252
rect 5632 13268 5684 13320
rect 5724 13311 5776 13320
rect 5724 13277 5733 13311
rect 5733 13277 5767 13311
rect 5767 13277 5776 13311
rect 5724 13268 5776 13277
rect 8392 13268 8444 13320
rect 9128 13311 9180 13320
rect 9128 13277 9137 13311
rect 9137 13277 9171 13311
rect 9171 13277 9180 13311
rect 9128 13268 9180 13277
rect 11888 13311 11940 13320
rect 11888 13277 11897 13311
rect 11897 13277 11931 13311
rect 11931 13277 11940 13311
rect 11888 13268 11940 13277
rect 16028 13379 16080 13388
rect 16028 13345 16037 13379
rect 16037 13345 16071 13379
rect 16071 13345 16080 13379
rect 16028 13336 16080 13345
rect 6000 13243 6052 13252
rect 6000 13209 6009 13243
rect 6009 13209 6043 13243
rect 6043 13209 6052 13243
rect 6000 13200 6052 13209
rect 7380 13200 7432 13252
rect 10692 13200 10744 13252
rect 12164 13243 12216 13252
rect 12164 13209 12173 13243
rect 12173 13209 12207 13243
rect 12207 13209 12216 13243
rect 12164 13200 12216 13209
rect 13452 13200 13504 13252
rect 15752 13268 15804 13320
rect 1584 13175 1636 13184
rect 1584 13141 1593 13175
rect 1593 13141 1627 13175
rect 1627 13141 1636 13175
rect 1584 13132 1636 13141
rect 6828 13132 6880 13184
rect 8668 13132 8720 13184
rect 12900 13132 12952 13184
rect 25688 13200 25740 13252
rect 28356 13243 28408 13252
rect 28356 13209 28365 13243
rect 28365 13209 28399 13243
rect 28399 13209 28408 13243
rect 28356 13200 28408 13209
rect 15844 13175 15896 13184
rect 15844 13141 15853 13175
rect 15853 13141 15887 13175
rect 15887 13141 15896 13175
rect 15844 13132 15896 13141
rect 16396 13175 16448 13184
rect 16396 13141 16405 13175
rect 16405 13141 16439 13175
rect 16439 13141 16448 13175
rect 16396 13132 16448 13141
rect 7896 13030 7948 13082
rect 7960 13030 8012 13082
rect 8024 13030 8076 13082
rect 8088 13030 8140 13082
rect 8152 13030 8204 13082
rect 14842 13030 14894 13082
rect 14906 13030 14958 13082
rect 14970 13030 15022 13082
rect 15034 13030 15086 13082
rect 15098 13030 15150 13082
rect 21788 13030 21840 13082
rect 21852 13030 21904 13082
rect 21916 13030 21968 13082
rect 21980 13030 22032 13082
rect 22044 13030 22096 13082
rect 28734 13030 28786 13082
rect 28798 13030 28850 13082
rect 28862 13030 28914 13082
rect 28926 13030 28978 13082
rect 28990 13030 29042 13082
rect 940 12792 992 12844
rect 1676 12835 1728 12844
rect 1676 12801 1685 12835
rect 1685 12801 1719 12835
rect 1719 12801 1728 12835
rect 1676 12792 1728 12801
rect 1860 12699 1912 12708
rect 1860 12665 1869 12699
rect 1869 12665 1903 12699
rect 1903 12665 1912 12699
rect 1860 12656 1912 12665
rect 6000 12928 6052 12980
rect 6736 12971 6788 12980
rect 6736 12937 6745 12971
rect 6745 12937 6779 12971
rect 6779 12937 6788 12971
rect 6736 12928 6788 12937
rect 6828 12971 6880 12980
rect 6828 12937 6837 12971
rect 6837 12937 6871 12971
rect 6871 12937 6880 12971
rect 6828 12928 6880 12937
rect 7380 12928 7432 12980
rect 7472 12928 7524 12980
rect 7656 12928 7708 12980
rect 7840 12928 7892 12980
rect 5632 12860 5684 12912
rect 5908 12860 5960 12912
rect 7104 12724 7156 12776
rect 7380 12724 7432 12776
rect 6000 12588 6052 12640
rect 8024 12792 8076 12844
rect 8760 12928 8812 12980
rect 8668 12860 8720 12912
rect 10416 12971 10468 12980
rect 10416 12937 10425 12971
rect 10425 12937 10459 12971
rect 10459 12937 10468 12971
rect 10416 12928 10468 12937
rect 10692 12928 10744 12980
rect 12164 12928 12216 12980
rect 13452 12928 13504 12980
rect 9680 12792 9732 12844
rect 10600 12835 10652 12844
rect 10600 12801 10609 12835
rect 10609 12801 10643 12835
rect 10643 12801 10652 12835
rect 10600 12792 10652 12801
rect 10324 12767 10376 12776
rect 10324 12733 10333 12767
rect 10333 12733 10367 12767
rect 10367 12733 10376 12767
rect 11060 12835 11112 12844
rect 11060 12801 11069 12835
rect 11069 12801 11103 12835
rect 11103 12801 11112 12835
rect 11060 12792 11112 12801
rect 10324 12724 10376 12733
rect 12440 12767 12492 12776
rect 12440 12733 12449 12767
rect 12449 12733 12483 12767
rect 12483 12733 12492 12767
rect 12440 12724 12492 12733
rect 12532 12767 12584 12776
rect 12532 12733 12541 12767
rect 12541 12733 12575 12767
rect 12575 12733 12584 12767
rect 12532 12724 12584 12733
rect 12900 12724 12952 12776
rect 7932 12699 7984 12708
rect 7932 12665 7941 12699
rect 7941 12665 7975 12699
rect 7975 12665 7984 12699
rect 7932 12656 7984 12665
rect 9772 12656 9824 12708
rect 13820 12792 13872 12844
rect 14740 12928 14792 12980
rect 16396 12928 16448 12980
rect 22836 12928 22888 12980
rect 14648 12860 14700 12912
rect 17776 12860 17828 12912
rect 15292 12835 15344 12844
rect 15292 12801 15301 12835
rect 15301 12801 15335 12835
rect 15335 12801 15344 12835
rect 15292 12792 15344 12801
rect 16120 12835 16172 12844
rect 16120 12801 16129 12835
rect 16129 12801 16163 12835
rect 16163 12801 16172 12835
rect 16120 12792 16172 12801
rect 25780 12724 25832 12776
rect 11428 12588 11480 12640
rect 15476 12631 15528 12640
rect 15476 12597 15485 12631
rect 15485 12597 15519 12631
rect 15519 12597 15528 12631
rect 15476 12588 15528 12597
rect 17224 12588 17276 12640
rect 4423 12486 4475 12538
rect 4487 12486 4539 12538
rect 4551 12486 4603 12538
rect 4615 12486 4667 12538
rect 4679 12486 4731 12538
rect 11369 12486 11421 12538
rect 11433 12486 11485 12538
rect 11497 12486 11549 12538
rect 11561 12486 11613 12538
rect 11625 12486 11677 12538
rect 18315 12486 18367 12538
rect 18379 12486 18431 12538
rect 18443 12486 18495 12538
rect 18507 12486 18559 12538
rect 18571 12486 18623 12538
rect 25261 12486 25313 12538
rect 25325 12486 25377 12538
rect 25389 12486 25441 12538
rect 25453 12486 25505 12538
rect 25517 12486 25569 12538
rect 5724 12359 5776 12368
rect 5724 12325 5733 12359
rect 5733 12325 5767 12359
rect 5767 12325 5776 12359
rect 5724 12316 5776 12325
rect 7840 12316 7892 12368
rect 9036 12316 9088 12368
rect 7012 12248 7064 12300
rect 7380 12291 7432 12300
rect 7380 12257 7389 12291
rect 7389 12257 7423 12291
rect 7423 12257 7432 12291
rect 7380 12248 7432 12257
rect 940 12180 992 12232
rect 1032 12112 1084 12164
rect 6644 12180 6696 12232
rect 7748 12112 7800 12164
rect 1860 12087 1912 12096
rect 1860 12053 1869 12087
rect 1869 12053 1903 12087
rect 1903 12053 1912 12087
rect 1860 12044 1912 12053
rect 5172 12087 5224 12096
rect 5172 12053 5181 12087
rect 5181 12053 5215 12087
rect 5215 12053 5224 12087
rect 5172 12044 5224 12053
rect 6828 12044 6880 12096
rect 7932 12044 7984 12096
rect 8760 12248 8812 12300
rect 9864 12223 9916 12232
rect 9864 12189 9873 12223
rect 9873 12189 9907 12223
rect 9907 12189 9916 12223
rect 9864 12180 9916 12189
rect 15200 12427 15252 12436
rect 15200 12393 15209 12427
rect 15209 12393 15243 12427
rect 15243 12393 15252 12427
rect 15200 12384 15252 12393
rect 16212 12384 16264 12436
rect 10600 12316 10652 12368
rect 11796 12316 11848 12368
rect 11520 12248 11572 12300
rect 12348 12248 12400 12300
rect 12440 12291 12492 12300
rect 12440 12257 12449 12291
rect 12449 12257 12483 12291
rect 12483 12257 12492 12291
rect 12440 12248 12492 12257
rect 11060 12180 11112 12232
rect 11428 12180 11480 12232
rect 9312 12112 9364 12164
rect 16672 12384 16724 12436
rect 23480 12384 23532 12436
rect 15568 12223 15620 12232
rect 15568 12189 15577 12223
rect 15577 12189 15611 12223
rect 15611 12189 15620 12223
rect 15568 12180 15620 12189
rect 8668 12044 8720 12096
rect 8852 12044 8904 12096
rect 9588 12044 9640 12096
rect 10416 12087 10468 12096
rect 10416 12053 10425 12087
rect 10425 12053 10459 12087
rect 10459 12053 10468 12087
rect 10416 12044 10468 12053
rect 11244 12044 11296 12096
rect 12440 12044 12492 12096
rect 13728 12112 13780 12164
rect 20076 12112 20128 12164
rect 20168 12112 20220 12164
rect 28356 12155 28408 12164
rect 28356 12121 28365 12155
rect 28365 12121 28399 12155
rect 28399 12121 28408 12155
rect 28356 12112 28408 12121
rect 12992 12044 13044 12096
rect 13084 12087 13136 12096
rect 13084 12053 13093 12087
rect 13093 12053 13127 12087
rect 13127 12053 13136 12087
rect 13084 12044 13136 12053
rect 13636 12044 13688 12096
rect 14188 12087 14240 12096
rect 14188 12053 14197 12087
rect 14197 12053 14231 12087
rect 14231 12053 14240 12087
rect 14188 12044 14240 12053
rect 18880 12044 18932 12096
rect 7896 11942 7948 11994
rect 7960 11942 8012 11994
rect 8024 11942 8076 11994
rect 8088 11942 8140 11994
rect 8152 11942 8204 11994
rect 14842 11942 14894 11994
rect 14906 11942 14958 11994
rect 14970 11942 15022 11994
rect 15034 11942 15086 11994
rect 15098 11942 15150 11994
rect 21788 11942 21840 11994
rect 21852 11942 21904 11994
rect 21916 11942 21968 11994
rect 21980 11942 22032 11994
rect 22044 11942 22096 11994
rect 28734 11942 28786 11994
rect 28798 11942 28850 11994
rect 28862 11942 28914 11994
rect 28926 11942 28978 11994
rect 28990 11942 29042 11994
rect 6000 11883 6052 11892
rect 6000 11849 6009 11883
rect 6009 11849 6043 11883
rect 6043 11849 6052 11883
rect 6000 11840 6052 11849
rect 6828 11883 6880 11892
rect 6828 11849 6837 11883
rect 6837 11849 6871 11883
rect 6871 11849 6880 11883
rect 6828 11840 6880 11849
rect 8024 11840 8076 11892
rect 3608 11772 3660 11824
rect 940 11704 992 11756
rect 1032 11636 1084 11688
rect 3792 11704 3844 11756
rect 6368 11704 6420 11756
rect 6920 11772 6972 11824
rect 7380 11772 7432 11824
rect 8852 11840 8904 11892
rect 8760 11772 8812 11824
rect 10048 11840 10100 11892
rect 10416 11840 10468 11892
rect 11520 11840 11572 11892
rect 9588 11772 9640 11824
rect 9496 11704 9548 11756
rect 9864 11704 9916 11756
rect 7932 11636 7984 11688
rect 8208 11636 8260 11688
rect 8668 11679 8720 11688
rect 8668 11645 8677 11679
rect 8677 11645 8711 11679
rect 8711 11645 8720 11679
rect 8668 11636 8720 11645
rect 1860 11543 1912 11552
rect 1860 11509 1869 11543
rect 1869 11509 1903 11543
rect 1903 11509 1912 11543
rect 1860 11500 1912 11509
rect 8668 11500 8720 11552
rect 9588 11568 9640 11620
rect 13084 11840 13136 11892
rect 16672 11840 16724 11892
rect 14188 11772 14240 11824
rect 11060 11704 11112 11756
rect 11428 11636 11480 11688
rect 11980 11747 12032 11756
rect 11980 11713 11989 11747
rect 11989 11713 12023 11747
rect 12023 11713 12032 11747
rect 11980 11704 12032 11713
rect 13728 11704 13780 11756
rect 17776 11840 17828 11892
rect 20168 11840 20220 11892
rect 17132 11747 17184 11756
rect 17132 11713 17141 11747
rect 17141 11713 17175 11747
rect 17175 11713 17184 11747
rect 17132 11704 17184 11713
rect 12348 11636 12400 11688
rect 13544 11636 13596 11688
rect 11888 11568 11940 11620
rect 28356 11679 28408 11688
rect 28356 11645 28365 11679
rect 28365 11645 28399 11679
rect 28399 11645 28408 11679
rect 28356 11636 28408 11645
rect 9036 11500 9088 11552
rect 9496 11500 9548 11552
rect 11704 11500 11756 11552
rect 12256 11500 12308 11552
rect 19248 11500 19300 11552
rect 26700 11543 26752 11552
rect 26700 11509 26709 11543
rect 26709 11509 26743 11543
rect 26743 11509 26752 11543
rect 26700 11500 26752 11509
rect 4423 11398 4475 11450
rect 4487 11398 4539 11450
rect 4551 11398 4603 11450
rect 4615 11398 4667 11450
rect 4679 11398 4731 11450
rect 11369 11398 11421 11450
rect 11433 11398 11485 11450
rect 11497 11398 11549 11450
rect 11561 11398 11613 11450
rect 11625 11398 11677 11450
rect 18315 11398 18367 11450
rect 18379 11398 18431 11450
rect 18443 11398 18495 11450
rect 18507 11398 18559 11450
rect 18571 11398 18623 11450
rect 25261 11398 25313 11450
rect 25325 11398 25377 11450
rect 25389 11398 25441 11450
rect 25453 11398 25505 11450
rect 25517 11398 25569 11450
rect 1860 11296 1912 11348
rect 5724 11228 5776 11280
rect 7380 11228 7432 11280
rect 3332 11160 3384 11212
rect 1400 11135 1452 11144
rect 1400 11101 1409 11135
rect 1409 11101 1443 11135
rect 1443 11101 1452 11135
rect 1400 11092 1452 11101
rect 1676 11135 1728 11144
rect 1676 11101 1685 11135
rect 1685 11101 1719 11135
rect 1719 11101 1728 11135
rect 1676 11092 1728 11101
rect 4896 11024 4948 11076
rect 5908 11135 5960 11144
rect 5908 11101 5917 11135
rect 5917 11101 5951 11135
rect 5951 11101 5960 11135
rect 5908 11092 5960 11101
rect 6000 11092 6052 11144
rect 7472 11092 7524 11144
rect 7656 11160 7708 11212
rect 8852 11160 8904 11212
rect 8944 11203 8996 11212
rect 8944 11169 8953 11203
rect 8953 11169 8987 11203
rect 8987 11169 8996 11203
rect 8944 11160 8996 11169
rect 9312 11203 9364 11212
rect 9312 11169 9321 11203
rect 9321 11169 9355 11203
rect 9355 11169 9364 11203
rect 9312 11160 9364 11169
rect 10048 11160 10100 11212
rect 5356 10999 5408 11008
rect 5356 10965 5365 10999
rect 5365 10965 5399 10999
rect 5399 10965 5408 10999
rect 5356 10956 5408 10965
rect 6644 11024 6696 11076
rect 8024 11024 8076 11076
rect 8392 11135 8444 11144
rect 8392 11101 8401 11135
rect 8401 11101 8435 11135
rect 8435 11101 8444 11135
rect 8392 11092 8444 11101
rect 9588 11092 9640 11144
rect 12440 11296 12492 11348
rect 11244 11092 11296 11144
rect 11520 11135 11572 11144
rect 11520 11101 11529 11135
rect 11529 11101 11563 11135
rect 11563 11101 11572 11135
rect 11520 11092 11572 11101
rect 13084 11092 13136 11144
rect 7380 10956 7432 11008
rect 9772 10956 9824 11008
rect 10232 10956 10284 11008
rect 11888 11024 11940 11076
rect 12256 11024 12308 11076
rect 16580 11160 16632 11212
rect 14464 11067 14516 11076
rect 14464 11033 14473 11067
rect 14473 11033 14507 11067
rect 14507 11033 14516 11067
rect 14464 11024 14516 11033
rect 13544 10956 13596 11008
rect 7896 10854 7948 10906
rect 7960 10854 8012 10906
rect 8024 10854 8076 10906
rect 8088 10854 8140 10906
rect 8152 10854 8204 10906
rect 14842 10854 14894 10906
rect 14906 10854 14958 10906
rect 14970 10854 15022 10906
rect 15034 10854 15086 10906
rect 15098 10854 15150 10906
rect 21788 10854 21840 10906
rect 21852 10854 21904 10906
rect 21916 10854 21968 10906
rect 21980 10854 22032 10906
rect 22044 10854 22096 10906
rect 28734 10854 28786 10906
rect 28798 10854 28850 10906
rect 28862 10854 28914 10906
rect 28926 10854 28978 10906
rect 28990 10854 29042 10906
rect 5908 10752 5960 10804
rect 6184 10752 6236 10804
rect 7012 10752 7064 10804
rect 7472 10752 7524 10804
rect 10508 10795 10560 10804
rect 10508 10761 10517 10795
rect 10517 10761 10551 10795
rect 10551 10761 10560 10795
rect 10508 10752 10560 10761
rect 5080 10684 5132 10736
rect 940 10616 992 10668
rect 1032 10548 1084 10600
rect 4160 10616 4212 10668
rect 5724 10684 5776 10736
rect 4344 10548 4396 10600
rect 6184 10548 6236 10600
rect 6552 10659 6604 10668
rect 6552 10625 6561 10659
rect 6561 10625 6595 10659
rect 6595 10625 6604 10659
rect 6552 10616 6604 10625
rect 6644 10616 6696 10668
rect 6828 10616 6880 10668
rect 7748 10616 7800 10668
rect 9680 10684 9732 10736
rect 10416 10684 10468 10736
rect 12808 10684 12860 10736
rect 13544 10727 13596 10736
rect 13544 10693 13553 10727
rect 13553 10693 13587 10727
rect 13587 10693 13596 10727
rect 13544 10684 13596 10693
rect 13728 10659 13780 10668
rect 13728 10625 13737 10659
rect 13737 10625 13771 10659
rect 13771 10625 13780 10659
rect 13728 10616 13780 10625
rect 8300 10548 8352 10600
rect 1584 10523 1636 10532
rect 1584 10489 1593 10523
rect 1593 10489 1627 10523
rect 1627 10489 1636 10523
rect 1584 10480 1636 10489
rect 6460 10480 6512 10532
rect 6552 10480 6604 10532
rect 10324 10591 10376 10600
rect 10324 10557 10333 10591
rect 10333 10557 10367 10591
rect 10367 10557 10376 10591
rect 10324 10548 10376 10557
rect 10876 10548 10928 10600
rect 11520 10591 11572 10600
rect 11520 10557 11529 10591
rect 11529 10557 11563 10591
rect 11563 10557 11572 10591
rect 11520 10548 11572 10557
rect 11796 10591 11848 10600
rect 11796 10557 11805 10591
rect 11805 10557 11839 10591
rect 11839 10557 11848 10591
rect 11796 10548 11848 10557
rect 9956 10480 10008 10532
rect 4160 10412 4212 10464
rect 10048 10412 10100 10464
rect 10140 10412 10192 10464
rect 26700 10752 26752 10804
rect 16028 10684 16080 10736
rect 15936 10659 15988 10668
rect 15936 10625 15945 10659
rect 15945 10625 15979 10659
rect 15979 10625 15988 10659
rect 15936 10616 15988 10625
rect 17132 10616 17184 10668
rect 28356 10591 28408 10600
rect 28356 10557 28365 10591
rect 28365 10557 28399 10591
rect 28399 10557 28408 10591
rect 28356 10548 28408 10557
rect 14004 10455 14056 10464
rect 14004 10421 14013 10455
rect 14013 10421 14047 10455
rect 14047 10421 14056 10455
rect 14004 10412 14056 10421
rect 16120 10455 16172 10464
rect 16120 10421 16129 10455
rect 16129 10421 16163 10455
rect 16163 10421 16172 10455
rect 16120 10412 16172 10421
rect 4423 10310 4475 10362
rect 4487 10310 4539 10362
rect 4551 10310 4603 10362
rect 4615 10310 4667 10362
rect 4679 10310 4731 10362
rect 11369 10310 11421 10362
rect 11433 10310 11485 10362
rect 11497 10310 11549 10362
rect 11561 10310 11613 10362
rect 11625 10310 11677 10362
rect 18315 10310 18367 10362
rect 18379 10310 18431 10362
rect 18443 10310 18495 10362
rect 18507 10310 18559 10362
rect 18571 10310 18623 10362
rect 25261 10310 25313 10362
rect 25325 10310 25377 10362
rect 25389 10310 25441 10362
rect 25453 10310 25505 10362
rect 25517 10310 25569 10362
rect 296 10208 348 10260
rect 664 10208 716 10260
rect 6460 10208 6512 10260
rect 7380 10208 7432 10260
rect 8484 10208 8536 10260
rect 9864 10251 9916 10260
rect 9864 10217 9873 10251
rect 9873 10217 9907 10251
rect 9907 10217 9916 10251
rect 9864 10208 9916 10217
rect 10048 10208 10100 10260
rect 11796 10208 11848 10260
rect 12808 10208 12860 10260
rect 17132 10208 17184 10260
rect 17224 10208 17276 10260
rect 9680 10140 9732 10192
rect 6000 10072 6052 10124
rect 7012 10072 7064 10124
rect 9956 10115 10008 10124
rect 9956 10081 9965 10115
rect 9965 10081 9999 10115
rect 9999 10081 10008 10115
rect 9956 10072 10008 10081
rect 12072 10140 12124 10192
rect 12440 10115 12492 10124
rect 12440 10081 12449 10115
rect 12449 10081 12483 10115
rect 12483 10081 12492 10115
rect 12440 10072 12492 10081
rect 940 10004 992 10056
rect 1676 10047 1728 10056
rect 1676 10013 1685 10047
rect 1685 10013 1719 10047
rect 1719 10013 1728 10047
rect 1676 10004 1728 10013
rect 6644 10004 6696 10056
rect 3148 9868 3200 9920
rect 4804 9911 4856 9920
rect 4804 9877 4813 9911
rect 4813 9877 4847 9911
rect 4847 9877 4856 9911
rect 4804 9868 4856 9877
rect 5356 9936 5408 9988
rect 5724 9936 5776 9988
rect 8668 10004 8720 10056
rect 9220 10004 9272 10056
rect 9864 10004 9916 10056
rect 12348 10004 12400 10056
rect 10140 9936 10192 9988
rect 11520 9936 11572 9988
rect 28356 9979 28408 9988
rect 28356 9945 28365 9979
rect 28365 9945 28399 9979
rect 28399 9945 28408 9979
rect 28356 9936 28408 9945
rect 11060 9868 11112 9920
rect 7896 9766 7948 9818
rect 7960 9766 8012 9818
rect 8024 9766 8076 9818
rect 8088 9766 8140 9818
rect 8152 9766 8204 9818
rect 14842 9766 14894 9818
rect 14906 9766 14958 9818
rect 14970 9766 15022 9818
rect 15034 9766 15086 9818
rect 15098 9766 15150 9818
rect 21788 9766 21840 9818
rect 21852 9766 21904 9818
rect 21916 9766 21968 9818
rect 21980 9766 22032 9818
rect 22044 9766 22096 9818
rect 28734 9766 28786 9818
rect 28798 9766 28850 9818
rect 28862 9766 28914 9818
rect 28926 9766 28978 9818
rect 28990 9766 29042 9818
rect 5908 9664 5960 9716
rect 6828 9664 6880 9716
rect 4620 9639 4672 9648
rect 4620 9605 4629 9639
rect 4629 9605 4663 9639
rect 4663 9605 4672 9639
rect 4620 9596 4672 9605
rect 4712 9596 4764 9648
rect 7840 9664 7892 9716
rect 17224 9664 17276 9716
rect 940 9528 992 9580
rect 1032 9460 1084 9512
rect 1768 9528 1820 9580
rect 2044 9528 2096 9580
rect 7196 9596 7248 9648
rect 7380 9596 7432 9648
rect 5080 9571 5132 9580
rect 5080 9537 5089 9571
rect 5089 9537 5123 9571
rect 5123 9537 5132 9571
rect 5080 9528 5132 9537
rect 5172 9569 5224 9580
rect 5172 9535 5181 9569
rect 5181 9535 5215 9569
rect 5215 9535 5224 9569
rect 5172 9528 5224 9535
rect 6184 9571 6236 9580
rect 6184 9537 6193 9571
rect 6193 9537 6227 9571
rect 6227 9537 6236 9571
rect 6184 9528 6236 9537
rect 6460 9528 6512 9580
rect 6552 9528 6604 9580
rect 8484 9528 8536 9580
rect 9404 9596 9456 9648
rect 10140 9596 10192 9648
rect 12072 9596 12124 9648
rect 5908 9460 5960 9512
rect 9680 9460 9732 9512
rect 10508 9460 10560 9512
rect 11704 9528 11756 9580
rect 14188 9571 14240 9580
rect 14188 9537 14197 9571
rect 14197 9537 14231 9571
rect 14231 9537 14240 9571
rect 14188 9528 14240 9537
rect 2136 9367 2188 9376
rect 2136 9333 2145 9367
rect 2145 9333 2179 9367
rect 2179 9333 2188 9367
rect 2136 9324 2188 9333
rect 2412 9367 2464 9376
rect 2412 9333 2421 9367
rect 2421 9333 2455 9367
rect 2455 9333 2464 9367
rect 2412 9324 2464 9333
rect 3792 9324 3844 9376
rect 4160 9367 4212 9376
rect 4160 9333 4169 9367
rect 4169 9333 4203 9367
rect 4203 9333 4212 9367
rect 4160 9324 4212 9333
rect 5632 9392 5684 9444
rect 10048 9392 10100 9444
rect 11428 9392 11480 9444
rect 13544 9392 13596 9444
rect 17224 9392 17276 9444
rect 23848 9392 23900 9444
rect 5172 9324 5224 9376
rect 5356 9367 5408 9376
rect 5356 9333 5365 9367
rect 5365 9333 5399 9367
rect 5399 9333 5408 9367
rect 5356 9324 5408 9333
rect 5816 9324 5868 9376
rect 7104 9324 7156 9376
rect 7748 9324 7800 9376
rect 9496 9324 9548 9376
rect 10324 9367 10376 9376
rect 10324 9333 10333 9367
rect 10333 9333 10367 9367
rect 10367 9333 10376 9367
rect 10324 9324 10376 9333
rect 11244 9324 11296 9376
rect 11796 9367 11848 9376
rect 11796 9333 11805 9367
rect 11805 9333 11839 9367
rect 11839 9333 11848 9367
rect 11796 9324 11848 9333
rect 13820 9324 13872 9376
rect 25780 9324 25832 9376
rect 4423 9222 4475 9274
rect 4487 9222 4539 9274
rect 4551 9222 4603 9274
rect 4615 9222 4667 9274
rect 4679 9222 4731 9274
rect 11369 9222 11421 9274
rect 11433 9222 11485 9274
rect 11497 9222 11549 9274
rect 11561 9222 11613 9274
rect 11625 9222 11677 9274
rect 18315 9222 18367 9274
rect 18379 9222 18431 9274
rect 18443 9222 18495 9274
rect 18507 9222 18559 9274
rect 18571 9222 18623 9274
rect 25261 9222 25313 9274
rect 25325 9222 25377 9274
rect 25389 9222 25441 9274
rect 25453 9222 25505 9274
rect 25517 9222 25569 9274
rect 1584 9095 1636 9104
rect 1584 9061 1593 9095
rect 1593 9061 1627 9095
rect 1627 9061 1636 9095
rect 1584 9052 1636 9061
rect 5448 9052 5500 9104
rect 5632 9163 5684 9172
rect 5632 9129 5641 9163
rect 5641 9129 5675 9163
rect 5675 9129 5684 9163
rect 5632 9120 5684 9129
rect 5816 9120 5868 9172
rect 6460 9120 6512 9172
rect 7472 9120 7524 9172
rect 7564 9120 7616 9172
rect 1308 8984 1360 9036
rect 940 8916 992 8968
rect 1032 8848 1084 8900
rect 1860 8916 1912 8968
rect 2228 8959 2280 8968
rect 2228 8925 2237 8959
rect 2237 8925 2271 8959
rect 2271 8925 2280 8959
rect 2228 8916 2280 8925
rect 848 8780 900 8832
rect 2320 8848 2372 8900
rect 1952 8823 2004 8832
rect 1952 8789 1961 8823
rect 1961 8789 1995 8823
rect 1995 8789 2004 8823
rect 1952 8780 2004 8789
rect 2504 8916 2556 8968
rect 3516 8984 3568 9036
rect 3608 8916 3660 8968
rect 5172 8916 5224 8968
rect 2780 8848 2832 8900
rect 3424 8848 3476 8900
rect 5448 8959 5500 8968
rect 5448 8925 5457 8959
rect 5457 8925 5491 8959
rect 5491 8925 5500 8959
rect 5448 8916 5500 8925
rect 2504 8823 2556 8832
rect 2504 8789 2513 8823
rect 2513 8789 2547 8823
rect 2547 8789 2556 8823
rect 2504 8780 2556 8789
rect 3148 8780 3200 8832
rect 3516 8780 3568 8832
rect 4712 8780 4764 8832
rect 5540 8780 5592 8832
rect 9864 9120 9916 9172
rect 10600 9120 10652 9172
rect 23480 9120 23532 9172
rect 10232 9052 10284 9104
rect 7840 9027 7892 9036
rect 7840 8993 7849 9027
rect 7849 8993 7883 9027
rect 7883 8993 7892 9027
rect 7840 8984 7892 8993
rect 9312 8984 9364 9036
rect 9680 8984 9732 9036
rect 8944 8959 8996 8968
rect 8944 8925 8953 8959
rect 8953 8925 8987 8959
rect 8987 8925 8996 8959
rect 8944 8916 8996 8925
rect 10600 8916 10652 8968
rect 6000 8848 6052 8900
rect 9220 8891 9272 8900
rect 9220 8857 9229 8891
rect 9229 8857 9263 8891
rect 9263 8857 9272 8891
rect 9220 8848 9272 8857
rect 9772 8848 9824 8900
rect 10508 8780 10560 8832
rect 10600 8780 10652 8832
rect 11060 8959 11112 8968
rect 11060 8925 11069 8959
rect 11069 8925 11103 8959
rect 11103 8925 11112 8959
rect 11060 8916 11112 8925
rect 12072 9027 12124 9036
rect 12072 8993 12081 9027
rect 12081 8993 12115 9027
rect 12115 8993 12124 9027
rect 12072 8984 12124 8993
rect 26608 8984 26660 9036
rect 28816 8984 28868 9036
rect 27160 8959 27212 8968
rect 27160 8925 27169 8959
rect 27169 8925 27203 8959
rect 27203 8925 27212 8959
rect 27160 8916 27212 8925
rect 26884 8848 26936 8900
rect 12440 8823 12492 8832
rect 12440 8789 12449 8823
rect 12449 8789 12483 8823
rect 12483 8789 12492 8823
rect 12440 8780 12492 8789
rect 7896 8678 7948 8730
rect 7960 8678 8012 8730
rect 8024 8678 8076 8730
rect 8088 8678 8140 8730
rect 8152 8678 8204 8730
rect 14842 8678 14894 8730
rect 14906 8678 14958 8730
rect 14970 8678 15022 8730
rect 15034 8678 15086 8730
rect 15098 8678 15150 8730
rect 21788 8678 21840 8730
rect 21852 8678 21904 8730
rect 21916 8678 21968 8730
rect 21980 8678 22032 8730
rect 22044 8678 22096 8730
rect 28734 8678 28786 8730
rect 28798 8678 28850 8730
rect 28862 8678 28914 8730
rect 28926 8678 28978 8730
rect 28990 8678 29042 8730
rect 1584 8619 1636 8628
rect 1584 8585 1593 8619
rect 1593 8585 1627 8619
rect 1627 8585 1636 8619
rect 1584 8576 1636 8585
rect 1492 8508 1544 8560
rect 2044 8508 2096 8560
rect 2780 8619 2832 8628
rect 2780 8585 2789 8619
rect 2789 8585 2823 8619
rect 2823 8585 2832 8619
rect 2780 8576 2832 8585
rect 1400 8483 1452 8492
rect 1400 8449 1409 8483
rect 1409 8449 1443 8483
rect 1443 8449 1452 8483
rect 1400 8440 1452 8449
rect 1676 8483 1728 8492
rect 1676 8449 1685 8483
rect 1685 8449 1719 8483
rect 1719 8449 1728 8483
rect 1676 8440 1728 8449
rect 756 8372 808 8424
rect 1032 8372 1084 8424
rect 2136 8440 2188 8492
rect 2320 8440 2372 8492
rect 2872 8440 2924 8492
rect 2964 8483 3016 8492
rect 2964 8449 2973 8483
rect 2973 8449 3007 8483
rect 3007 8449 3016 8483
rect 2964 8440 3016 8449
rect 3148 8440 3200 8492
rect 3332 8483 3384 8492
rect 3332 8449 3341 8483
rect 3341 8449 3375 8483
rect 3375 8449 3384 8483
rect 3332 8440 3384 8449
rect 5908 8576 5960 8628
rect 6184 8576 6236 8628
rect 4988 8508 5040 8560
rect 5540 8508 5592 8560
rect 7288 8576 7340 8628
rect 7748 8576 7800 8628
rect 8576 8619 8628 8628
rect 8576 8585 8585 8619
rect 8585 8585 8619 8619
rect 8619 8585 8628 8619
rect 8576 8576 8628 8585
rect 9220 8576 9272 8628
rect 10600 8576 10652 8628
rect 10784 8576 10836 8628
rect 11152 8576 11204 8628
rect 27160 8576 27212 8628
rect 3700 8440 3752 8492
rect 5172 8440 5224 8492
rect 7380 8440 7432 8492
rect 17224 8508 17276 8560
rect 2320 8304 2372 8356
rect 3056 8347 3108 8356
rect 3056 8313 3065 8347
rect 3065 8313 3099 8347
rect 3099 8313 3108 8347
rect 3056 8304 3108 8313
rect 6092 8415 6144 8424
rect 6092 8381 6101 8415
rect 6101 8381 6135 8415
rect 6135 8381 6144 8415
rect 6092 8372 6144 8381
rect 6276 8372 6328 8424
rect 7748 8415 7800 8424
rect 7748 8381 7757 8415
rect 7757 8381 7791 8415
rect 7791 8381 7800 8415
rect 7748 8372 7800 8381
rect 8576 8372 8628 8424
rect 4712 8304 4764 8356
rect 1032 8236 1084 8288
rect 1584 8236 1636 8288
rect 1952 8236 2004 8288
rect 2044 8236 2096 8288
rect 4252 8236 4304 8288
rect 10508 8440 10560 8492
rect 11060 8372 11112 8424
rect 11244 8415 11296 8424
rect 11244 8381 11253 8415
rect 11253 8381 11287 8415
rect 11287 8381 11296 8415
rect 11244 8372 11296 8381
rect 12164 8415 12216 8424
rect 12164 8381 12173 8415
rect 12173 8381 12207 8415
rect 12207 8381 12216 8415
rect 12164 8372 12216 8381
rect 28356 8415 28408 8424
rect 28356 8381 28365 8415
rect 28365 8381 28399 8415
rect 28399 8381 28408 8415
rect 28356 8372 28408 8381
rect 7656 8236 7708 8288
rect 23388 8236 23440 8288
rect 4423 8134 4475 8186
rect 4487 8134 4539 8186
rect 4551 8134 4603 8186
rect 4615 8134 4667 8186
rect 4679 8134 4731 8186
rect 11369 8134 11421 8186
rect 11433 8134 11485 8186
rect 11497 8134 11549 8186
rect 11561 8134 11613 8186
rect 11625 8134 11677 8186
rect 18315 8134 18367 8186
rect 18379 8134 18431 8186
rect 18443 8134 18495 8186
rect 18507 8134 18559 8186
rect 18571 8134 18623 8186
rect 25261 8134 25313 8186
rect 25325 8134 25377 8186
rect 25389 8134 25441 8186
rect 25453 8134 25505 8186
rect 25517 8134 25569 8186
rect 1400 8032 1452 8084
rect 1676 8032 1728 8084
rect 480 7964 532 8016
rect 1400 7828 1452 7880
rect 1584 7828 1636 7880
rect 2044 7828 2096 7880
rect 3240 7939 3292 7948
rect 3240 7905 3249 7939
rect 3249 7905 3283 7939
rect 3283 7905 3292 7939
rect 3240 7896 3292 7905
rect 3884 7896 3936 7948
rect 4160 7896 4212 7948
rect 5080 8032 5132 8084
rect 5632 8032 5684 8084
rect 5908 8032 5960 8084
rect 7196 8032 7248 8084
rect 9128 8032 9180 8084
rect 10968 8032 11020 8084
rect 13176 8032 13228 8084
rect 27160 8032 27212 8084
rect 1952 7803 2004 7812
rect 1952 7769 1961 7803
rect 1961 7769 1995 7803
rect 1995 7769 2004 7803
rect 1952 7760 2004 7769
rect 756 7556 808 7608
rect 664 7488 716 7540
rect 1584 7735 1636 7744
rect 1584 7701 1593 7735
rect 1593 7701 1627 7735
rect 1627 7701 1636 7735
rect 1584 7692 1636 7701
rect 2136 7692 2188 7744
rect 2412 7735 2464 7744
rect 2412 7701 2421 7735
rect 2421 7701 2455 7735
rect 2455 7701 2464 7735
rect 2412 7692 2464 7701
rect 2688 7735 2740 7744
rect 2688 7701 2697 7735
rect 2697 7701 2731 7735
rect 2731 7701 2740 7735
rect 2688 7692 2740 7701
rect 3148 7692 3200 7744
rect 3424 7871 3476 7880
rect 3424 7837 3433 7871
rect 3433 7837 3467 7871
rect 3467 7837 3476 7871
rect 3424 7828 3476 7837
rect 3976 7871 4028 7880
rect 3976 7837 3985 7871
rect 3985 7837 4019 7871
rect 4019 7837 4028 7871
rect 3976 7828 4028 7837
rect 6460 7964 6512 8016
rect 4988 7896 5040 7948
rect 7656 7896 7708 7948
rect 8208 7896 8260 7948
rect 8300 7896 8352 7948
rect 12256 7964 12308 8016
rect 23388 7964 23440 8016
rect 5080 7828 5132 7880
rect 6736 7828 6788 7880
rect 5540 7760 5592 7812
rect 7012 7760 7064 7812
rect 3516 7692 3568 7744
rect 3884 7692 3936 7744
rect 4160 7735 4212 7744
rect 4160 7701 4169 7735
rect 4169 7701 4203 7735
rect 4203 7701 4212 7735
rect 4160 7692 4212 7701
rect 4804 7692 4856 7744
rect 4988 7735 5040 7744
rect 4988 7701 4997 7735
rect 4997 7701 5031 7735
rect 5031 7701 5040 7735
rect 4988 7692 5040 7701
rect 5724 7692 5776 7744
rect 7288 7760 7340 7812
rect 9680 7828 9732 7880
rect 8576 7760 8628 7812
rect 9128 7760 9180 7812
rect 10416 7871 10468 7880
rect 10416 7837 10425 7871
rect 10425 7837 10459 7871
rect 10459 7837 10468 7871
rect 10416 7828 10468 7837
rect 10508 7828 10560 7880
rect 10692 7828 10744 7880
rect 12532 7828 12584 7880
rect 27620 7939 27672 7948
rect 27620 7905 27629 7939
rect 27629 7905 27663 7939
rect 27663 7905 27672 7939
rect 27620 7896 27672 7905
rect 15476 7828 15528 7880
rect 14648 7760 14700 7812
rect 10048 7735 10100 7744
rect 10048 7701 10057 7735
rect 10057 7701 10091 7735
rect 10091 7701 10100 7735
rect 10048 7692 10100 7701
rect 7896 7590 7948 7642
rect 7960 7590 8012 7642
rect 8024 7590 8076 7642
rect 8088 7590 8140 7642
rect 8152 7590 8204 7642
rect 14842 7590 14894 7642
rect 14906 7590 14958 7642
rect 14970 7590 15022 7642
rect 15034 7590 15086 7642
rect 15098 7590 15150 7642
rect 21788 7590 21840 7642
rect 21852 7590 21904 7642
rect 21916 7590 21968 7642
rect 21980 7590 22032 7642
rect 22044 7590 22096 7642
rect 28734 7590 28786 7642
rect 28798 7590 28850 7642
rect 28862 7590 28914 7642
rect 28926 7590 28978 7642
rect 28990 7590 29042 7642
rect 1768 7531 1820 7540
rect 1768 7497 1777 7531
rect 1777 7497 1811 7531
rect 1811 7497 1820 7531
rect 1768 7488 1820 7497
rect 3976 7488 4028 7540
rect 4252 7488 4304 7540
rect 4988 7488 5040 7540
rect 6184 7488 6236 7540
rect 6920 7488 6972 7540
rect 7012 7488 7064 7540
rect 8392 7488 8444 7540
rect 1216 7420 1268 7472
rect 940 7352 992 7404
rect 2504 7352 2556 7404
rect 3608 7420 3660 7472
rect 5724 7420 5776 7472
rect 6828 7420 6880 7472
rect 1952 7327 2004 7336
rect 1952 7293 1961 7327
rect 1961 7293 1995 7327
rect 1995 7293 2004 7327
rect 1952 7284 2004 7293
rect 3608 7284 3660 7336
rect 4068 7284 4120 7336
rect 4712 7284 4764 7336
rect 6276 7352 6328 7404
rect 6460 7352 6512 7404
rect 8576 7420 8628 7472
rect 1584 7216 1636 7268
rect 2504 7259 2556 7268
rect 2504 7225 2513 7259
rect 2513 7225 2547 7259
rect 2547 7225 2556 7259
rect 2504 7216 2556 7225
rect 6092 7284 6144 7336
rect 5908 7216 5960 7268
rect 3700 7148 3752 7200
rect 4988 7148 5040 7200
rect 7012 7327 7064 7336
rect 7012 7293 7021 7327
rect 7021 7293 7055 7327
rect 7055 7293 7064 7327
rect 7012 7284 7064 7293
rect 6552 7216 6604 7268
rect 9772 7531 9824 7540
rect 9772 7497 9781 7531
rect 9781 7497 9815 7531
rect 9815 7497 9824 7531
rect 9772 7488 9824 7497
rect 10048 7488 10100 7540
rect 24400 7488 24452 7540
rect 9128 7395 9180 7404
rect 9128 7361 9137 7395
rect 9137 7361 9171 7395
rect 9171 7361 9180 7395
rect 9128 7352 9180 7361
rect 9220 7352 9272 7404
rect 9404 7352 9456 7404
rect 9864 7352 9916 7404
rect 10508 7463 10560 7472
rect 10508 7429 10517 7463
rect 10517 7429 10551 7463
rect 10551 7429 10560 7463
rect 10508 7420 10560 7429
rect 12256 7420 12308 7472
rect 29184 7420 29236 7472
rect 10324 7352 10376 7404
rect 11796 7352 11848 7404
rect 16304 7352 16356 7404
rect 27160 7395 27212 7404
rect 27160 7361 27169 7395
rect 27169 7361 27203 7395
rect 27203 7361 27212 7395
rect 27160 7352 27212 7361
rect 8760 7327 8812 7336
rect 8760 7293 8769 7327
rect 8769 7293 8803 7327
rect 8803 7293 8812 7327
rect 8760 7284 8812 7293
rect 9036 7284 9088 7336
rect 9772 7284 9824 7336
rect 28356 7327 28408 7336
rect 28356 7293 28365 7327
rect 28365 7293 28399 7327
rect 28399 7293 28408 7327
rect 28356 7284 28408 7293
rect 10508 7216 10560 7268
rect 8668 7148 8720 7200
rect 9312 7191 9364 7200
rect 9312 7157 9321 7191
rect 9321 7157 9355 7191
rect 9355 7157 9364 7191
rect 9312 7148 9364 7157
rect 10784 7148 10836 7200
rect 11152 7191 11204 7200
rect 11152 7157 11161 7191
rect 11161 7157 11195 7191
rect 11195 7157 11204 7191
rect 11152 7148 11204 7157
rect 4423 7046 4475 7098
rect 4487 7046 4539 7098
rect 4551 7046 4603 7098
rect 4615 7046 4667 7098
rect 4679 7046 4731 7098
rect 11369 7046 11421 7098
rect 11433 7046 11485 7098
rect 11497 7046 11549 7098
rect 11561 7046 11613 7098
rect 11625 7046 11677 7098
rect 18315 7046 18367 7098
rect 18379 7046 18431 7098
rect 18443 7046 18495 7098
rect 18507 7046 18559 7098
rect 18571 7046 18623 7098
rect 25261 7046 25313 7098
rect 25325 7046 25377 7098
rect 25389 7046 25441 7098
rect 25453 7046 25505 7098
rect 25517 7046 25569 7098
rect 7840 6944 7892 6996
rect 3240 6876 3292 6928
rect 3608 6876 3660 6928
rect 9312 6944 9364 6996
rect 1124 6808 1176 6860
rect 296 6740 348 6792
rect 4896 6808 4948 6860
rect 5080 6851 5132 6860
rect 5080 6817 5089 6851
rect 5089 6817 5123 6851
rect 5123 6817 5132 6851
rect 5080 6808 5132 6817
rect 2504 6783 2556 6792
rect 2504 6749 2513 6783
rect 2513 6749 2547 6783
rect 2547 6749 2556 6783
rect 2504 6740 2556 6749
rect 1308 6672 1360 6724
rect 2872 6740 2924 6792
rect 3792 6740 3844 6792
rect 3516 6672 3568 6724
rect 1860 6647 1912 6656
rect 1860 6613 1869 6647
rect 1869 6613 1903 6647
rect 1903 6613 1912 6647
rect 1860 6604 1912 6613
rect 3884 6604 3936 6656
rect 6460 6740 6512 6792
rect 6828 6808 6880 6860
rect 11980 6876 12032 6928
rect 24952 6876 25004 6928
rect 8668 6851 8720 6860
rect 8668 6817 8677 6851
rect 8677 6817 8711 6851
rect 8711 6817 8720 6851
rect 8668 6808 8720 6817
rect 9036 6808 9088 6860
rect 9588 6851 9640 6860
rect 9588 6817 9597 6851
rect 9597 6817 9631 6851
rect 9631 6817 9640 6851
rect 9588 6808 9640 6817
rect 4896 6604 4948 6656
rect 5356 6715 5408 6724
rect 5356 6681 5365 6715
rect 5365 6681 5399 6715
rect 5399 6681 5408 6715
rect 5356 6672 5408 6681
rect 6736 6672 6788 6724
rect 8024 6740 8076 6792
rect 8116 6740 8168 6792
rect 9772 6808 9824 6860
rect 7656 6604 7708 6656
rect 8024 6647 8076 6656
rect 8024 6613 8033 6647
rect 8033 6613 8067 6647
rect 8067 6613 8076 6647
rect 8024 6604 8076 6613
rect 8484 6604 8536 6656
rect 10324 6715 10376 6724
rect 10324 6681 10333 6715
rect 10333 6681 10367 6715
rect 10367 6681 10376 6715
rect 10324 6672 10376 6681
rect 10784 6647 10836 6656
rect 10784 6613 10793 6647
rect 10793 6613 10827 6647
rect 10827 6613 10836 6647
rect 10784 6604 10836 6613
rect 12624 6672 12676 6724
rect 26884 6715 26936 6724
rect 26884 6681 26893 6715
rect 26893 6681 26927 6715
rect 26927 6681 26936 6715
rect 26884 6672 26936 6681
rect 28356 6715 28408 6724
rect 28356 6681 28365 6715
rect 28365 6681 28399 6715
rect 28399 6681 28408 6715
rect 28356 6672 28408 6681
rect 22376 6604 22428 6656
rect 7896 6502 7948 6554
rect 7960 6502 8012 6554
rect 8024 6502 8076 6554
rect 8088 6502 8140 6554
rect 8152 6502 8204 6554
rect 14842 6502 14894 6554
rect 14906 6502 14958 6554
rect 14970 6502 15022 6554
rect 15034 6502 15086 6554
rect 15098 6502 15150 6554
rect 21788 6502 21840 6554
rect 21852 6502 21904 6554
rect 21916 6502 21968 6554
rect 21980 6502 22032 6554
rect 22044 6502 22096 6554
rect 28734 6502 28786 6554
rect 28798 6502 28850 6554
rect 28862 6502 28914 6554
rect 28926 6502 28978 6554
rect 28990 6502 29042 6554
rect 2228 6400 2280 6452
rect 3884 6400 3936 6452
rect 4344 6400 4396 6452
rect 5356 6443 5408 6452
rect 5356 6409 5365 6443
rect 5365 6409 5399 6443
rect 5399 6409 5408 6443
rect 5356 6400 5408 6409
rect 6368 6443 6420 6452
rect 6368 6409 6377 6443
rect 6377 6409 6411 6443
rect 6411 6409 6420 6443
rect 6368 6400 6420 6409
rect 7380 6400 7432 6452
rect 7656 6400 7708 6452
rect 7196 6332 7248 6384
rect 2228 6239 2280 6248
rect 2228 6205 2237 6239
rect 2237 6205 2271 6239
rect 2271 6205 2280 6239
rect 2228 6196 2280 6205
rect 3608 6264 3660 6316
rect 3700 6196 3752 6248
rect 5908 6307 5960 6316
rect 5908 6273 5917 6307
rect 5917 6273 5951 6307
rect 5951 6273 5960 6307
rect 5908 6264 5960 6273
rect 4252 6196 4304 6248
rect 5080 6196 5132 6248
rect 6644 6196 6696 6248
rect 4344 6128 4396 6180
rect 2780 6103 2832 6112
rect 2780 6069 2789 6103
rect 2789 6069 2823 6103
rect 2823 6069 2832 6103
rect 2780 6060 2832 6069
rect 3884 6103 3936 6112
rect 3884 6069 3893 6103
rect 3893 6069 3927 6103
rect 3927 6069 3936 6103
rect 3884 6060 3936 6069
rect 5908 6060 5960 6112
rect 8300 6400 8352 6452
rect 8944 6400 8996 6452
rect 9772 6400 9824 6452
rect 9864 6400 9916 6452
rect 10324 6400 10376 6452
rect 9036 6332 9088 6384
rect 9220 6196 9272 6248
rect 23756 6264 23808 6316
rect 24584 6264 24636 6316
rect 24676 6239 24728 6248
rect 24676 6205 24685 6239
rect 24685 6205 24719 6239
rect 24719 6205 24728 6239
rect 24676 6196 24728 6205
rect 26148 6239 26200 6248
rect 26148 6205 26157 6239
rect 26157 6205 26191 6239
rect 26191 6205 26200 6239
rect 26148 6196 26200 6205
rect 28632 6196 28684 6248
rect 7472 6103 7524 6112
rect 7472 6069 7481 6103
rect 7481 6069 7515 6103
rect 7515 6069 7524 6103
rect 7472 6060 7524 6069
rect 9496 6128 9548 6180
rect 24860 6128 24912 6180
rect 8576 6060 8628 6112
rect 10232 6060 10284 6112
rect 17224 6060 17276 6112
rect 23756 6103 23808 6112
rect 23756 6069 23765 6103
rect 23765 6069 23799 6103
rect 23799 6069 23808 6103
rect 23756 6060 23808 6069
rect 4423 5958 4475 6010
rect 4487 5958 4539 6010
rect 4551 5958 4603 6010
rect 4615 5958 4667 6010
rect 4679 5958 4731 6010
rect 11369 5958 11421 6010
rect 11433 5958 11485 6010
rect 11497 5958 11549 6010
rect 11561 5958 11613 6010
rect 11625 5958 11677 6010
rect 18315 5958 18367 6010
rect 18379 5958 18431 6010
rect 18443 5958 18495 6010
rect 18507 5958 18559 6010
rect 18571 5958 18623 6010
rect 25261 5958 25313 6010
rect 25325 5958 25377 6010
rect 25389 5958 25441 6010
rect 25453 5958 25505 6010
rect 25517 5958 25569 6010
rect 2964 5856 3016 5908
rect 3424 5856 3476 5908
rect 3884 5856 3936 5908
rect 6736 5856 6788 5908
rect 8300 5856 8352 5908
rect 8392 5856 8444 5908
rect 9036 5899 9088 5908
rect 9036 5865 9045 5899
rect 9045 5865 9079 5899
rect 9079 5865 9088 5899
rect 9036 5856 9088 5865
rect 9128 5856 9180 5908
rect 9864 5899 9916 5908
rect 9864 5865 9873 5899
rect 9873 5865 9907 5899
rect 9907 5865 9916 5899
rect 9864 5856 9916 5865
rect 10232 5899 10284 5908
rect 10232 5865 10241 5899
rect 10241 5865 10275 5899
rect 10275 5865 10284 5899
rect 10232 5856 10284 5865
rect 17224 5856 17276 5908
rect 26700 5856 26752 5908
rect 3332 5788 3384 5840
rect 6644 5788 6696 5840
rect 7840 5788 7892 5840
rect 7932 5831 7984 5840
rect 7932 5797 7941 5831
rect 7941 5797 7975 5831
rect 7975 5797 7984 5831
rect 7932 5788 7984 5797
rect 8024 5788 8076 5840
rect 11704 5788 11756 5840
rect 2596 5720 2648 5772
rect 3700 5720 3752 5772
rect 6000 5720 6052 5772
rect 1768 5652 1820 5704
rect 10232 5720 10284 5772
rect 14004 5720 14056 5772
rect 7472 5652 7524 5704
rect 7564 5652 7616 5704
rect 8668 5652 8720 5704
rect 9864 5652 9916 5704
rect 22836 5695 22888 5704
rect 22836 5661 22845 5695
rect 22845 5661 22879 5695
rect 22879 5661 22888 5695
rect 22836 5652 22888 5661
rect 26424 5763 26476 5772
rect 26424 5729 26433 5763
rect 26433 5729 26467 5763
rect 26467 5729 26476 5763
rect 26424 5720 26476 5729
rect 28816 5720 28868 5772
rect 4804 5584 4856 5636
rect 6000 5627 6052 5636
rect 6000 5593 6009 5627
rect 6009 5593 6043 5627
rect 6043 5593 6052 5627
rect 6000 5584 6052 5593
rect 6092 5627 6144 5636
rect 6092 5593 6101 5627
rect 6101 5593 6135 5627
rect 6135 5593 6144 5627
rect 6092 5584 6144 5593
rect 7104 5584 7156 5636
rect 4436 5516 4488 5568
rect 5816 5516 5868 5568
rect 9680 5516 9732 5568
rect 11796 5516 11848 5568
rect 27252 5584 27304 5636
rect 13084 5516 13136 5568
rect 7896 5414 7948 5466
rect 7960 5414 8012 5466
rect 8024 5414 8076 5466
rect 8088 5414 8140 5466
rect 8152 5414 8204 5466
rect 14842 5414 14894 5466
rect 14906 5414 14958 5466
rect 14970 5414 15022 5466
rect 15034 5414 15086 5466
rect 15098 5414 15150 5466
rect 21788 5414 21840 5466
rect 21852 5414 21904 5466
rect 21916 5414 21968 5466
rect 21980 5414 22032 5466
rect 22044 5414 22096 5466
rect 28734 5414 28786 5466
rect 28798 5414 28850 5466
rect 28862 5414 28914 5466
rect 28926 5414 28978 5466
rect 28990 5414 29042 5466
rect 664 5312 716 5364
rect 3056 5355 3108 5364
rect 3056 5321 3065 5355
rect 3065 5321 3099 5355
rect 3099 5321 3108 5355
rect 3056 5312 3108 5321
rect 3700 5312 3752 5364
rect 4252 5312 4304 5364
rect 5448 5355 5500 5364
rect 5448 5321 5457 5355
rect 5457 5321 5491 5355
rect 5491 5321 5500 5355
rect 5448 5312 5500 5321
rect 3332 5244 3384 5296
rect 6092 5312 6144 5364
rect 6460 5355 6512 5364
rect 6460 5321 6469 5355
rect 6469 5321 6503 5355
rect 6503 5321 6512 5355
rect 6460 5312 6512 5321
rect 388 5176 440 5228
rect 1584 5219 1636 5228
rect 1584 5185 1593 5219
rect 1593 5185 1627 5219
rect 1627 5185 1636 5219
rect 1584 5176 1636 5185
rect 2136 5176 2188 5228
rect 3976 5176 4028 5228
rect 6000 5244 6052 5296
rect 7748 5287 7800 5296
rect 7748 5253 7757 5287
rect 7757 5253 7791 5287
rect 7791 5253 7800 5287
rect 7748 5244 7800 5253
rect 8484 5312 8536 5364
rect 8760 5312 8812 5364
rect 9036 5312 9088 5364
rect 24584 5312 24636 5364
rect 26700 5355 26752 5364
rect 26700 5321 26709 5355
rect 26709 5321 26743 5355
rect 26743 5321 26752 5355
rect 26700 5312 26752 5321
rect 9864 5287 9916 5296
rect 6552 5219 6604 5228
rect 1952 5151 2004 5160
rect 1952 5117 1961 5151
rect 1961 5117 1995 5151
rect 1995 5117 2004 5151
rect 1952 5108 2004 5117
rect 4988 5151 5040 5160
rect 4988 5117 4997 5151
rect 4997 5117 5031 5151
rect 5031 5117 5040 5151
rect 4988 5108 5040 5117
rect 5356 5108 5408 5160
rect 6552 5185 6561 5219
rect 6561 5185 6595 5219
rect 6595 5185 6604 5219
rect 6552 5176 6604 5185
rect 6092 5151 6144 5160
rect 6092 5117 6101 5151
rect 6101 5117 6135 5151
rect 6135 5117 6144 5151
rect 6092 5108 6144 5117
rect 7840 5151 7892 5160
rect 7840 5117 7849 5151
rect 7849 5117 7883 5151
rect 7883 5117 7892 5151
rect 7840 5108 7892 5117
rect 8254 5176 8306 5228
rect 8392 5219 8444 5228
rect 8392 5185 8401 5219
rect 8401 5185 8435 5219
rect 8435 5185 8444 5219
rect 8392 5176 8444 5185
rect 8484 5219 8536 5228
rect 8484 5185 8493 5219
rect 8493 5185 8527 5219
rect 8527 5185 8536 5219
rect 8484 5176 8536 5185
rect 8944 5219 8996 5228
rect 8944 5185 8953 5219
rect 8953 5185 8987 5219
rect 8987 5185 8996 5219
rect 8944 5176 8996 5185
rect 9220 5219 9272 5228
rect 9220 5185 9229 5219
rect 9229 5185 9263 5219
rect 9263 5185 9272 5219
rect 9220 5176 9272 5185
rect 9864 5253 9873 5287
rect 9873 5253 9907 5287
rect 9907 5253 9916 5287
rect 9864 5244 9916 5253
rect 14464 5244 14516 5296
rect 17408 5176 17460 5228
rect 23480 5219 23532 5228
rect 23480 5185 23489 5219
rect 23489 5185 23523 5219
rect 23523 5185 23532 5219
rect 23480 5176 23532 5185
rect 24860 5219 24912 5228
rect 24860 5185 24869 5219
rect 24869 5185 24903 5219
rect 24903 5185 24912 5219
rect 24860 5176 24912 5185
rect 10968 5108 11020 5160
rect 8116 5040 8168 5092
rect 2504 5015 2556 5024
rect 2504 4981 2513 5015
rect 2513 4981 2547 5015
rect 2547 4981 2556 5015
rect 2504 4972 2556 4981
rect 2688 4972 2740 5024
rect 4896 4972 4948 5024
rect 6644 5015 6696 5024
rect 6644 4981 6653 5015
rect 6653 4981 6687 5015
rect 6687 4981 6696 5015
rect 6644 4972 6696 4981
rect 8208 5015 8260 5024
rect 8208 4981 8217 5015
rect 8217 4981 8251 5015
rect 8251 4981 8260 5015
rect 8208 4972 8260 4981
rect 8576 4972 8628 5024
rect 8852 4972 8904 5024
rect 10784 4972 10836 5024
rect 11152 4972 11204 5024
rect 24768 5108 24820 5160
rect 25964 5108 26016 5160
rect 26516 5040 26568 5092
rect 28080 4972 28132 5024
rect 4423 4870 4475 4922
rect 4487 4870 4539 4922
rect 4551 4870 4603 4922
rect 4615 4870 4667 4922
rect 4679 4870 4731 4922
rect 11369 4870 11421 4922
rect 11433 4870 11485 4922
rect 11497 4870 11549 4922
rect 11561 4870 11613 4922
rect 11625 4870 11677 4922
rect 18315 4870 18367 4922
rect 18379 4870 18431 4922
rect 18443 4870 18495 4922
rect 18507 4870 18559 4922
rect 18571 4870 18623 4922
rect 25261 4870 25313 4922
rect 25325 4870 25377 4922
rect 25389 4870 25441 4922
rect 25453 4870 25505 4922
rect 25517 4870 25569 4922
rect 2228 4768 2280 4820
rect 3976 4811 4028 4820
rect 3976 4777 3985 4811
rect 3985 4777 4019 4811
rect 4019 4777 4028 4811
rect 3976 4768 4028 4777
rect 4068 4768 4120 4820
rect 5172 4768 5224 4820
rect 5540 4768 5592 4820
rect 3516 4700 3568 4752
rect 4344 4743 4396 4752
rect 4344 4709 4353 4743
rect 4353 4709 4387 4743
rect 4387 4709 4396 4743
rect 4344 4700 4396 4709
rect 1216 4632 1268 4684
rect 1308 4564 1360 4616
rect 3976 4632 4028 4684
rect 5356 4632 5408 4684
rect 5816 4675 5868 4684
rect 5816 4641 5825 4675
rect 5825 4641 5859 4675
rect 5859 4641 5868 4675
rect 5816 4632 5868 4641
rect 8024 4700 8076 4752
rect 9404 4811 9456 4820
rect 9404 4777 9413 4811
rect 9413 4777 9447 4811
rect 9447 4777 9456 4811
rect 9404 4768 9456 4777
rect 9864 4768 9916 4820
rect 12440 4768 12492 4820
rect 22928 4768 22980 4820
rect 6644 4632 6696 4684
rect 7104 4632 7156 4684
rect 12348 4700 12400 4752
rect 12624 4700 12676 4752
rect 19248 4700 19300 4752
rect 3884 4564 3936 4616
rect 4068 4564 4120 4616
rect 5264 4564 5316 4616
rect 5908 4564 5960 4616
rect 6736 4607 6788 4616
rect 6736 4573 6745 4607
rect 6745 4573 6779 4607
rect 6779 4573 6788 4607
rect 6736 4564 6788 4573
rect 9036 4632 9088 4684
rect 10784 4632 10836 4684
rect 16120 4632 16172 4684
rect 20904 4632 20956 4684
rect 9404 4564 9456 4616
rect 9680 4564 9732 4616
rect 16488 4564 16540 4616
rect 22928 4564 22980 4616
rect 1492 4428 1544 4480
rect 7104 4496 7156 4548
rect 8760 4496 8812 4548
rect 9312 4471 9364 4480
rect 9312 4437 9321 4471
rect 9321 4437 9355 4471
rect 9355 4437 9364 4471
rect 9312 4428 9364 4437
rect 22560 4539 22612 4548
rect 22560 4505 22569 4539
rect 22569 4505 22603 4539
rect 22603 4505 22612 4539
rect 22560 4496 22612 4505
rect 24860 4496 24912 4548
rect 11152 4428 11204 4480
rect 12072 4428 12124 4480
rect 23664 4428 23716 4480
rect 25136 4632 25188 4684
rect 25872 4607 25924 4616
rect 25872 4573 25881 4607
rect 25881 4573 25915 4607
rect 25915 4573 25924 4607
rect 25872 4564 25924 4573
rect 7896 4326 7948 4378
rect 7960 4326 8012 4378
rect 8024 4326 8076 4378
rect 8088 4326 8140 4378
rect 8152 4326 8204 4378
rect 14842 4326 14894 4378
rect 14906 4326 14958 4378
rect 14970 4326 15022 4378
rect 15034 4326 15086 4378
rect 15098 4326 15150 4378
rect 21788 4326 21840 4378
rect 21852 4326 21904 4378
rect 21916 4326 21968 4378
rect 21980 4326 22032 4378
rect 22044 4326 22096 4378
rect 28734 4326 28786 4378
rect 28798 4326 28850 4378
rect 28862 4326 28914 4378
rect 28926 4326 28978 4378
rect 28990 4326 29042 4378
rect 1584 4224 1636 4276
rect 2504 4224 2556 4276
rect 848 4156 900 4208
rect 1308 4156 1360 4208
rect 3148 4156 3200 4208
rect 1584 4131 1636 4140
rect 1584 4097 1593 4131
rect 1593 4097 1627 4131
rect 1627 4097 1636 4131
rect 1584 4088 1636 4097
rect 2320 4131 2372 4140
rect 2320 4097 2329 4131
rect 2329 4097 2363 4131
rect 2363 4097 2372 4131
rect 2320 4088 2372 4097
rect 2320 3884 2372 3936
rect 3700 4020 3752 4072
rect 4160 4088 4212 4140
rect 6184 4156 6236 4208
rect 5448 4088 5500 4140
rect 5632 4088 5684 4140
rect 5816 4131 5868 4140
rect 5816 4097 5825 4131
rect 5825 4097 5859 4131
rect 5859 4097 5868 4131
rect 5816 4088 5868 4097
rect 8576 4156 8628 4208
rect 9220 4267 9272 4276
rect 9220 4233 9229 4267
rect 9229 4233 9263 4267
rect 9263 4233 9272 4267
rect 9220 4224 9272 4233
rect 9312 4224 9364 4276
rect 9680 4156 9732 4208
rect 9772 4156 9824 4208
rect 9864 4199 9916 4208
rect 9864 4165 9873 4199
rect 9873 4165 9907 4199
rect 9907 4165 9916 4199
rect 9864 4156 9916 4165
rect 10784 4199 10836 4208
rect 10784 4165 10793 4199
rect 10793 4165 10827 4199
rect 10827 4165 10836 4199
rect 10784 4156 10836 4165
rect 22560 4224 22612 4276
rect 28356 4224 28408 4276
rect 23296 4156 23348 4208
rect 5172 3952 5224 4004
rect 9312 4131 9364 4140
rect 9312 4097 9321 4131
rect 9321 4097 9355 4131
rect 9355 4097 9364 4131
rect 9312 4088 9364 4097
rect 6828 3952 6880 4004
rect 8300 3952 8352 4004
rect 8760 3952 8812 4004
rect 10232 4131 10284 4140
rect 10232 4097 10241 4131
rect 10241 4097 10275 4131
rect 10275 4097 10284 4131
rect 10232 4088 10284 4097
rect 10048 4020 10100 4072
rect 11336 4088 11388 4140
rect 22376 4131 22428 4140
rect 22376 4097 22385 4131
rect 22385 4097 22419 4131
rect 22419 4097 22428 4131
rect 22376 4088 22428 4097
rect 23848 4131 23900 4140
rect 23848 4097 23857 4131
rect 23857 4097 23891 4131
rect 23891 4097 23900 4131
rect 23848 4088 23900 4097
rect 24124 4088 24176 4140
rect 26608 4088 26660 4140
rect 27160 4131 27212 4140
rect 27160 4097 27169 4131
rect 27169 4097 27203 4131
rect 27203 4097 27212 4131
rect 27160 4088 27212 4097
rect 10692 4020 10744 4072
rect 3056 3884 3108 3936
rect 4252 3884 4304 3936
rect 4988 3884 5040 3936
rect 5908 3884 5960 3936
rect 9588 3884 9640 3936
rect 10140 3884 10192 3936
rect 10508 3952 10560 4004
rect 12072 3952 12124 4004
rect 22284 4020 22336 4072
rect 23112 4020 23164 4072
rect 10600 3884 10652 3936
rect 11888 3884 11940 3936
rect 23756 3884 23808 3936
rect 23940 3952 23992 4004
rect 25136 3952 25188 4004
rect 25596 3884 25648 3936
rect 4423 3782 4475 3834
rect 4487 3782 4539 3834
rect 4551 3782 4603 3834
rect 4615 3782 4667 3834
rect 4679 3782 4731 3834
rect 11369 3782 11421 3834
rect 11433 3782 11485 3834
rect 11497 3782 11549 3834
rect 11561 3782 11613 3834
rect 11625 3782 11677 3834
rect 18315 3782 18367 3834
rect 18379 3782 18431 3834
rect 18443 3782 18495 3834
rect 18507 3782 18559 3834
rect 18571 3782 18623 3834
rect 25261 3782 25313 3834
rect 25325 3782 25377 3834
rect 25389 3782 25441 3834
rect 25453 3782 25505 3834
rect 25517 3782 25569 3834
rect 2688 3680 2740 3732
rect 3056 3680 3108 3732
rect 4528 3680 4580 3732
rect 4988 3680 5040 3732
rect 7748 3680 7800 3732
rect 8484 3680 8536 3732
rect 8852 3680 8904 3732
rect 10232 3680 10284 3732
rect 10876 3680 10928 3732
rect 10968 3680 11020 3732
rect 11888 3723 11940 3732
rect 11888 3689 11897 3723
rect 11897 3689 11931 3723
rect 11931 3689 11940 3723
rect 11888 3680 11940 3689
rect 12072 3680 12124 3732
rect 24124 3723 24176 3732
rect 24124 3689 24133 3723
rect 24133 3689 24167 3723
rect 24167 3689 24176 3723
rect 24124 3680 24176 3689
rect 27160 3680 27212 3732
rect 4068 3544 4120 3596
rect 5908 3544 5960 3596
rect 2596 3476 2648 3528
rect 2780 3476 2832 3528
rect 3332 3476 3384 3528
rect 3884 3476 3936 3528
rect 1584 3408 1636 3460
rect 2044 3383 2096 3392
rect 2044 3349 2053 3383
rect 2053 3349 2087 3383
rect 2087 3349 2096 3383
rect 2044 3340 2096 3349
rect 2872 3408 2924 3460
rect 3056 3408 3108 3460
rect 4528 3451 4580 3460
rect 4528 3417 4537 3451
rect 4537 3417 4571 3451
rect 4571 3417 4580 3451
rect 4528 3408 4580 3417
rect 4804 3519 4856 3528
rect 4804 3485 4813 3519
rect 4813 3485 4847 3519
rect 4847 3485 4856 3519
rect 4804 3476 4856 3485
rect 10048 3612 10100 3664
rect 20352 3612 20404 3664
rect 21456 3612 21508 3664
rect 3884 3340 3936 3392
rect 4896 3340 4948 3392
rect 7104 3476 7156 3528
rect 7472 3519 7524 3528
rect 7472 3485 7481 3519
rect 7481 3485 7515 3519
rect 7515 3485 7524 3519
rect 7472 3476 7524 3485
rect 7656 3476 7708 3528
rect 7932 3519 7984 3528
rect 7932 3485 7941 3519
rect 7941 3485 7975 3519
rect 7975 3485 7984 3519
rect 7932 3476 7984 3485
rect 9588 3476 9640 3528
rect 7196 3408 7248 3460
rect 10968 3519 11020 3528
rect 10968 3485 10977 3519
rect 10977 3485 11011 3519
rect 11011 3485 11020 3519
rect 10968 3476 11020 3485
rect 11336 3476 11388 3528
rect 11152 3408 11204 3460
rect 20076 3519 20128 3528
rect 20076 3485 20085 3519
rect 20085 3485 20119 3519
rect 20119 3485 20128 3519
rect 20076 3476 20128 3485
rect 22836 3544 22888 3596
rect 24400 3519 24452 3528
rect 24400 3485 24409 3519
rect 24409 3485 24443 3519
rect 24443 3485 24452 3519
rect 24400 3476 24452 3485
rect 8760 3340 8812 3392
rect 10416 3340 10468 3392
rect 10508 3340 10560 3392
rect 10784 3383 10836 3392
rect 10784 3349 10793 3383
rect 10793 3349 10827 3383
rect 10827 3349 10836 3383
rect 10784 3340 10836 3349
rect 11060 3383 11112 3392
rect 11060 3349 11069 3383
rect 11069 3349 11103 3383
rect 11103 3349 11112 3383
rect 11060 3340 11112 3349
rect 24216 3408 24268 3460
rect 25872 3519 25924 3528
rect 25872 3485 25881 3519
rect 25881 3485 25915 3519
rect 25915 3485 25924 3519
rect 25872 3476 25924 3485
rect 29460 3476 29512 3528
rect 27068 3340 27120 3392
rect 7896 3238 7948 3290
rect 7960 3238 8012 3290
rect 8024 3238 8076 3290
rect 8088 3238 8140 3290
rect 8152 3238 8204 3290
rect 14842 3238 14894 3290
rect 14906 3238 14958 3290
rect 14970 3238 15022 3290
rect 15034 3238 15086 3290
rect 15098 3238 15150 3290
rect 21788 3238 21840 3290
rect 21852 3238 21904 3290
rect 21916 3238 21968 3290
rect 21980 3238 22032 3290
rect 22044 3238 22096 3290
rect 28734 3238 28786 3290
rect 28798 3238 28850 3290
rect 28862 3238 28914 3290
rect 28926 3238 28978 3290
rect 28990 3238 29042 3290
rect 1952 3136 2004 3188
rect 2320 3136 2372 3188
rect 5448 3136 5500 3188
rect 1860 2932 1912 2984
rect 2872 2975 2924 2984
rect 2872 2941 2881 2975
rect 2881 2941 2915 2975
rect 2915 2941 2924 2975
rect 2872 2932 2924 2941
rect 3056 3043 3108 3052
rect 3056 3009 3065 3043
rect 3065 3009 3099 3043
rect 3099 3009 3108 3043
rect 3056 3000 3108 3009
rect 3700 3000 3752 3052
rect 3884 3043 3936 3052
rect 3884 3009 3893 3043
rect 3893 3009 3927 3043
rect 3927 3009 3936 3043
rect 3884 3000 3936 3009
rect 6184 3111 6236 3120
rect 6184 3077 6193 3111
rect 6193 3077 6227 3111
rect 6227 3077 6236 3111
rect 6184 3068 6236 3077
rect 7564 3179 7616 3188
rect 7564 3145 7573 3179
rect 7573 3145 7607 3179
rect 7607 3145 7616 3179
rect 7564 3136 7616 3145
rect 8392 3136 8444 3188
rect 9404 3136 9456 3188
rect 9312 3068 9364 3120
rect 4068 3000 4120 3052
rect 6552 3043 6604 3052
rect 6552 3009 6561 3043
rect 6561 3009 6595 3043
rect 6595 3009 6604 3043
rect 6552 3000 6604 3009
rect 7472 3000 7524 3052
rect 10140 3136 10192 3188
rect 10416 3136 10468 3188
rect 10508 3136 10560 3188
rect 11244 3136 11296 3188
rect 11888 3136 11940 3188
rect 11980 3136 12032 3188
rect 12348 3179 12400 3188
rect 12348 3145 12357 3179
rect 12357 3145 12391 3179
rect 12391 3145 12400 3179
rect 12348 3136 12400 3145
rect 9956 3068 10008 3120
rect 10784 3000 10836 3052
rect 11704 3043 11756 3052
rect 11704 3009 11713 3043
rect 11713 3009 11747 3043
rect 11747 3009 11756 3043
rect 11704 3000 11756 3009
rect 7380 2932 7432 2984
rect 8208 2932 8260 2984
rect 8760 2932 8812 2984
rect 9220 2975 9272 2984
rect 9220 2941 9229 2975
rect 9229 2941 9263 2975
rect 9263 2941 9272 2975
rect 9220 2932 9272 2941
rect 9496 2932 9548 2984
rect 10140 2932 10192 2984
rect 10600 2932 10652 2984
rect 6736 2907 6788 2916
rect 6736 2873 6745 2907
rect 6745 2873 6779 2907
rect 6779 2873 6788 2907
rect 6736 2864 6788 2873
rect 9680 2864 9732 2916
rect 12256 3043 12308 3052
rect 12256 3009 12265 3043
rect 12265 3009 12299 3043
rect 12299 3009 12308 3043
rect 12256 3000 12308 3009
rect 23388 3136 23440 3188
rect 15844 3000 15896 3052
rect 18880 3000 18932 3052
rect 21824 3043 21876 3052
rect 21824 3009 21833 3043
rect 21833 3009 21867 3043
rect 21867 3009 21876 3043
rect 21824 3000 21876 3009
rect 26792 3068 26844 3120
rect 23296 3043 23348 3052
rect 23296 3009 23305 3043
rect 23305 3009 23339 3043
rect 23339 3009 23348 3043
rect 23296 3000 23348 3009
rect 21364 2864 21416 2916
rect 22560 2932 22612 2984
rect 24952 3043 25004 3052
rect 24952 3009 24961 3043
rect 24961 3009 24995 3043
rect 24995 3009 25004 3043
rect 24952 3000 25004 3009
rect 26976 3043 27028 3052
rect 26976 3009 26985 3043
rect 26985 3009 27019 3043
rect 27019 3009 27028 3043
rect 26976 3000 27028 3009
rect 1768 2796 1820 2848
rect 3792 2796 3844 2848
rect 4252 2796 4304 2848
rect 4804 2796 4856 2848
rect 8300 2796 8352 2848
rect 11336 2796 11388 2848
rect 21548 2796 21600 2848
rect 24676 2864 24728 2916
rect 4423 2694 4475 2746
rect 4487 2694 4539 2746
rect 4551 2694 4603 2746
rect 4615 2694 4667 2746
rect 4679 2694 4731 2746
rect 11369 2694 11421 2746
rect 11433 2694 11485 2746
rect 11497 2694 11549 2746
rect 11561 2694 11613 2746
rect 11625 2694 11677 2746
rect 18315 2694 18367 2746
rect 18379 2694 18431 2746
rect 18443 2694 18495 2746
rect 18507 2694 18559 2746
rect 18571 2694 18623 2746
rect 25261 2694 25313 2746
rect 25325 2694 25377 2746
rect 25389 2694 25441 2746
rect 25453 2694 25505 2746
rect 25517 2694 25569 2746
rect 6276 2592 6328 2644
rect 7012 2592 7064 2644
rect 9680 2592 9732 2644
rect 10508 2592 10560 2644
rect 11704 2592 11756 2644
rect 12164 2592 12216 2644
rect 12532 2635 12584 2644
rect 12532 2601 12541 2635
rect 12541 2601 12575 2635
rect 12575 2601 12584 2635
rect 12532 2592 12584 2601
rect 2320 2499 2372 2508
rect 2320 2465 2329 2499
rect 2329 2465 2363 2499
rect 2363 2465 2372 2499
rect 2320 2456 2372 2465
rect 2596 2456 2648 2508
rect 7104 2524 7156 2576
rect 10968 2524 11020 2576
rect 3056 2431 3108 2440
rect 3056 2397 3065 2431
rect 3065 2397 3099 2431
rect 3099 2397 3108 2431
rect 3056 2388 3108 2397
rect 5356 2388 5408 2440
rect 6184 2499 6236 2508
rect 6184 2465 6193 2499
rect 6193 2465 6227 2499
rect 6227 2465 6236 2499
rect 6184 2456 6236 2465
rect 6276 2388 6328 2440
rect 2136 2295 2188 2304
rect 2136 2261 2145 2295
rect 2145 2261 2179 2295
rect 2179 2261 2188 2295
rect 2136 2252 2188 2261
rect 2872 2295 2924 2304
rect 2872 2261 2881 2295
rect 2881 2261 2915 2295
rect 2915 2261 2924 2295
rect 2872 2252 2924 2261
rect 3608 2295 3660 2304
rect 3608 2261 3617 2295
rect 3617 2261 3651 2295
rect 3651 2261 3660 2295
rect 3608 2252 3660 2261
rect 8484 2388 8536 2440
rect 8852 2388 8904 2440
rect 9496 2456 9548 2508
rect 9864 2388 9916 2440
rect 10692 2388 10744 2440
rect 10784 2431 10836 2440
rect 10784 2397 10793 2431
rect 10793 2397 10827 2431
rect 10827 2397 10836 2431
rect 10784 2388 10836 2397
rect 11060 2388 11112 2440
rect 11244 2388 11296 2440
rect 13084 2524 13136 2576
rect 20720 2499 20772 2508
rect 20720 2465 20729 2499
rect 20729 2465 20763 2499
rect 20763 2465 20772 2499
rect 20720 2456 20772 2465
rect 21180 2456 21232 2508
rect 13268 2431 13320 2440
rect 13268 2397 13277 2431
rect 13277 2397 13311 2431
rect 13311 2397 13320 2431
rect 13268 2388 13320 2397
rect 17684 2431 17736 2440
rect 17684 2397 17693 2431
rect 17693 2397 17727 2431
rect 17727 2397 17736 2431
rect 17684 2388 17736 2397
rect 7656 2320 7708 2372
rect 5264 2252 5316 2304
rect 8944 2252 8996 2304
rect 18880 2363 18932 2372
rect 18880 2329 18889 2363
rect 18889 2329 18923 2363
rect 18923 2329 18932 2363
rect 18880 2320 18932 2329
rect 11980 2252 12032 2304
rect 13084 2295 13136 2304
rect 13084 2261 13093 2295
rect 13093 2261 13127 2295
rect 13127 2261 13136 2295
rect 13084 2252 13136 2261
rect 15200 2252 15252 2304
rect 20352 2388 20404 2440
rect 24584 2456 24636 2508
rect 23388 2320 23440 2372
rect 26240 2252 26292 2304
rect 7896 2150 7948 2202
rect 7960 2150 8012 2202
rect 8024 2150 8076 2202
rect 8088 2150 8140 2202
rect 8152 2150 8204 2202
rect 14842 2150 14894 2202
rect 14906 2150 14958 2202
rect 14970 2150 15022 2202
rect 15034 2150 15086 2202
rect 15098 2150 15150 2202
rect 21788 2150 21840 2202
rect 21852 2150 21904 2202
rect 21916 2150 21968 2202
rect 21980 2150 22032 2202
rect 22044 2150 22096 2202
rect 28734 2150 28786 2202
rect 28798 2150 28850 2202
rect 28862 2150 28914 2202
rect 28926 2150 28978 2202
rect 28990 2150 29042 2202
rect 5356 2048 5408 2100
rect 6552 2048 6604 2100
rect 13084 2048 13136 2100
rect 18880 2048 18932 2100
rect 3056 1980 3108 2032
rect 6000 1980 6052 2032
rect 6184 1980 6236 2032
rect 10876 1980 10928 2032
rect 2320 1912 2372 1964
rect 5724 1912 5776 1964
rect 2412 1844 2464 1896
rect 25596 2048 25648 2100
rect 26424 2048 26476 2100
rect 27252 2048 27304 2100
rect 27804 2048 27856 2100
rect 28908 1980 28960 2032
rect 14648 1912 14700 1964
rect 26240 1912 26292 1964
rect 24860 1844 24912 1896
rect 26424 1844 26476 1896
rect 3608 1776 3660 1828
rect 10968 1708 11020 1760
rect 2136 1640 2188 1692
rect 8668 1640 8720 1692
rect 2872 1504 2924 1556
rect 11152 1504 11204 1556
rect 24584 1504 24636 1556
rect 22008 1368 22060 1420
<< metal2 >>
rect 4423 27772 4731 27781
rect 4423 27770 4429 27772
rect 4485 27770 4509 27772
rect 4565 27770 4589 27772
rect 4645 27770 4669 27772
rect 4725 27770 4731 27772
rect 4485 27718 4487 27770
rect 4667 27718 4669 27770
rect 4423 27716 4429 27718
rect 4485 27716 4509 27718
rect 4565 27716 4589 27718
rect 4645 27716 4669 27718
rect 4725 27716 4731 27718
rect 4423 27707 4731 27716
rect 11369 27772 11677 27781
rect 11369 27770 11375 27772
rect 11431 27770 11455 27772
rect 11511 27770 11535 27772
rect 11591 27770 11615 27772
rect 11671 27770 11677 27772
rect 11431 27718 11433 27770
rect 11613 27718 11615 27770
rect 11369 27716 11375 27718
rect 11431 27716 11455 27718
rect 11511 27716 11535 27718
rect 11591 27716 11615 27718
rect 11671 27716 11677 27718
rect 11369 27707 11677 27716
rect 18315 27772 18623 27781
rect 18315 27770 18321 27772
rect 18377 27770 18401 27772
rect 18457 27770 18481 27772
rect 18537 27770 18561 27772
rect 18617 27770 18623 27772
rect 18377 27718 18379 27770
rect 18559 27718 18561 27770
rect 18315 27716 18321 27718
rect 18377 27716 18401 27718
rect 18457 27716 18481 27718
rect 18537 27716 18561 27718
rect 18617 27716 18623 27718
rect 18315 27707 18623 27716
rect 25261 27772 25569 27781
rect 25261 27770 25267 27772
rect 25323 27770 25347 27772
rect 25403 27770 25427 27772
rect 25483 27770 25507 27772
rect 25563 27770 25569 27772
rect 25323 27718 25325 27770
rect 25505 27718 25507 27770
rect 25261 27716 25267 27718
rect 25323 27716 25347 27718
rect 25403 27716 25427 27718
rect 25483 27716 25507 27718
rect 25563 27716 25569 27718
rect 25261 27707 25569 27716
rect 28538 27568 28594 27577
rect 28538 27503 28540 27512
rect 28592 27503 28594 27512
rect 28540 27474 28592 27480
rect 7896 27228 8204 27237
rect 7896 27226 7902 27228
rect 7958 27226 7982 27228
rect 8038 27226 8062 27228
rect 8118 27226 8142 27228
rect 8198 27226 8204 27228
rect 7958 27174 7960 27226
rect 8140 27174 8142 27226
rect 7896 27172 7902 27174
rect 7958 27172 7982 27174
rect 8038 27172 8062 27174
rect 8118 27172 8142 27174
rect 8198 27172 8204 27174
rect 7896 27163 8204 27172
rect 14842 27228 15150 27237
rect 14842 27226 14848 27228
rect 14904 27226 14928 27228
rect 14984 27226 15008 27228
rect 15064 27226 15088 27228
rect 15144 27226 15150 27228
rect 14904 27174 14906 27226
rect 15086 27174 15088 27226
rect 14842 27172 14848 27174
rect 14904 27172 14928 27174
rect 14984 27172 15008 27174
rect 15064 27172 15088 27174
rect 15144 27172 15150 27174
rect 14842 27163 15150 27172
rect 21788 27228 22096 27237
rect 21788 27226 21794 27228
rect 21850 27226 21874 27228
rect 21930 27226 21954 27228
rect 22010 27226 22034 27228
rect 22090 27226 22096 27228
rect 21850 27174 21852 27226
rect 22032 27174 22034 27226
rect 21788 27172 21794 27174
rect 21850 27172 21874 27174
rect 21930 27172 21954 27174
rect 22010 27172 22034 27174
rect 22090 27172 22096 27174
rect 21788 27163 22096 27172
rect 28734 27228 29042 27237
rect 28734 27226 28740 27228
rect 28796 27226 28820 27228
rect 28876 27226 28900 27228
rect 28956 27226 28980 27228
rect 29036 27226 29042 27228
rect 28796 27174 28798 27226
rect 28978 27174 28980 27226
rect 28734 27172 28740 27174
rect 28796 27172 28820 27174
rect 28876 27172 28900 27174
rect 28956 27172 28980 27174
rect 29036 27172 29042 27174
rect 28734 27163 29042 27172
rect 28356 26920 28408 26926
rect 28356 26862 28408 26868
rect 22744 26784 22796 26790
rect 28368 26761 28396 26862
rect 22744 26726 22796 26732
rect 28354 26752 28410 26761
rect 4423 26684 4731 26693
rect 4423 26682 4429 26684
rect 4485 26682 4509 26684
rect 4565 26682 4589 26684
rect 4645 26682 4669 26684
rect 4725 26682 4731 26684
rect 4485 26630 4487 26682
rect 4667 26630 4669 26682
rect 4423 26628 4429 26630
rect 4485 26628 4509 26630
rect 4565 26628 4589 26630
rect 4645 26628 4669 26630
rect 4725 26628 4731 26630
rect 4423 26619 4731 26628
rect 11369 26684 11677 26693
rect 11369 26682 11375 26684
rect 11431 26682 11455 26684
rect 11511 26682 11535 26684
rect 11591 26682 11615 26684
rect 11671 26682 11677 26684
rect 11431 26630 11433 26682
rect 11613 26630 11615 26682
rect 11369 26628 11375 26630
rect 11431 26628 11455 26630
rect 11511 26628 11535 26630
rect 11591 26628 11615 26630
rect 11671 26628 11677 26630
rect 11369 26619 11677 26628
rect 18315 26684 18623 26693
rect 18315 26682 18321 26684
rect 18377 26682 18401 26684
rect 18457 26682 18481 26684
rect 18537 26682 18561 26684
rect 18617 26682 18623 26684
rect 18377 26630 18379 26682
rect 18559 26630 18561 26682
rect 18315 26628 18321 26630
rect 18377 26628 18401 26630
rect 18457 26628 18481 26630
rect 18537 26628 18561 26630
rect 18617 26628 18623 26630
rect 18315 26619 18623 26628
rect 14280 26308 14332 26314
rect 14280 26250 14332 26256
rect 7896 26140 8204 26149
rect 7896 26138 7902 26140
rect 7958 26138 7982 26140
rect 8038 26138 8062 26140
rect 8118 26138 8142 26140
rect 8198 26138 8204 26140
rect 7958 26086 7960 26138
rect 8140 26086 8142 26138
rect 7896 26084 7902 26086
rect 7958 26084 7982 26086
rect 8038 26084 8062 26086
rect 8118 26084 8142 26086
rect 8198 26084 8204 26086
rect 7896 26075 8204 26084
rect 4423 25596 4731 25605
rect 4423 25594 4429 25596
rect 4485 25594 4509 25596
rect 4565 25594 4589 25596
rect 4645 25594 4669 25596
rect 4725 25594 4731 25596
rect 4485 25542 4487 25594
rect 4667 25542 4669 25594
rect 4423 25540 4429 25542
rect 4485 25540 4509 25542
rect 4565 25540 4589 25542
rect 4645 25540 4669 25542
rect 4725 25540 4731 25542
rect 4423 25531 4731 25540
rect 11369 25596 11677 25605
rect 11369 25594 11375 25596
rect 11431 25594 11455 25596
rect 11511 25594 11535 25596
rect 11591 25594 11615 25596
rect 11671 25594 11677 25596
rect 11431 25542 11433 25594
rect 11613 25542 11615 25594
rect 11369 25540 11375 25542
rect 11431 25540 11455 25542
rect 11511 25540 11535 25542
rect 11591 25540 11615 25542
rect 11671 25540 11677 25542
rect 11369 25531 11677 25540
rect 7896 25052 8204 25061
rect 7896 25050 7902 25052
rect 7958 25050 7982 25052
rect 8038 25050 8062 25052
rect 8118 25050 8142 25052
rect 8198 25050 8204 25052
rect 7958 24998 7960 25050
rect 8140 24998 8142 25050
rect 7896 24996 7902 24998
rect 7958 24996 7982 24998
rect 8038 24996 8062 24998
rect 8118 24996 8142 24998
rect 8198 24996 8204 24998
rect 7896 24987 8204 24996
rect 12808 24608 12860 24614
rect 12808 24550 12860 24556
rect 4423 24508 4731 24517
rect 4423 24506 4429 24508
rect 4485 24506 4509 24508
rect 4565 24506 4589 24508
rect 4645 24506 4669 24508
rect 4725 24506 4731 24508
rect 4485 24454 4487 24506
rect 4667 24454 4669 24506
rect 4423 24452 4429 24454
rect 4485 24452 4509 24454
rect 4565 24452 4589 24454
rect 4645 24452 4669 24454
rect 4725 24452 4731 24454
rect 4423 24443 4731 24452
rect 11369 24508 11677 24517
rect 11369 24506 11375 24508
rect 11431 24506 11455 24508
rect 11511 24506 11535 24508
rect 11591 24506 11615 24508
rect 11671 24506 11677 24508
rect 11431 24454 11433 24506
rect 11613 24454 11615 24506
rect 11369 24452 11375 24454
rect 11431 24452 11455 24454
rect 11511 24452 11535 24454
rect 11591 24452 11615 24454
rect 11671 24452 11677 24454
rect 11369 24443 11677 24452
rect 7896 23964 8204 23973
rect 7896 23962 7902 23964
rect 7958 23962 7982 23964
rect 8038 23962 8062 23964
rect 8118 23962 8142 23964
rect 8198 23962 8204 23964
rect 7958 23910 7960 23962
rect 8140 23910 8142 23962
rect 7896 23908 7902 23910
rect 7958 23908 7982 23910
rect 8038 23908 8062 23910
rect 8118 23908 8142 23910
rect 8198 23908 8204 23910
rect 7896 23899 8204 23908
rect 1400 23724 1452 23730
rect 1400 23666 1452 23672
rect 1412 23497 1440 23666
rect 1584 23520 1636 23526
rect 1398 23488 1454 23497
rect 1584 23462 1636 23468
rect 1398 23423 1454 23432
rect 940 23112 992 23118
rect 940 23054 992 23060
rect 952 22681 980 23054
rect 1032 23044 1084 23050
rect 1032 22986 1084 22992
rect 1044 22953 1072 22986
rect 1030 22944 1086 22953
rect 1030 22879 1086 22888
rect 938 22672 994 22681
rect 938 22607 994 22616
rect 1032 22636 1084 22642
rect 1032 22578 1084 22584
rect 940 22568 992 22574
rect 940 22510 992 22516
rect 952 22409 980 22510
rect 938 22400 994 22409
rect 938 22335 994 22344
rect 1044 22137 1072 22578
rect 1030 22128 1086 22137
rect 1030 22063 1086 22072
rect 940 22024 992 22030
rect 940 21966 992 21972
rect 952 21593 980 21966
rect 1032 21956 1084 21962
rect 1032 21898 1084 21904
rect 1044 21865 1072 21898
rect 1030 21856 1086 21865
rect 1030 21791 1086 21800
rect 938 21584 994 21593
rect 938 21519 994 21528
rect 1032 21548 1084 21554
rect 1032 21490 1084 21496
rect 940 21480 992 21486
rect 940 21422 992 21428
rect 952 21321 980 21422
rect 938 21312 994 21321
rect 938 21247 994 21256
rect 1044 21049 1072 21490
rect 1030 21040 1086 21049
rect 1030 20975 1086 20984
rect 1400 20936 1452 20942
rect 1400 20878 1452 20884
rect 940 20868 992 20874
rect 940 20810 992 20816
rect 952 20777 980 20810
rect 938 20768 994 20777
rect 938 20703 994 20712
rect 1412 20641 1440 20878
rect 1398 20632 1454 20641
rect 1398 20567 1454 20576
rect 940 20460 992 20466
rect 940 20402 992 20408
rect 952 19961 980 20402
rect 1032 20392 1084 20398
rect 1032 20334 1084 20340
rect 1596 20346 1624 23462
rect 4423 23420 4731 23429
rect 4423 23418 4429 23420
rect 4485 23418 4509 23420
rect 4565 23418 4589 23420
rect 4645 23418 4669 23420
rect 4725 23418 4731 23420
rect 4485 23366 4487 23418
rect 4667 23366 4669 23418
rect 4423 23364 4429 23366
rect 4485 23364 4509 23366
rect 4565 23364 4589 23366
rect 4645 23364 4669 23366
rect 4725 23364 4731 23366
rect 4423 23355 4731 23364
rect 11369 23420 11677 23429
rect 11369 23418 11375 23420
rect 11431 23418 11455 23420
rect 11511 23418 11535 23420
rect 11591 23418 11615 23420
rect 11671 23418 11677 23420
rect 11431 23366 11433 23418
rect 11613 23366 11615 23418
rect 11369 23364 11375 23366
rect 11431 23364 11455 23366
rect 11511 23364 11535 23366
rect 11591 23364 11615 23366
rect 11671 23364 11677 23366
rect 11369 23355 11677 23364
rect 4252 23248 4304 23254
rect 4252 23190 4304 23196
rect 1860 22976 1912 22982
rect 1860 22918 1912 22924
rect 1044 20233 1072 20334
rect 1596 20318 1808 20346
rect 1584 20256 1636 20262
rect 1030 20224 1086 20233
rect 1584 20198 1636 20204
rect 1030 20159 1086 20168
rect 938 19952 994 19961
rect 938 19887 994 19896
rect 940 19848 992 19854
rect 940 19790 992 19796
rect 952 19417 980 19790
rect 1032 19780 1084 19786
rect 1032 19722 1084 19728
rect 1044 19689 1072 19722
rect 1030 19680 1086 19689
rect 1030 19615 1086 19624
rect 938 19408 994 19417
rect 938 19343 994 19352
rect 1400 19372 1452 19378
rect 1400 19314 1452 19320
rect 1412 19009 1440 19314
rect 1398 19000 1454 19009
rect 1398 18935 1454 18944
rect 940 18760 992 18766
rect 940 18702 992 18708
rect 952 18329 980 18702
rect 1032 18692 1084 18698
rect 1032 18634 1084 18640
rect 1044 18601 1072 18634
rect 1030 18592 1086 18601
rect 1030 18527 1086 18536
rect 938 18320 994 18329
rect 938 18255 994 18264
rect 1400 18284 1452 18290
rect 1400 18226 1452 18232
rect 940 18216 992 18222
rect 940 18158 992 18164
rect 952 18057 980 18158
rect 938 18048 994 18057
rect 938 17983 994 17992
rect 1412 17921 1440 18226
rect 1398 17912 1454 17921
rect 1398 17847 1454 17856
rect 1032 17672 1084 17678
rect 1032 17614 1084 17620
rect 940 17604 992 17610
rect 940 17546 992 17552
rect 952 17513 980 17546
rect 938 17504 994 17513
rect 938 17439 994 17448
rect 1044 17241 1072 17614
rect 1030 17232 1086 17241
rect 940 17196 992 17202
rect 1030 17167 1086 17176
rect 940 17138 992 17144
rect 952 16969 980 17138
rect 1032 17128 1084 17134
rect 1032 17070 1084 17076
rect 938 16960 994 16969
rect 938 16895 994 16904
rect 1044 16697 1072 17070
rect 1308 17060 1360 17066
rect 1308 17002 1360 17008
rect 1030 16688 1086 16697
rect 1030 16623 1086 16632
rect 940 16584 992 16590
rect 1320 16574 1348 17002
rect 940 16526 992 16532
rect 1228 16546 1348 16574
rect 664 16448 716 16454
rect 952 16425 980 16526
rect 1032 16516 1084 16522
rect 1032 16458 1084 16464
rect 664 16390 716 16396
rect 938 16416 994 16425
rect 388 16244 440 16250
rect 388 16186 440 16192
rect 296 10260 348 10266
rect 296 10202 348 10208
rect 308 6798 336 10202
rect 296 6792 348 6798
rect 296 6734 348 6740
rect 400 5234 428 16186
rect 480 15360 532 15366
rect 480 15302 532 15308
rect 492 8022 520 15302
rect 676 10266 704 16390
rect 938 16351 994 16360
rect 1044 16153 1072 16458
rect 1030 16144 1086 16153
rect 940 16108 992 16114
rect 1030 16079 1086 16088
rect 940 16050 992 16056
rect 952 15881 980 16050
rect 1032 16040 1084 16046
rect 1032 15982 1084 15988
rect 938 15872 994 15881
rect 938 15807 994 15816
rect 940 15632 992 15638
rect 860 15580 940 15586
rect 1044 15609 1072 15982
rect 860 15574 992 15580
rect 1030 15600 1086 15609
rect 860 15558 980 15574
rect 860 12434 888 15558
rect 1030 15535 1086 15544
rect 940 15496 992 15502
rect 940 15438 992 15444
rect 952 15337 980 15438
rect 938 15328 994 15337
rect 938 15263 994 15272
rect 940 15020 992 15026
rect 940 14962 992 14968
rect 952 14521 980 14962
rect 938 14512 994 14521
rect 938 14447 994 14456
rect 940 14408 992 14414
rect 940 14350 992 14356
rect 952 14249 980 14350
rect 1032 14340 1084 14346
rect 1032 14282 1084 14288
rect 938 14240 994 14249
rect 938 14175 994 14184
rect 1044 13977 1072 14282
rect 1030 13968 1086 13977
rect 1030 13903 1086 13912
rect 940 13320 992 13326
rect 940 13262 992 13268
rect 952 13161 980 13262
rect 1032 13252 1084 13258
rect 1032 13194 1084 13200
rect 938 13152 994 13161
rect 938 13087 994 13096
rect 1044 12889 1072 13194
rect 1030 12880 1086 12889
rect 940 12844 992 12850
rect 1030 12815 1086 12824
rect 940 12786 992 12792
rect 952 12617 980 12786
rect 938 12608 994 12617
rect 938 12543 994 12552
rect 860 12406 1164 12434
rect 940 12232 992 12238
rect 940 12174 992 12180
rect 952 12073 980 12174
rect 1032 12164 1084 12170
rect 1032 12106 1084 12112
rect 938 12064 994 12073
rect 938 11999 994 12008
rect 1044 11801 1072 12106
rect 1030 11792 1086 11801
rect 940 11756 992 11762
rect 1030 11727 1086 11736
rect 940 11698 992 11704
rect 952 11529 980 11698
rect 1032 11688 1084 11694
rect 1032 11630 1084 11636
rect 938 11520 994 11529
rect 938 11455 994 11464
rect 1044 11257 1072 11630
rect 1030 11248 1086 11257
rect 1030 11183 1086 11192
rect 940 10668 992 10674
rect 940 10610 992 10616
rect 952 10441 980 10610
rect 1032 10600 1084 10606
rect 1032 10542 1084 10548
rect 938 10432 994 10441
rect 938 10367 994 10376
rect 664 10260 716 10266
rect 664 10202 716 10208
rect 1044 10169 1072 10542
rect 1030 10160 1086 10169
rect 1030 10095 1086 10104
rect 940 10056 992 10062
rect 940 9998 992 10004
rect 952 9897 980 9998
rect 938 9888 994 9897
rect 938 9823 994 9832
rect 940 9580 992 9586
rect 940 9522 992 9528
rect 952 9353 980 9522
rect 1032 9512 1084 9518
rect 1032 9454 1084 9460
rect 938 9344 994 9353
rect 938 9279 994 9288
rect 1044 9081 1072 9454
rect 1030 9072 1086 9081
rect 1030 9007 1086 9016
rect 940 8968 992 8974
rect 940 8910 992 8916
rect 848 8832 900 8838
rect 952 8809 980 8910
rect 1032 8900 1084 8906
rect 1032 8842 1084 8848
rect 848 8774 900 8780
rect 938 8800 994 8809
rect 756 8424 808 8430
rect 756 8366 808 8372
rect 480 8016 532 8022
rect 480 7958 532 7964
rect 768 7732 796 8366
rect 492 7704 796 7732
rect 388 5228 440 5234
rect 388 5170 440 5176
rect 492 800 520 7704
rect 756 7608 808 7614
rect 756 7550 808 7556
rect 664 7540 716 7546
rect 664 7482 716 7488
rect 676 5370 704 7482
rect 664 5364 716 5370
rect 664 5306 716 5312
rect 768 800 796 7550
rect 860 4214 888 8774
rect 938 8735 994 8744
rect 1044 8537 1072 8842
rect 1030 8528 1086 8537
rect 1030 8463 1086 8472
rect 1032 8424 1084 8430
rect 1030 8392 1032 8401
rect 1084 8392 1086 8401
rect 1030 8327 1086 8336
rect 1032 8288 1084 8294
rect 1032 8230 1084 8236
rect 940 7404 992 7410
rect 940 7346 992 7352
rect 952 7177 980 7346
rect 938 7168 994 7177
rect 938 7103 994 7112
rect 1044 4264 1072 8230
rect 1136 6866 1164 12406
rect 1228 7478 1256 16546
rect 1596 15502 1624 20198
rect 1676 19372 1728 19378
rect 1676 19314 1728 19320
rect 1688 19281 1716 19314
rect 1674 19272 1730 19281
rect 1674 19207 1730 19216
rect 1676 16448 1728 16454
rect 1676 16390 1728 16396
rect 1688 16250 1716 16390
rect 1676 16244 1728 16250
rect 1676 16186 1728 16192
rect 1676 15904 1728 15910
rect 1676 15846 1728 15852
rect 1584 15496 1636 15502
rect 1584 15438 1636 15444
rect 1688 15337 1716 15846
rect 1674 15328 1730 15337
rect 1674 15263 1730 15272
rect 1780 15094 1808 20318
rect 1872 19802 1900 22918
rect 2044 22500 2096 22506
rect 2044 22442 2096 22448
rect 1872 19774 1992 19802
rect 1860 19712 1912 19718
rect 1860 19654 1912 19660
rect 1872 17270 1900 19654
rect 1860 17264 1912 17270
rect 1860 17206 1912 17212
rect 1860 15496 1912 15502
rect 1860 15438 1912 15444
rect 1872 15201 1900 15438
rect 1858 15192 1914 15201
rect 1858 15127 1914 15136
rect 1768 15088 1820 15094
rect 1768 15030 1820 15036
rect 1584 14884 1636 14890
rect 1584 14826 1636 14832
rect 1596 14074 1624 14826
rect 1858 14376 1914 14385
rect 1858 14311 1914 14320
rect 1872 14278 1900 14311
rect 1964 14278 1992 19774
rect 1860 14272 1912 14278
rect 1860 14214 1912 14220
rect 1952 14272 2004 14278
rect 1952 14214 2004 14220
rect 1584 14068 1636 14074
rect 1584 14010 1636 14016
rect 1860 14068 1912 14074
rect 1860 14010 1912 14016
rect 1400 13932 1452 13938
rect 1400 13874 1452 13880
rect 1676 13932 1728 13938
rect 1676 13874 1728 13880
rect 1412 13705 1440 13874
rect 1688 13705 1716 13874
rect 1872 13841 1900 14010
rect 1858 13832 1914 13841
rect 2056 13802 2084 22442
rect 4068 21072 4120 21078
rect 4068 21014 4120 21020
rect 3608 19508 3660 19514
rect 3608 19450 3660 19456
rect 3332 18896 3384 18902
rect 3332 18838 3384 18844
rect 3240 15904 3292 15910
rect 3240 15846 3292 15852
rect 1858 13767 1914 13776
rect 2044 13796 2096 13802
rect 2044 13738 2096 13744
rect 1398 13696 1454 13705
rect 1398 13631 1454 13640
rect 1674 13696 1730 13705
rect 1674 13631 1730 13640
rect 1860 13456 1912 13462
rect 1858 13424 1860 13433
rect 1912 13424 1914 13433
rect 1858 13359 1914 13368
rect 1582 13288 1638 13297
rect 1582 13223 1638 13232
rect 1596 13190 1624 13223
rect 1584 13184 1636 13190
rect 1584 13126 1636 13132
rect 1676 12844 1728 12850
rect 1676 12786 1728 12792
rect 1688 12345 1716 12786
rect 1858 12744 1914 12753
rect 1858 12679 1860 12688
rect 1912 12679 1914 12688
rect 1860 12650 1912 12656
rect 1674 12336 1730 12345
rect 1674 12271 1730 12280
rect 1858 12200 1914 12209
rect 1858 12135 1914 12144
rect 1872 12102 1900 12135
rect 1860 12096 1912 12102
rect 1860 12038 1912 12044
rect 1860 11552 1912 11558
rect 1860 11494 1912 11500
rect 1872 11354 1900 11494
rect 1860 11348 1912 11354
rect 1860 11290 1912 11296
rect 1400 11144 1452 11150
rect 1400 11086 1452 11092
rect 1676 11144 1728 11150
rect 1676 11086 1728 11092
rect 1412 10985 1440 11086
rect 1688 10985 1716 11086
rect 1398 10976 1454 10985
rect 1398 10911 1454 10920
rect 1674 10976 1730 10985
rect 1674 10911 1730 10920
rect 1582 10568 1638 10577
rect 1582 10503 1584 10512
rect 1636 10503 1638 10512
rect 1584 10474 1636 10480
rect 1676 10056 1728 10062
rect 1676 9998 1728 10004
rect 1688 9625 1716 9998
rect 3148 9920 3200 9926
rect 3148 9862 3200 9868
rect 1674 9616 1730 9625
rect 1674 9551 1730 9560
rect 1768 9580 1820 9586
rect 1768 9522 1820 9528
rect 2044 9580 2096 9586
rect 2044 9522 2096 9528
rect 1584 9104 1636 9110
rect 1584 9046 1636 9052
rect 1308 9036 1360 9042
rect 1308 8978 1360 8984
rect 1216 7472 1268 7478
rect 1216 7414 1268 7420
rect 1320 7290 1348 8978
rect 1596 8809 1624 9046
rect 1582 8800 1638 8809
rect 1582 8735 1638 8744
rect 1584 8628 1636 8634
rect 1584 8570 1636 8576
rect 1492 8560 1544 8566
rect 1596 8537 1624 8570
rect 1492 8502 1544 8508
rect 1582 8528 1638 8537
rect 1400 8492 1452 8498
rect 1400 8434 1452 8440
rect 1412 8265 1440 8434
rect 1398 8256 1454 8265
rect 1398 8191 1454 8200
rect 1400 8084 1452 8090
rect 1400 8026 1452 8032
rect 1412 7886 1440 8026
rect 1400 7880 1452 7886
rect 1400 7822 1452 7828
rect 1320 7262 1440 7290
rect 1306 7168 1362 7177
rect 1228 7126 1306 7154
rect 1124 6860 1176 6866
rect 1124 6802 1176 6808
rect 1228 4690 1256 7126
rect 1306 7103 1362 7112
rect 1308 6724 1360 6730
rect 1308 6666 1360 6672
rect 1320 6361 1348 6666
rect 1306 6352 1362 6361
rect 1306 6287 1362 6296
rect 1412 6202 1440 7262
rect 1504 6905 1532 8502
rect 1582 8463 1638 8472
rect 1676 8492 1728 8498
rect 1676 8434 1728 8440
rect 1584 8288 1636 8294
rect 1688 8265 1716 8434
rect 1584 8230 1636 8236
rect 1674 8256 1730 8265
rect 1596 7886 1624 8230
rect 1674 8191 1730 8200
rect 1676 8084 1728 8090
rect 1676 8026 1728 8032
rect 1584 7880 1636 7886
rect 1584 7822 1636 7828
rect 1584 7744 1636 7750
rect 1584 7686 1636 7692
rect 1596 7274 1624 7686
rect 1584 7268 1636 7274
rect 1584 7210 1636 7216
rect 1688 7154 1716 8026
rect 1780 7721 1808 9522
rect 1860 8968 1912 8974
rect 1860 8910 1912 8916
rect 1766 7712 1822 7721
rect 1766 7647 1822 7656
rect 1768 7540 1820 7546
rect 1768 7482 1820 7488
rect 1596 7126 1716 7154
rect 1490 6896 1546 6905
rect 1490 6831 1546 6840
rect 1596 6746 1624 7126
rect 1780 6905 1808 7482
rect 1766 6896 1822 6905
rect 1766 6831 1822 6840
rect 1872 6746 1900 8910
rect 1952 8832 2004 8838
rect 1952 8774 2004 8780
rect 1964 8294 1992 8774
rect 2056 8566 2084 9522
rect 2136 9376 2188 9382
rect 2136 9318 2188 9324
rect 2412 9376 2464 9382
rect 2412 9318 2464 9324
rect 2148 8945 2176 9318
rect 2228 8968 2280 8974
rect 2134 8936 2190 8945
rect 2228 8910 2280 8916
rect 2134 8871 2190 8880
rect 2044 8560 2096 8566
rect 2044 8502 2096 8508
rect 2136 8492 2188 8498
rect 2136 8434 2188 8440
rect 1952 8288 2004 8294
rect 1952 8230 2004 8236
rect 2044 8288 2096 8294
rect 2044 8230 2096 8236
rect 2056 8106 2084 8230
rect 1964 8078 2084 8106
rect 1964 7818 1992 8078
rect 2044 7880 2096 7886
rect 2044 7822 2096 7828
rect 1952 7812 2004 7818
rect 1952 7754 2004 7760
rect 1952 7336 2004 7342
rect 1952 7278 2004 7284
rect 1320 6174 1440 6202
rect 1504 6718 1624 6746
rect 1688 6718 1900 6746
rect 1216 4684 1268 4690
rect 1216 4626 1268 4632
rect 1320 4622 1348 6174
rect 1308 4616 1360 4622
rect 1308 4558 1360 4564
rect 1504 4486 1532 6718
rect 1584 5228 1636 5234
rect 1584 5170 1636 5176
rect 1492 4480 1544 4486
rect 1492 4422 1544 4428
rect 1596 4282 1624 5170
rect 952 4236 1072 4264
rect 1584 4276 1636 4282
rect 848 4208 900 4214
rect 848 4150 900 4156
rect 952 4128 980 4236
rect 1584 4218 1636 4224
rect 1308 4208 1360 4214
rect 1308 4150 1360 4156
rect 952 4100 1072 4128
rect 1044 800 1072 4100
rect 1320 800 1348 4150
rect 1584 4140 1636 4146
rect 1584 4082 1636 4088
rect 1596 3466 1624 4082
rect 1584 3460 1636 3466
rect 1584 3402 1636 3408
rect 1688 2774 1716 6718
rect 1860 6656 1912 6662
rect 1860 6598 1912 6604
rect 1768 5704 1820 5710
rect 1768 5646 1820 5652
rect 1780 2854 1808 5646
rect 1872 2990 1900 6598
rect 1964 5545 1992 7278
rect 2056 6633 2084 7822
rect 2148 7750 2176 8434
rect 2136 7744 2188 7750
rect 2136 7686 2188 7692
rect 2042 6624 2098 6633
rect 2042 6559 2098 6568
rect 1950 5536 2006 5545
rect 1950 5471 2006 5480
rect 2148 5234 2176 7686
rect 2240 6458 2268 8910
rect 2320 8900 2372 8906
rect 2320 8842 2372 8848
rect 2332 8498 2360 8842
rect 2424 8673 2452 9318
rect 2504 8968 2556 8974
rect 2556 8928 2636 8956
rect 2504 8910 2556 8916
rect 2504 8832 2556 8838
rect 2504 8774 2556 8780
rect 2410 8664 2466 8673
rect 2410 8599 2466 8608
rect 2320 8492 2372 8498
rect 2320 8434 2372 8440
rect 2320 8356 2372 8362
rect 2320 8298 2372 8304
rect 2228 6452 2280 6458
rect 2228 6394 2280 6400
rect 2228 6248 2280 6254
rect 2228 6190 2280 6196
rect 2136 5228 2188 5234
rect 2136 5170 2188 5176
rect 1952 5160 2004 5166
rect 1952 5102 2004 5108
rect 1964 3194 1992 5102
rect 2240 4826 2268 6190
rect 2228 4820 2280 4826
rect 2228 4762 2280 4768
rect 2332 4146 2360 8298
rect 2412 7744 2464 7750
rect 2412 7686 2464 7692
rect 2424 5273 2452 7686
rect 2516 7410 2544 8774
rect 2504 7404 2556 7410
rect 2504 7346 2556 7352
rect 2502 7304 2558 7313
rect 2502 7239 2504 7248
rect 2556 7239 2558 7248
rect 2504 7210 2556 7216
rect 2504 6792 2556 6798
rect 2504 6734 2556 6740
rect 2410 5264 2466 5273
rect 2410 5199 2466 5208
rect 2516 5114 2544 6734
rect 2608 5778 2636 8928
rect 2780 8900 2832 8906
rect 2780 8842 2832 8848
rect 2792 8634 2820 8842
rect 3160 8838 3188 9862
rect 3148 8832 3200 8838
rect 3148 8774 3200 8780
rect 2780 8628 2832 8634
rect 2780 8570 2832 8576
rect 2872 8492 2924 8498
rect 2872 8434 2924 8440
rect 2964 8492 3016 8498
rect 2964 8434 3016 8440
rect 3148 8492 3200 8498
rect 3148 8434 3200 8440
rect 2688 7744 2740 7750
rect 2688 7686 2740 7692
rect 2778 7712 2834 7721
rect 2700 6914 2728 7686
rect 2778 7647 2834 7656
rect 2792 7449 2820 7647
rect 2778 7440 2834 7449
rect 2778 7375 2834 7384
rect 2700 6886 2820 6914
rect 2792 6610 2820 6886
rect 2884 6798 2912 8434
rect 2872 6792 2924 6798
rect 2872 6734 2924 6740
rect 2792 6582 2912 6610
rect 2780 6112 2832 6118
rect 2780 6054 2832 6060
rect 2596 5772 2648 5778
rect 2596 5714 2648 5720
rect 2424 5086 2544 5114
rect 2320 4140 2372 4146
rect 2320 4082 2372 4088
rect 2320 3936 2372 3942
rect 2320 3878 2372 3884
rect 2042 3496 2098 3505
rect 2042 3431 2098 3440
rect 2056 3398 2084 3431
rect 2044 3392 2096 3398
rect 2044 3334 2096 3340
rect 2332 3194 2360 3878
rect 1952 3188 2004 3194
rect 1952 3130 2004 3136
rect 2320 3188 2372 3194
rect 2320 3130 2372 3136
rect 1860 2984 1912 2990
rect 1860 2926 1912 2932
rect 1768 2848 1820 2854
rect 1768 2790 1820 2796
rect 1596 2746 1716 2774
rect 1596 800 1624 2746
rect 2320 2508 2372 2514
rect 2320 2450 2372 2456
rect 2136 2304 2188 2310
rect 2136 2246 2188 2252
rect 2148 1698 2176 2246
rect 2332 1970 2360 2450
rect 2320 1964 2372 1970
rect 2320 1906 2372 1912
rect 2424 1902 2452 5086
rect 2504 5024 2556 5030
rect 2504 4966 2556 4972
rect 2688 5024 2740 5030
rect 2688 4966 2740 4972
rect 2516 4282 2544 4966
rect 2504 4276 2556 4282
rect 2504 4218 2556 4224
rect 2700 3738 2728 4966
rect 2688 3732 2740 3738
rect 2688 3674 2740 3680
rect 2792 3534 2820 6054
rect 2596 3528 2648 3534
rect 2596 3470 2648 3476
rect 2780 3528 2832 3534
rect 2780 3470 2832 3476
rect 2608 2514 2636 3470
rect 2884 3466 2912 6582
rect 2976 5914 3004 8434
rect 3056 8356 3108 8362
rect 3056 8298 3108 8304
rect 3068 7177 3096 8298
rect 3160 7834 3188 8434
rect 3252 7954 3280 15846
rect 3344 11218 3372 18838
rect 3424 18148 3476 18154
rect 3424 18090 3476 18096
rect 3332 11212 3384 11218
rect 3332 11154 3384 11160
rect 3436 8906 3464 18090
rect 3516 17536 3568 17542
rect 3516 17478 3568 17484
rect 3528 9042 3556 17478
rect 3620 11830 3648 19450
rect 3976 19440 4028 19446
rect 3976 19382 4028 19388
rect 3792 18624 3844 18630
rect 3792 18566 3844 18572
rect 3700 17808 3752 17814
rect 3700 17750 3752 17756
rect 3608 11824 3660 11830
rect 3608 11766 3660 11772
rect 3516 9036 3568 9042
rect 3516 8978 3568 8984
rect 3608 8968 3660 8974
rect 3608 8910 3660 8916
rect 3424 8900 3476 8906
rect 3424 8842 3476 8848
rect 3516 8832 3568 8838
rect 3516 8774 3568 8780
rect 3332 8492 3384 8498
rect 3332 8434 3384 8440
rect 3240 7948 3292 7954
rect 3240 7890 3292 7896
rect 3160 7806 3280 7834
rect 3148 7744 3200 7750
rect 3148 7686 3200 7692
rect 3054 7168 3110 7177
rect 3054 7103 3110 7112
rect 2964 5908 3016 5914
rect 2964 5850 3016 5856
rect 2962 5536 3018 5545
rect 2962 5471 3018 5480
rect 2872 3460 2924 3466
rect 2872 3402 2924 3408
rect 2870 3360 2926 3369
rect 2870 3295 2926 3304
rect 2884 2990 2912 3295
rect 2872 2984 2924 2990
rect 2872 2926 2924 2932
rect 2596 2508 2648 2514
rect 2596 2450 2648 2456
rect 2872 2304 2924 2310
rect 2872 2246 2924 2252
rect 2412 1896 2464 1902
rect 2412 1838 2464 1844
rect 2136 1692 2188 1698
rect 2136 1634 2188 1640
rect 2884 1562 2912 2246
rect 2872 1556 2924 1562
rect 2872 1498 2924 1504
rect 2976 800 3004 5471
rect 3056 5364 3108 5370
rect 3056 5306 3108 5312
rect 3068 3942 3096 5306
rect 3160 4214 3188 7686
rect 3252 7392 3280 7806
rect 3344 7721 3372 8434
rect 3424 7880 3476 7886
rect 3424 7822 3476 7828
rect 3330 7712 3386 7721
rect 3330 7647 3386 7656
rect 3252 7364 3372 7392
rect 3240 6928 3292 6934
rect 3240 6870 3292 6876
rect 3148 4208 3200 4214
rect 3148 4150 3200 4156
rect 3056 3936 3108 3942
rect 3056 3878 3108 3884
rect 3068 3738 3096 3878
rect 3056 3732 3108 3738
rect 3056 3674 3108 3680
rect 3056 3460 3108 3466
rect 3056 3402 3108 3408
rect 3068 3058 3096 3402
rect 3056 3052 3108 3058
rect 3056 2994 3108 3000
rect 3056 2440 3108 2446
rect 3056 2382 3108 2388
rect 3068 2038 3096 2382
rect 3056 2032 3108 2038
rect 3056 1974 3108 1980
rect 3252 800 3280 6870
rect 3344 5846 3372 7364
rect 3436 5914 3464 7822
rect 3528 7750 3556 8774
rect 3516 7744 3568 7750
rect 3516 7686 3568 7692
rect 3620 7478 3648 8910
rect 3712 8498 3740 17750
rect 3804 11762 3832 18566
rect 3988 13394 4016 19382
rect 4080 18873 4108 21014
rect 4066 18864 4122 18873
rect 4066 18799 4122 18808
rect 4264 18222 4292 23190
rect 7896 22876 8204 22885
rect 7896 22874 7902 22876
rect 7958 22874 7982 22876
rect 8038 22874 8062 22876
rect 8118 22874 8142 22876
rect 8198 22874 8204 22876
rect 7958 22822 7960 22874
rect 8140 22822 8142 22874
rect 7896 22820 7902 22822
rect 7958 22820 7982 22822
rect 8038 22820 8062 22822
rect 8118 22820 8142 22822
rect 8198 22820 8204 22822
rect 7896 22811 8204 22820
rect 10232 22432 10284 22438
rect 10232 22374 10284 22380
rect 4423 22332 4731 22341
rect 4423 22330 4429 22332
rect 4485 22330 4509 22332
rect 4565 22330 4589 22332
rect 4645 22330 4669 22332
rect 4725 22330 4731 22332
rect 4485 22278 4487 22330
rect 4667 22278 4669 22330
rect 4423 22276 4429 22278
rect 4485 22276 4509 22278
rect 4565 22276 4589 22278
rect 4645 22276 4669 22278
rect 4725 22276 4731 22278
rect 4423 22267 4731 22276
rect 9220 21956 9272 21962
rect 9220 21898 9272 21904
rect 7896 21788 8204 21797
rect 7896 21786 7902 21788
rect 7958 21786 7982 21788
rect 8038 21786 8062 21788
rect 8118 21786 8142 21788
rect 8198 21786 8204 21788
rect 7958 21734 7960 21786
rect 8140 21734 8142 21786
rect 7896 21732 7902 21734
rect 7958 21732 7982 21734
rect 8038 21732 8062 21734
rect 8118 21732 8142 21734
rect 8198 21732 8204 21734
rect 7896 21723 8204 21732
rect 7472 21412 7524 21418
rect 7472 21354 7524 21360
rect 4423 21244 4731 21253
rect 4423 21242 4429 21244
rect 4485 21242 4509 21244
rect 4565 21242 4589 21244
rect 4645 21242 4669 21244
rect 4725 21242 4731 21244
rect 4485 21190 4487 21242
rect 4667 21190 4669 21242
rect 4423 21188 4429 21190
rect 4485 21188 4509 21190
rect 4565 21188 4589 21190
rect 4645 21188 4669 21190
rect 4725 21188 4731 21190
rect 4423 21179 4731 21188
rect 5540 20256 5592 20262
rect 5540 20198 5592 20204
rect 4423 20156 4731 20165
rect 4423 20154 4429 20156
rect 4485 20154 4509 20156
rect 4565 20154 4589 20156
rect 4645 20154 4669 20156
rect 4725 20154 4731 20156
rect 4485 20102 4487 20154
rect 4667 20102 4669 20154
rect 4423 20100 4429 20102
rect 4485 20100 4509 20102
rect 4565 20100 4589 20102
rect 4645 20100 4669 20102
rect 4725 20100 4731 20102
rect 4423 20091 4731 20100
rect 4423 19068 4731 19077
rect 4423 19066 4429 19068
rect 4485 19066 4509 19068
rect 4565 19066 4589 19068
rect 4645 19066 4669 19068
rect 4725 19066 4731 19068
rect 4485 19014 4487 19066
rect 4667 19014 4669 19066
rect 4423 19012 4429 19014
rect 4485 19012 4509 19014
rect 4565 19012 4589 19014
rect 4645 19012 4669 19014
rect 4725 19012 4731 19014
rect 4423 19003 4731 19012
rect 4252 18216 4304 18222
rect 4252 18158 4304 18164
rect 4160 18080 4212 18086
rect 4160 18022 4212 18028
rect 3976 13388 4028 13394
rect 3976 13330 4028 13336
rect 3792 11756 3844 11762
rect 3792 11698 3844 11704
rect 4172 10674 4200 18022
rect 4423 17980 4731 17989
rect 4423 17978 4429 17980
rect 4485 17978 4509 17980
rect 4565 17978 4589 17980
rect 4645 17978 4669 17980
rect 4725 17978 4731 17980
rect 4485 17926 4487 17978
rect 4667 17926 4669 17978
rect 4423 17924 4429 17926
rect 4485 17924 4509 17926
rect 4565 17924 4589 17926
rect 4645 17924 4669 17926
rect 4725 17924 4731 17926
rect 4423 17915 4731 17924
rect 5264 17332 5316 17338
rect 5264 17274 5316 17280
rect 4423 16892 4731 16901
rect 4423 16890 4429 16892
rect 4485 16890 4509 16892
rect 4565 16890 4589 16892
rect 4645 16890 4669 16892
rect 4725 16890 4731 16892
rect 4485 16838 4487 16890
rect 4667 16838 4669 16890
rect 4423 16836 4429 16838
rect 4485 16836 4509 16838
rect 4565 16836 4589 16838
rect 4645 16836 4669 16838
rect 4725 16836 4731 16838
rect 4423 16827 4731 16836
rect 4423 15804 4731 15813
rect 4423 15802 4429 15804
rect 4485 15802 4509 15804
rect 4565 15802 4589 15804
rect 4645 15802 4669 15804
rect 4725 15802 4731 15804
rect 4485 15750 4487 15802
rect 4667 15750 4669 15802
rect 4423 15748 4429 15750
rect 4485 15748 4509 15750
rect 4565 15748 4589 15750
rect 4645 15748 4669 15750
rect 4725 15748 4731 15750
rect 4423 15739 4731 15748
rect 4423 14716 4731 14725
rect 4423 14714 4429 14716
rect 4485 14714 4509 14716
rect 4565 14714 4589 14716
rect 4645 14714 4669 14716
rect 4725 14714 4731 14716
rect 4485 14662 4487 14714
rect 4667 14662 4669 14714
rect 4423 14660 4429 14662
rect 4485 14660 4509 14662
rect 4565 14660 4589 14662
rect 4645 14660 4669 14662
rect 4725 14660 4731 14662
rect 4423 14651 4731 14660
rect 4423 13628 4731 13637
rect 4423 13626 4429 13628
rect 4485 13626 4509 13628
rect 4565 13626 4589 13628
rect 4645 13626 4669 13628
rect 4725 13626 4731 13628
rect 4485 13574 4487 13626
rect 4667 13574 4669 13626
rect 4423 13572 4429 13574
rect 4485 13572 4509 13574
rect 4565 13572 4589 13574
rect 4645 13572 4669 13574
rect 4725 13572 4731 13574
rect 4423 13563 4731 13572
rect 4423 12540 4731 12549
rect 4423 12538 4429 12540
rect 4485 12538 4509 12540
rect 4565 12538 4589 12540
rect 4645 12538 4669 12540
rect 4725 12538 4731 12540
rect 4485 12486 4487 12538
rect 4667 12486 4669 12538
rect 4423 12484 4429 12486
rect 4485 12484 4509 12486
rect 4565 12484 4589 12486
rect 4645 12484 4669 12486
rect 4725 12484 4731 12486
rect 4423 12475 4731 12484
rect 5172 12096 5224 12102
rect 5172 12038 5224 12044
rect 5184 11801 5212 12038
rect 5170 11792 5226 11801
rect 5170 11727 5226 11736
rect 4423 11452 4731 11461
rect 4423 11450 4429 11452
rect 4485 11450 4509 11452
rect 4565 11450 4589 11452
rect 4645 11450 4669 11452
rect 4725 11450 4731 11452
rect 4485 11398 4487 11450
rect 4667 11398 4669 11450
rect 4423 11396 4429 11398
rect 4485 11396 4509 11398
rect 4565 11396 4589 11398
rect 4645 11396 4669 11398
rect 4725 11396 4731 11398
rect 4423 11387 4731 11396
rect 4896 11076 4948 11082
rect 4896 11018 4948 11024
rect 4160 10668 4212 10674
rect 4160 10610 4212 10616
rect 4344 10600 4396 10606
rect 4344 10542 4396 10548
rect 4160 10464 4212 10470
rect 4160 10406 4212 10412
rect 4172 9382 4200 10406
rect 3792 9376 3844 9382
rect 3792 9318 3844 9324
rect 4160 9376 4212 9382
rect 4160 9318 4212 9324
rect 3700 8492 3752 8498
rect 3700 8434 3752 8440
rect 3804 8344 3832 9318
rect 3712 8316 3832 8344
rect 3608 7472 3660 7478
rect 3608 7414 3660 7420
rect 3608 7336 3660 7342
rect 3608 7278 3660 7284
rect 3620 6934 3648 7278
rect 3712 7206 3740 8316
rect 4172 7954 4200 9318
rect 4252 8288 4304 8294
rect 4252 8230 4304 8236
rect 3884 7948 3936 7954
rect 3884 7890 3936 7896
rect 4160 7948 4212 7954
rect 4160 7890 4212 7896
rect 3896 7750 3924 7890
rect 3976 7880 4028 7886
rect 3976 7822 4028 7828
rect 3884 7744 3936 7750
rect 3884 7686 3936 7692
rect 3896 7426 3924 7686
rect 3988 7546 4016 7822
rect 4160 7744 4212 7750
rect 4160 7686 4212 7692
rect 3976 7540 4028 7546
rect 3976 7482 4028 7488
rect 3896 7398 4016 7426
rect 3700 7200 3752 7206
rect 3700 7142 3752 7148
rect 3608 6928 3660 6934
rect 3608 6870 3660 6876
rect 3516 6724 3568 6730
rect 3516 6666 3568 6672
rect 3424 5908 3476 5914
rect 3424 5850 3476 5856
rect 3332 5840 3384 5846
rect 3332 5782 3384 5788
rect 3332 5296 3384 5302
rect 3332 5238 3384 5244
rect 3344 3534 3372 5238
rect 3528 4758 3556 6666
rect 3608 6316 3660 6322
rect 3608 6258 3660 6264
rect 3516 4752 3568 4758
rect 3516 4694 3568 4700
rect 3332 3528 3384 3534
rect 3332 3470 3384 3476
rect 3620 2774 3648 6258
rect 3712 6254 3740 7142
rect 3792 6792 3844 6798
rect 3792 6734 3844 6740
rect 3700 6248 3752 6254
rect 3700 6190 3752 6196
rect 3700 5772 3752 5778
rect 3700 5714 3752 5720
rect 3712 5370 3740 5714
rect 3700 5364 3752 5370
rect 3700 5306 3752 5312
rect 3700 4072 3752 4078
rect 3700 4014 3752 4020
rect 3712 3058 3740 4014
rect 3700 3052 3752 3058
rect 3700 2994 3752 3000
rect 3804 2938 3832 6734
rect 3884 6656 3936 6662
rect 3884 6598 3936 6604
rect 3896 6458 3924 6598
rect 3884 6452 3936 6458
rect 3884 6394 3936 6400
rect 3884 6112 3936 6118
rect 3884 6054 3936 6060
rect 3896 5914 3924 6054
rect 3884 5908 3936 5914
rect 3884 5850 3936 5856
rect 3988 5794 4016 7398
rect 4068 7336 4120 7342
rect 4068 7278 4120 7284
rect 3896 5766 4016 5794
rect 3896 4706 3924 5766
rect 3976 5228 4028 5234
rect 3976 5170 4028 5176
rect 3988 4826 4016 5170
rect 4080 4826 4108 7278
rect 3976 4820 4028 4826
rect 3976 4762 4028 4768
rect 4068 4820 4120 4826
rect 4068 4762 4120 4768
rect 4066 4720 4122 4729
rect 3896 4690 4016 4706
rect 3896 4684 4028 4690
rect 3896 4678 3976 4684
rect 4066 4655 4122 4664
rect 3976 4626 4028 4632
rect 3884 4616 3936 4622
rect 3884 4558 3936 4564
rect 3896 3534 3924 4558
rect 3884 3528 3936 3534
rect 3884 3470 3936 3476
rect 3884 3392 3936 3398
rect 3988 3380 4016 4626
rect 4080 4622 4108 4655
rect 4068 4616 4120 4622
rect 4068 4558 4120 4564
rect 4172 4146 4200 7686
rect 4264 7546 4292 8230
rect 4252 7540 4304 7546
rect 4252 7482 4304 7488
rect 4356 6458 4384 10542
rect 4423 10364 4731 10373
rect 4423 10362 4429 10364
rect 4485 10362 4509 10364
rect 4565 10362 4589 10364
rect 4645 10362 4669 10364
rect 4725 10362 4731 10364
rect 4485 10310 4487 10362
rect 4667 10310 4669 10362
rect 4423 10308 4429 10310
rect 4485 10308 4509 10310
rect 4565 10308 4589 10310
rect 4645 10308 4669 10310
rect 4725 10308 4731 10310
rect 4423 10299 4731 10308
rect 4802 10024 4858 10033
rect 4724 9982 4802 10010
rect 4724 9654 4752 9982
rect 4802 9959 4858 9968
rect 4804 9920 4856 9926
rect 4804 9862 4856 9868
rect 4620 9648 4672 9654
rect 4618 9616 4620 9625
rect 4712 9648 4764 9654
rect 4672 9616 4674 9625
rect 4712 9590 4764 9596
rect 4618 9551 4674 9560
rect 4423 9276 4731 9285
rect 4423 9274 4429 9276
rect 4485 9274 4509 9276
rect 4565 9274 4589 9276
rect 4645 9274 4669 9276
rect 4725 9274 4731 9276
rect 4485 9222 4487 9274
rect 4667 9222 4669 9274
rect 4423 9220 4429 9222
rect 4485 9220 4509 9222
rect 4565 9220 4589 9222
rect 4645 9220 4669 9222
rect 4725 9220 4731 9222
rect 4423 9211 4731 9220
rect 4712 8832 4764 8838
rect 4816 8820 4844 9862
rect 4764 8792 4844 8820
rect 4712 8774 4764 8780
rect 4724 8362 4752 8774
rect 4712 8356 4764 8362
rect 4764 8316 4844 8344
rect 4712 8298 4764 8304
rect 4423 8188 4731 8197
rect 4423 8186 4429 8188
rect 4485 8186 4509 8188
rect 4565 8186 4589 8188
rect 4645 8186 4669 8188
rect 4725 8186 4731 8188
rect 4485 8134 4487 8186
rect 4667 8134 4669 8186
rect 4423 8132 4429 8134
rect 4485 8132 4509 8134
rect 4565 8132 4589 8134
rect 4645 8132 4669 8134
rect 4725 8132 4731 8134
rect 4423 8123 4731 8132
rect 4816 7834 4844 8316
rect 4724 7806 4844 7834
rect 4724 7342 4752 7806
rect 4804 7744 4856 7750
rect 4804 7686 4856 7692
rect 4712 7336 4764 7342
rect 4712 7278 4764 7284
rect 4423 7100 4731 7109
rect 4423 7098 4429 7100
rect 4485 7098 4509 7100
rect 4565 7098 4589 7100
rect 4645 7098 4669 7100
rect 4725 7098 4731 7100
rect 4485 7046 4487 7098
rect 4667 7046 4669 7098
rect 4423 7044 4429 7046
rect 4485 7044 4509 7046
rect 4565 7044 4589 7046
rect 4645 7044 4669 7046
rect 4725 7044 4731 7046
rect 4423 7035 4731 7044
rect 4344 6452 4396 6458
rect 4344 6394 4396 6400
rect 4252 6248 4304 6254
rect 4252 6190 4304 6196
rect 4264 5370 4292 6190
rect 4344 6180 4396 6186
rect 4344 6122 4396 6128
rect 4356 5658 4384 6122
rect 4423 6012 4731 6021
rect 4423 6010 4429 6012
rect 4485 6010 4509 6012
rect 4565 6010 4589 6012
rect 4645 6010 4669 6012
rect 4725 6010 4731 6012
rect 4485 5958 4487 6010
rect 4667 5958 4669 6010
rect 4423 5956 4429 5958
rect 4485 5956 4509 5958
rect 4565 5956 4589 5958
rect 4645 5956 4669 5958
rect 4725 5956 4731 5958
rect 4423 5947 4731 5956
rect 4356 5630 4568 5658
rect 4816 5642 4844 7686
rect 4908 6866 4936 11018
rect 5080 10736 5132 10742
rect 5080 10678 5132 10684
rect 5092 9625 5120 10678
rect 5078 9616 5134 9625
rect 5078 9551 5080 9560
rect 5132 9551 5134 9560
rect 5172 9580 5224 9586
rect 5080 9522 5132 9528
rect 5172 9522 5224 9528
rect 5184 9382 5212 9522
rect 5172 9376 5224 9382
rect 5172 9318 5224 9324
rect 5276 9194 5304 17274
rect 5552 17202 5580 20198
rect 5632 19984 5684 19990
rect 5632 19926 5684 19932
rect 5540 17196 5592 17202
rect 5540 17138 5592 17144
rect 5644 15026 5672 19926
rect 7380 17196 7432 17202
rect 7380 17138 7432 17144
rect 7196 17128 7248 17134
rect 7392 17082 7420 17138
rect 7196 17070 7248 17076
rect 6460 16992 6512 16998
rect 6460 16934 6512 16940
rect 6472 16658 6500 16934
rect 6460 16652 6512 16658
rect 6460 16594 6512 16600
rect 5724 16584 5776 16590
rect 5724 16526 5776 16532
rect 5632 15020 5684 15026
rect 5632 14962 5684 14968
rect 5736 14414 5764 16526
rect 6644 16516 6696 16522
rect 6644 16458 6696 16464
rect 6656 16250 6684 16458
rect 7208 16250 7236 17070
rect 7300 17054 7420 17082
rect 6644 16244 6696 16250
rect 6644 16186 6696 16192
rect 7196 16244 7248 16250
rect 7196 16186 7248 16192
rect 7012 16040 7064 16046
rect 7012 15982 7064 15988
rect 6920 14952 6972 14958
rect 6920 14894 6972 14900
rect 6276 14816 6328 14822
rect 6276 14758 6328 14764
rect 6288 14482 6316 14758
rect 6276 14476 6328 14482
rect 6276 14418 6328 14424
rect 5724 14408 5776 14414
rect 5724 14350 5776 14356
rect 5736 13326 5764 14350
rect 6932 14074 6960 14894
rect 6920 14068 6972 14074
rect 6920 14010 6972 14016
rect 6736 13796 6788 13802
rect 6736 13738 6788 13744
rect 6748 13530 6776 13738
rect 6736 13524 6788 13530
rect 6736 13466 6788 13472
rect 6736 13388 6788 13394
rect 6736 13330 6788 13336
rect 5632 13320 5684 13326
rect 5632 13262 5684 13268
rect 5724 13320 5776 13326
rect 5724 13262 5776 13268
rect 5644 12918 5672 13262
rect 5632 12912 5684 12918
rect 5632 12854 5684 12860
rect 5736 12374 5764 13262
rect 6000 13252 6052 13258
rect 6000 13194 6052 13200
rect 6012 12986 6040 13194
rect 6748 12986 6776 13330
rect 6828 13184 6880 13190
rect 6828 13126 6880 13132
rect 6840 12986 6868 13126
rect 6000 12980 6052 12986
rect 6000 12922 6052 12928
rect 6736 12980 6788 12986
rect 6736 12922 6788 12928
rect 6828 12980 6880 12986
rect 6828 12922 6880 12928
rect 5908 12912 5960 12918
rect 5908 12854 5960 12860
rect 5724 12368 5776 12374
rect 5724 12310 5776 12316
rect 5724 11280 5776 11286
rect 5724 11222 5776 11228
rect 5920 11234 5948 12854
rect 6000 12640 6052 12646
rect 6000 12582 6052 12588
rect 6012 11898 6040 12582
rect 7024 12434 7052 15982
rect 7300 15178 7328 17054
rect 7380 16992 7432 16998
rect 7380 16934 7432 16940
rect 7392 16250 7420 16934
rect 7380 16244 7432 16250
rect 7380 16186 7432 16192
rect 7484 16046 7512 21354
rect 8392 21344 8444 21350
rect 8392 21286 8444 21292
rect 7656 20800 7708 20806
rect 7656 20742 7708 20748
rect 7668 17202 7696 20742
rect 7896 20700 8204 20709
rect 7896 20698 7902 20700
rect 7958 20698 7982 20700
rect 8038 20698 8062 20700
rect 8118 20698 8142 20700
rect 8198 20698 8204 20700
rect 7958 20646 7960 20698
rect 8140 20646 8142 20698
rect 7896 20644 7902 20646
rect 7958 20644 7982 20646
rect 8038 20644 8062 20646
rect 8118 20644 8142 20646
rect 8198 20644 8204 20646
rect 7896 20635 8204 20644
rect 7896 19612 8204 19621
rect 7896 19610 7902 19612
rect 7958 19610 7982 19612
rect 8038 19610 8062 19612
rect 8118 19610 8142 19612
rect 8198 19610 8204 19612
rect 7958 19558 7960 19610
rect 8140 19558 8142 19610
rect 7896 19556 7902 19558
rect 7958 19556 7982 19558
rect 8038 19556 8062 19558
rect 8118 19556 8142 19558
rect 8198 19556 8204 19558
rect 7896 19547 8204 19556
rect 7896 18524 8204 18533
rect 7896 18522 7902 18524
rect 7958 18522 7982 18524
rect 8038 18522 8062 18524
rect 8118 18522 8142 18524
rect 8198 18522 8204 18524
rect 7958 18470 7960 18522
rect 8140 18470 8142 18522
rect 7896 18468 7902 18470
rect 7958 18468 7982 18470
rect 8038 18468 8062 18470
rect 8118 18468 8142 18470
rect 8198 18468 8204 18470
rect 7896 18459 8204 18468
rect 8300 18352 8352 18358
rect 8300 18294 8352 18300
rect 7896 17436 8204 17445
rect 7896 17434 7902 17436
rect 7958 17434 7982 17436
rect 8038 17434 8062 17436
rect 8118 17434 8142 17436
rect 8198 17434 8204 17436
rect 7958 17382 7960 17434
rect 8140 17382 8142 17434
rect 7896 17380 7902 17382
rect 7958 17380 7982 17382
rect 8038 17380 8062 17382
rect 8118 17380 8142 17382
rect 8198 17380 8204 17382
rect 7896 17371 8204 17380
rect 7656 17196 7708 17202
rect 7656 17138 7708 17144
rect 7564 17060 7616 17066
rect 7564 17002 7616 17008
rect 7380 16040 7432 16046
rect 7380 15982 7432 15988
rect 7472 16040 7524 16046
rect 7472 15982 7524 15988
rect 7392 15910 7420 15982
rect 7380 15904 7432 15910
rect 7380 15846 7432 15852
rect 7208 15150 7328 15178
rect 7104 14816 7156 14822
rect 7104 14758 7156 14764
rect 7116 14074 7144 14758
rect 7104 14068 7156 14074
rect 7104 14010 7156 14016
rect 7104 13864 7156 13870
rect 7104 13806 7156 13812
rect 7116 12782 7144 13806
rect 7104 12776 7156 12782
rect 7104 12718 7156 12724
rect 7024 12406 7144 12434
rect 7012 12300 7064 12306
rect 7012 12242 7064 12248
rect 6644 12232 6696 12238
rect 6644 12174 6696 12180
rect 6000 11892 6052 11898
rect 6000 11834 6052 11840
rect 6368 11756 6420 11762
rect 6368 11698 6420 11704
rect 5356 11008 5408 11014
rect 5356 10950 5408 10956
rect 5368 9994 5396 10950
rect 5736 10742 5764 11222
rect 5920 11206 6132 11234
rect 5908 11144 5960 11150
rect 5908 11086 5960 11092
rect 6000 11144 6052 11150
rect 6000 11086 6052 11092
rect 5920 10810 5948 11086
rect 5908 10804 5960 10810
rect 5908 10746 5960 10752
rect 5724 10736 5776 10742
rect 5724 10678 5776 10684
rect 6012 10130 6040 11086
rect 6000 10124 6052 10130
rect 6000 10066 6052 10072
rect 5722 10024 5778 10033
rect 5356 9988 5408 9994
rect 5722 9959 5724 9968
rect 5356 9930 5408 9936
rect 5776 9959 5778 9968
rect 5724 9930 5776 9936
rect 5908 9716 5960 9722
rect 5908 9658 5960 9664
rect 5920 9518 5948 9658
rect 5908 9512 5960 9518
rect 5908 9454 5960 9460
rect 5632 9444 5684 9450
rect 5632 9386 5684 9392
rect 5356 9376 5408 9382
rect 5356 9318 5408 9324
rect 5368 9217 5396 9318
rect 5092 9166 5304 9194
rect 5354 9208 5410 9217
rect 4988 8560 5040 8566
rect 4988 8502 5040 8508
rect 5000 7954 5028 8502
rect 5092 8090 5120 9166
rect 5644 9178 5672 9386
rect 5816 9376 5868 9382
rect 5816 9318 5868 9324
rect 5828 9178 5856 9318
rect 5354 9143 5410 9152
rect 5632 9172 5684 9178
rect 5632 9114 5684 9120
rect 5816 9172 5868 9178
rect 5816 9114 5868 9120
rect 5448 9104 5500 9110
rect 5500 9064 5580 9092
rect 5448 9046 5500 9052
rect 5172 8968 5224 8974
rect 5448 8968 5500 8974
rect 5224 8928 5304 8956
rect 5172 8910 5224 8916
rect 5172 8492 5224 8498
rect 5172 8434 5224 8440
rect 5080 8084 5132 8090
rect 5080 8026 5132 8032
rect 4988 7948 5040 7954
rect 4988 7890 5040 7896
rect 5080 7880 5132 7886
rect 5080 7822 5132 7828
rect 4988 7744 5040 7750
rect 4988 7686 5040 7692
rect 5000 7546 5028 7686
rect 4988 7540 5040 7546
rect 4988 7482 5040 7488
rect 4988 7200 5040 7206
rect 4988 7142 5040 7148
rect 4896 6860 4948 6866
rect 4896 6802 4948 6808
rect 4896 6656 4948 6662
rect 4896 6598 4948 6604
rect 4436 5568 4488 5574
rect 4436 5510 4488 5516
rect 4252 5364 4304 5370
rect 4252 5306 4304 5312
rect 4448 5250 4476 5510
rect 4264 5222 4476 5250
rect 4264 4570 4292 5222
rect 4540 5114 4568 5630
rect 4804 5636 4856 5642
rect 4804 5578 4856 5584
rect 4356 5086 4568 5114
rect 4356 4758 4384 5086
rect 4908 5030 4936 6598
rect 5000 5166 5028 7142
rect 5092 6866 5120 7822
rect 5080 6860 5132 6866
rect 5080 6802 5132 6808
rect 5080 6248 5132 6254
rect 5080 6190 5132 6196
rect 4988 5160 5040 5166
rect 4988 5102 5040 5108
rect 4896 5024 4948 5030
rect 4896 4966 4948 4972
rect 4423 4924 4731 4933
rect 4423 4922 4429 4924
rect 4485 4922 4509 4924
rect 4565 4922 4589 4924
rect 4645 4922 4669 4924
rect 4725 4922 4731 4924
rect 4485 4870 4487 4922
rect 4667 4870 4669 4922
rect 4423 4868 4429 4870
rect 4485 4868 4509 4870
rect 4565 4868 4589 4870
rect 4645 4868 4669 4870
rect 4725 4868 4731 4870
rect 4423 4859 4731 4868
rect 4344 4752 4396 4758
rect 4344 4694 4396 4700
rect 4264 4542 4384 4570
rect 4160 4140 4212 4146
rect 4160 4082 4212 4088
rect 4252 3936 4304 3942
rect 4252 3878 4304 3884
rect 4068 3596 4120 3602
rect 4068 3538 4120 3544
rect 3936 3352 4016 3380
rect 3884 3334 3936 3340
rect 3896 3058 3924 3334
rect 4080 3058 4108 3538
rect 3884 3052 3936 3058
rect 3884 2994 3936 3000
rect 4068 3052 4120 3058
rect 4068 2994 4120 3000
rect 3804 2910 4108 2938
rect 3792 2848 3844 2854
rect 3792 2790 3844 2796
rect 3528 2746 3648 2774
rect 3528 800 3556 2746
rect 3608 2304 3660 2310
rect 3608 2246 3660 2252
rect 3620 1834 3648 2246
rect 3608 1828 3660 1834
rect 3608 1770 3660 1776
rect 3804 800 3832 2790
rect 4080 800 4108 2910
rect 4264 2854 4292 3878
rect 4252 2848 4304 2854
rect 4252 2790 4304 2796
rect 4356 800 4384 4542
rect 4802 4040 4858 4049
rect 4802 3975 4858 3984
rect 4423 3836 4731 3845
rect 4423 3834 4429 3836
rect 4485 3834 4509 3836
rect 4565 3834 4589 3836
rect 4645 3834 4669 3836
rect 4725 3834 4731 3836
rect 4485 3782 4487 3834
rect 4667 3782 4669 3834
rect 4423 3780 4429 3782
rect 4485 3780 4509 3782
rect 4565 3780 4589 3782
rect 4645 3780 4669 3782
rect 4725 3780 4731 3782
rect 4423 3771 4731 3780
rect 4528 3732 4580 3738
rect 4528 3674 4580 3680
rect 4540 3466 4568 3674
rect 4816 3534 4844 3975
rect 5000 3942 5028 5102
rect 4988 3936 5040 3942
rect 4988 3878 5040 3884
rect 5000 3738 5028 3878
rect 4988 3732 5040 3738
rect 4988 3674 5040 3680
rect 4804 3528 4856 3534
rect 5092 3505 5120 6190
rect 5184 4826 5212 8434
rect 5172 4820 5224 4826
rect 5172 4762 5224 4768
rect 5276 4622 5304 8928
rect 5368 8916 5448 8922
rect 5368 8910 5500 8916
rect 5552 8922 5580 9064
rect 5368 8894 5488 8910
rect 5552 8894 5764 8922
rect 6012 8906 6040 10066
rect 5368 6914 5396 8894
rect 5540 8832 5592 8838
rect 5540 8774 5592 8780
rect 5552 8566 5580 8774
rect 5540 8560 5592 8566
rect 5540 8502 5592 8508
rect 5632 8084 5684 8090
rect 5632 8026 5684 8032
rect 5540 7812 5592 7818
rect 5540 7754 5592 7760
rect 5368 6886 5488 6914
rect 5356 6724 5408 6730
rect 5356 6666 5408 6672
rect 5368 6458 5396 6666
rect 5356 6452 5408 6458
rect 5356 6394 5408 6400
rect 5460 5370 5488 6886
rect 5448 5364 5500 5370
rect 5448 5306 5500 5312
rect 5356 5160 5408 5166
rect 5356 5102 5408 5108
rect 5368 4690 5396 5102
rect 5552 4826 5580 7754
rect 5540 4820 5592 4826
rect 5540 4762 5592 4768
rect 5356 4684 5408 4690
rect 5356 4626 5408 4632
rect 5264 4616 5316 4622
rect 5264 4558 5316 4564
rect 5644 4146 5672 8026
rect 5736 7750 5764 8894
rect 6000 8900 6052 8906
rect 6000 8842 6052 8848
rect 5908 8628 5960 8634
rect 5908 8570 5960 8576
rect 5920 8090 5948 8570
rect 5908 8084 5960 8090
rect 5908 8026 5960 8032
rect 5724 7744 5776 7750
rect 5724 7686 5776 7692
rect 5736 7478 5764 7686
rect 5724 7472 5776 7478
rect 5724 7414 5776 7420
rect 5908 7268 5960 7274
rect 5908 7210 5960 7216
rect 5920 6322 5948 7210
rect 5908 6316 5960 6322
rect 5908 6258 5960 6264
rect 5908 6112 5960 6118
rect 5908 6054 5960 6060
rect 5920 5624 5948 6054
rect 6012 5778 6040 8842
rect 6104 8514 6132 11206
rect 6184 10804 6236 10810
rect 6184 10746 6236 10752
rect 6196 10606 6224 10746
rect 6184 10600 6236 10606
rect 6184 10542 6236 10548
rect 6184 9580 6236 9586
rect 6184 9522 6236 9528
rect 6196 8634 6224 9522
rect 6184 8628 6236 8634
rect 6184 8570 6236 8576
rect 6104 8486 6224 8514
rect 6092 8424 6144 8430
rect 6092 8366 6144 8372
rect 6104 7342 6132 8366
rect 6196 7546 6224 8486
rect 6276 8424 6328 8430
rect 6276 8366 6328 8372
rect 6184 7540 6236 7546
rect 6184 7482 6236 7488
rect 6288 7410 6316 8366
rect 6276 7404 6328 7410
rect 6276 7346 6328 7352
rect 6092 7336 6144 7342
rect 6092 7278 6144 7284
rect 6274 6760 6330 6769
rect 6274 6695 6330 6704
rect 6000 5772 6052 5778
rect 6000 5714 6052 5720
rect 6000 5636 6052 5642
rect 5920 5596 6000 5624
rect 6000 5578 6052 5584
rect 6092 5636 6144 5642
rect 6092 5578 6144 5584
rect 5816 5568 5868 5574
rect 5816 5510 5868 5516
rect 5828 4690 5856 5510
rect 6012 5302 6040 5578
rect 6104 5370 6132 5578
rect 6092 5364 6144 5370
rect 6092 5306 6144 5312
rect 6000 5296 6052 5302
rect 6000 5238 6052 5244
rect 6090 5264 6146 5273
rect 6090 5199 6146 5208
rect 6104 5166 6132 5199
rect 6092 5160 6144 5166
rect 6092 5102 6144 5108
rect 5816 4684 5868 4690
rect 5816 4626 5868 4632
rect 5908 4616 5960 4622
rect 5908 4558 5960 4564
rect 5920 4264 5948 4558
rect 5828 4236 5948 4264
rect 5828 4146 5856 4236
rect 6184 4208 6236 4214
rect 6184 4150 6236 4156
rect 5448 4140 5500 4146
rect 5448 4082 5500 4088
rect 5632 4140 5684 4146
rect 5632 4082 5684 4088
rect 5816 4140 5868 4146
rect 5816 4082 5868 4088
rect 5172 4004 5224 4010
rect 5172 3946 5224 3952
rect 4804 3470 4856 3476
rect 5078 3496 5134 3505
rect 4528 3460 4580 3466
rect 5078 3431 5134 3440
rect 4528 3402 4580 3408
rect 4540 3369 4568 3402
rect 4896 3392 4948 3398
rect 4526 3360 4582 3369
rect 4896 3334 4948 3340
rect 4526 3295 4582 3304
rect 4804 2848 4856 2854
rect 4804 2790 4856 2796
rect 4423 2748 4731 2757
rect 4423 2746 4429 2748
rect 4485 2746 4509 2748
rect 4565 2746 4589 2748
rect 4645 2746 4669 2748
rect 4725 2746 4731 2748
rect 4485 2694 4487 2746
rect 4667 2694 4669 2746
rect 4423 2692 4429 2694
rect 4485 2692 4509 2694
rect 4565 2692 4589 2694
rect 4645 2692 4669 2694
rect 4725 2692 4731 2694
rect 4423 2683 4731 2692
rect 4816 1306 4844 2790
rect 4632 1278 4844 1306
rect 4632 800 4660 1278
rect 4908 800 4936 3334
rect 5184 800 5212 3946
rect 5460 3194 5488 4082
rect 5908 3936 5960 3942
rect 5908 3878 5960 3884
rect 5920 3602 5948 3878
rect 5908 3596 5960 3602
rect 5908 3538 5960 3544
rect 5448 3188 5500 3194
rect 5448 3130 5500 3136
rect 6196 3126 6224 4150
rect 6184 3120 6236 3126
rect 6184 3062 6236 3068
rect 6288 2650 6316 6695
rect 6380 6458 6408 11698
rect 6656 11082 6684 12174
rect 6828 12096 6880 12102
rect 6828 12038 6880 12044
rect 6840 11898 6868 12038
rect 6828 11892 6880 11898
rect 6828 11834 6880 11840
rect 6920 11824 6972 11830
rect 6920 11766 6972 11772
rect 6644 11076 6696 11082
rect 6644 11018 6696 11024
rect 6552 10668 6604 10674
rect 6552 10610 6604 10616
rect 6644 10668 6696 10674
rect 6644 10610 6696 10616
rect 6828 10668 6880 10674
rect 6828 10610 6880 10616
rect 6564 10538 6592 10610
rect 6460 10532 6512 10538
rect 6460 10474 6512 10480
rect 6552 10532 6604 10538
rect 6552 10474 6604 10480
rect 6472 10266 6500 10474
rect 6460 10260 6512 10266
rect 6460 10202 6512 10208
rect 6656 10062 6684 10610
rect 6644 10056 6696 10062
rect 6644 9998 6696 10004
rect 6840 9722 6868 10610
rect 6828 9716 6880 9722
rect 6828 9658 6880 9664
rect 6460 9580 6512 9586
rect 6460 9522 6512 9528
rect 6552 9580 6604 9586
rect 6552 9522 6604 9528
rect 6472 9178 6500 9522
rect 6460 9172 6512 9178
rect 6460 9114 6512 9120
rect 6564 8401 6592 9522
rect 6642 8800 6698 8809
rect 6698 8758 6776 8786
rect 6642 8735 6698 8744
rect 6550 8392 6606 8401
rect 6550 8327 6606 8336
rect 6460 8016 6512 8022
rect 6460 7958 6512 7964
rect 6472 7410 6500 7958
rect 6748 7886 6776 8758
rect 6736 7880 6788 7886
rect 6736 7822 6788 7828
rect 6932 7546 6960 11766
rect 7024 10810 7052 12242
rect 7012 10804 7064 10810
rect 7012 10746 7064 10752
rect 7024 10130 7052 10746
rect 7012 10124 7064 10130
rect 7012 10066 7064 10072
rect 7116 9466 7144 12406
rect 7208 9654 7236 15150
rect 7288 15020 7340 15026
rect 7288 14962 7340 14968
rect 7196 9648 7248 9654
rect 7196 9590 7248 9596
rect 7116 9438 7236 9466
rect 7104 9376 7156 9382
rect 7104 9318 7156 9324
rect 7012 7812 7064 7818
rect 7012 7754 7064 7760
rect 7024 7546 7052 7754
rect 6920 7540 6972 7546
rect 6920 7482 6972 7488
rect 7012 7540 7064 7546
rect 7012 7482 7064 7488
rect 6828 7472 6880 7478
rect 6828 7414 6880 7420
rect 6460 7404 6512 7410
rect 6460 7346 6512 7352
rect 6552 7268 6604 7274
rect 6552 7210 6604 7216
rect 6460 6792 6512 6798
rect 6460 6734 6512 6740
rect 6368 6452 6420 6458
rect 6368 6394 6420 6400
rect 6472 5370 6500 6734
rect 6460 5364 6512 5370
rect 6460 5306 6512 5312
rect 6564 5234 6592 7210
rect 6840 6866 6868 7414
rect 7012 7336 7064 7342
rect 7012 7278 7064 7284
rect 7024 7177 7052 7278
rect 7010 7168 7066 7177
rect 7010 7103 7066 7112
rect 6918 6896 6974 6905
rect 6828 6860 6880 6866
rect 6974 6854 7052 6882
rect 6918 6831 6974 6840
rect 6828 6802 6880 6808
rect 6736 6724 6788 6730
rect 6736 6666 6788 6672
rect 6644 6248 6696 6254
rect 6644 6190 6696 6196
rect 6656 5846 6684 6190
rect 6748 5914 6776 6666
rect 6736 5908 6788 5914
rect 6736 5850 6788 5856
rect 6644 5840 6696 5846
rect 6644 5782 6696 5788
rect 6552 5228 6604 5234
rect 6552 5170 6604 5176
rect 6550 5128 6606 5137
rect 6550 5063 6606 5072
rect 6564 3058 6592 5063
rect 6644 5024 6696 5030
rect 6644 4966 6696 4972
rect 6656 4690 6684 4966
rect 6644 4684 6696 4690
rect 6644 4626 6696 4632
rect 6748 4622 6776 5850
rect 7024 4672 7052 6854
rect 7116 5642 7144 9318
rect 7208 8090 7236 9438
rect 7300 8634 7328 14962
rect 7392 13870 7420 15846
rect 7472 14340 7524 14346
rect 7472 14282 7524 14288
rect 7484 14006 7512 14282
rect 7472 14000 7524 14006
rect 7472 13942 7524 13948
rect 7380 13864 7432 13870
rect 7380 13806 7432 13812
rect 7380 13252 7432 13258
rect 7380 13194 7432 13200
rect 7392 12986 7420 13194
rect 7380 12980 7432 12986
rect 7380 12922 7432 12928
rect 7472 12980 7524 12986
rect 7472 12922 7524 12928
rect 7380 12776 7432 12782
rect 7380 12718 7432 12724
rect 7392 12306 7420 12718
rect 7380 12300 7432 12306
rect 7380 12242 7432 12248
rect 7484 11914 7512 12922
rect 7392 11886 7512 11914
rect 7392 11830 7420 11886
rect 7380 11824 7432 11830
rect 7380 11766 7432 11772
rect 7380 11280 7432 11286
rect 7380 11222 7432 11228
rect 7392 11014 7420 11222
rect 7472 11144 7524 11150
rect 7472 11086 7524 11092
rect 7380 11008 7432 11014
rect 7380 10950 7432 10956
rect 7484 10810 7512 11086
rect 7472 10804 7524 10810
rect 7472 10746 7524 10752
rect 7380 10260 7432 10266
rect 7380 10202 7432 10208
rect 7392 9654 7420 10202
rect 7380 9648 7432 9654
rect 7380 9590 7432 9596
rect 7576 9178 7604 17002
rect 7748 16992 7800 16998
rect 7748 16934 7800 16940
rect 7760 15978 7788 16934
rect 8312 16658 8340 18294
rect 8404 16658 8432 21286
rect 9232 18290 9260 21898
rect 9680 21888 9732 21894
rect 9680 21830 9732 21836
rect 9692 18290 9720 21830
rect 9220 18284 9272 18290
rect 9220 18226 9272 18232
rect 9404 18284 9456 18290
rect 9404 18226 9456 18232
rect 9680 18284 9732 18290
rect 9680 18226 9732 18232
rect 9864 18284 9916 18290
rect 9864 18226 9916 18232
rect 8760 17536 8812 17542
rect 8760 17478 8812 17484
rect 9312 17536 9364 17542
rect 9312 17478 9364 17484
rect 8772 17134 8800 17478
rect 8852 17332 8904 17338
rect 8852 17274 8904 17280
rect 8760 17128 8812 17134
rect 8760 17070 8812 17076
rect 8300 16652 8352 16658
rect 8300 16594 8352 16600
rect 8392 16652 8444 16658
rect 8392 16594 8444 16600
rect 8312 16538 8340 16594
rect 8576 16584 8628 16590
rect 8312 16510 8432 16538
rect 8576 16526 8628 16532
rect 8300 16448 8352 16454
rect 8300 16390 8352 16396
rect 7896 16348 8204 16357
rect 7896 16346 7902 16348
rect 7958 16346 7982 16348
rect 8038 16346 8062 16348
rect 8118 16346 8142 16348
rect 8198 16346 8204 16348
rect 7958 16294 7960 16346
rect 8140 16294 8142 16346
rect 7896 16292 7902 16294
rect 7958 16292 7982 16294
rect 8038 16292 8062 16294
rect 8118 16292 8142 16294
rect 8198 16292 8204 16294
rect 7896 16283 8204 16292
rect 8312 16114 8340 16390
rect 8404 16250 8432 16510
rect 8392 16244 8444 16250
rect 8392 16186 8444 16192
rect 8300 16108 8352 16114
rect 8300 16050 8352 16056
rect 7656 15972 7708 15978
rect 7656 15914 7708 15920
rect 7748 15972 7800 15978
rect 7748 15914 7800 15920
rect 7668 15026 7696 15914
rect 8208 15904 8260 15910
rect 8208 15846 8260 15852
rect 8220 15706 8248 15846
rect 8208 15700 8260 15706
rect 8208 15642 8260 15648
rect 8404 15570 8432 16186
rect 8392 15564 8444 15570
rect 8392 15506 8444 15512
rect 7748 15428 7800 15434
rect 7748 15370 7800 15376
rect 7656 15020 7708 15026
rect 7656 14962 7708 14968
rect 7656 14816 7708 14822
rect 7656 14758 7708 14764
rect 7668 14414 7696 14758
rect 7656 14408 7708 14414
rect 7656 14350 7708 14356
rect 7656 13456 7708 13462
rect 7656 13398 7708 13404
rect 7668 12986 7696 13398
rect 7656 12980 7708 12986
rect 7656 12922 7708 12928
rect 7760 12434 7788 15370
rect 7896 15260 8204 15269
rect 7896 15258 7902 15260
rect 7958 15258 7982 15260
rect 8038 15258 8062 15260
rect 8118 15258 8142 15260
rect 8198 15258 8204 15260
rect 7958 15206 7960 15258
rect 8140 15206 8142 15258
rect 7896 15204 7902 15206
rect 7958 15204 7982 15206
rect 8038 15204 8062 15206
rect 8118 15204 8142 15206
rect 8198 15204 8204 15206
rect 7896 15195 8204 15204
rect 8300 14612 8352 14618
rect 8300 14554 8352 14560
rect 7896 14172 8204 14181
rect 7896 14170 7902 14172
rect 7958 14170 7982 14172
rect 8038 14170 8062 14172
rect 8118 14170 8142 14172
rect 8198 14170 8204 14172
rect 7958 14118 7960 14170
rect 8140 14118 8142 14170
rect 7896 14116 7902 14118
rect 7958 14116 7982 14118
rect 8038 14116 8062 14118
rect 8118 14116 8142 14118
rect 8198 14116 8204 14118
rect 7896 14107 8204 14116
rect 8116 13728 8168 13734
rect 8116 13670 8168 13676
rect 8128 13462 8156 13670
rect 8116 13456 8168 13462
rect 8116 13398 8168 13404
rect 8312 13394 8340 14554
rect 8404 13938 8432 15506
rect 8392 13932 8444 13938
rect 8392 13874 8444 13880
rect 8390 13696 8446 13705
rect 8390 13631 8446 13640
rect 8300 13388 8352 13394
rect 8300 13330 8352 13336
rect 8312 13138 8340 13330
rect 8404 13326 8432 13631
rect 8392 13320 8444 13326
rect 8392 13262 8444 13268
rect 8312 13110 8524 13138
rect 7896 13084 8204 13093
rect 7896 13082 7902 13084
rect 7958 13082 7982 13084
rect 8038 13082 8062 13084
rect 8118 13082 8142 13084
rect 8198 13082 8204 13084
rect 7958 13030 7960 13082
rect 8140 13030 8142 13082
rect 7896 13028 7902 13030
rect 7958 13028 7982 13030
rect 8038 13028 8062 13030
rect 8118 13028 8142 13030
rect 8198 13028 8204 13030
rect 7896 13019 8204 13028
rect 7840 12980 7892 12986
rect 7840 12922 7892 12928
rect 7668 12406 7788 12434
rect 7668 11218 7696 12406
rect 7852 12374 7880 12922
rect 8022 12880 8078 12889
rect 8078 12824 8432 12832
rect 8022 12815 8024 12824
rect 8076 12804 8432 12824
rect 8024 12786 8076 12792
rect 7932 12708 7984 12714
rect 7932 12650 7984 12656
rect 7944 12481 7972 12650
rect 7930 12472 7986 12481
rect 7930 12407 7986 12416
rect 7840 12368 7892 12374
rect 7840 12310 7892 12316
rect 7748 12164 7800 12170
rect 7748 12106 7800 12112
rect 7656 11212 7708 11218
rect 7656 11154 7708 11160
rect 7760 10674 7788 12106
rect 7932 12096 7984 12102
rect 7984 12056 8340 12084
rect 7932 12038 7984 12044
rect 7896 11996 8204 12005
rect 7896 11994 7902 11996
rect 7958 11994 7982 11996
rect 8038 11994 8062 11996
rect 8118 11994 8142 11996
rect 8198 11994 8204 11996
rect 7958 11942 7960 11994
rect 8140 11942 8142 11994
rect 7896 11940 7902 11942
rect 7958 11940 7982 11942
rect 8038 11940 8062 11942
rect 8118 11940 8142 11942
rect 8198 11940 8204 11942
rect 7896 11931 8204 11940
rect 8024 11892 8076 11898
rect 8024 11834 8076 11840
rect 7930 11792 7986 11801
rect 7930 11727 7986 11736
rect 7944 11694 7972 11727
rect 7932 11688 7984 11694
rect 7932 11630 7984 11636
rect 8036 11082 8064 11834
rect 8312 11778 8340 12056
rect 8220 11750 8340 11778
rect 8220 11694 8248 11750
rect 8208 11688 8260 11694
rect 8208 11630 8260 11636
rect 8404 11234 8432 12804
rect 8312 11206 8432 11234
rect 8024 11076 8076 11082
rect 8024 11018 8076 11024
rect 7896 10908 8204 10917
rect 7896 10906 7902 10908
rect 7958 10906 7982 10908
rect 8038 10906 8062 10908
rect 8118 10906 8142 10908
rect 8198 10906 8204 10908
rect 7958 10854 7960 10906
rect 8140 10854 8142 10906
rect 7896 10852 7902 10854
rect 7958 10852 7982 10854
rect 8038 10852 8062 10854
rect 8118 10852 8142 10854
rect 8198 10852 8204 10854
rect 7896 10843 8204 10852
rect 7748 10668 7800 10674
rect 7748 10610 7800 10616
rect 7760 9382 7788 10610
rect 8312 10606 8340 11206
rect 8392 11144 8444 11150
rect 8392 11086 8444 11092
rect 8300 10600 8352 10606
rect 8300 10542 8352 10548
rect 7896 9820 8204 9829
rect 7896 9818 7902 9820
rect 7958 9818 7982 9820
rect 8038 9818 8062 9820
rect 8118 9818 8142 9820
rect 8198 9818 8204 9820
rect 7958 9766 7960 9818
rect 8140 9766 8142 9818
rect 7896 9764 7902 9766
rect 7958 9764 7982 9766
rect 8038 9764 8062 9766
rect 8118 9764 8142 9766
rect 8198 9764 8204 9766
rect 7896 9755 8204 9764
rect 7840 9716 7892 9722
rect 7840 9658 7892 9664
rect 7748 9376 7800 9382
rect 7748 9318 7800 9324
rect 7472 9172 7524 9178
rect 7472 9114 7524 9120
rect 7564 9172 7616 9178
rect 7564 9114 7616 9120
rect 7288 8628 7340 8634
rect 7288 8570 7340 8576
rect 7380 8492 7432 8498
rect 7380 8434 7432 8440
rect 7196 8084 7248 8090
rect 7196 8026 7248 8032
rect 7288 7812 7340 7818
rect 7288 7754 7340 7760
rect 7196 6384 7248 6390
rect 7196 6326 7248 6332
rect 7104 5636 7156 5642
rect 7104 5578 7156 5584
rect 7104 4684 7156 4690
rect 7024 4644 7104 4672
rect 7104 4626 7156 4632
rect 6736 4616 6788 4622
rect 6736 4558 6788 4564
rect 7104 4548 7156 4554
rect 7104 4490 7156 4496
rect 6828 4004 6880 4010
rect 6828 3946 6880 3952
rect 6552 3052 6604 3058
rect 6552 2994 6604 3000
rect 6734 2952 6790 2961
rect 6734 2887 6736 2896
rect 6788 2887 6790 2896
rect 6736 2858 6788 2864
rect 6276 2644 6328 2650
rect 6276 2586 6328 2592
rect 6184 2508 6236 2514
rect 6184 2450 6236 2456
rect 5356 2440 5408 2446
rect 5356 2382 5408 2388
rect 5264 2304 5316 2310
rect 5264 2246 5316 2252
rect 5276 1306 5304 2246
rect 5368 2106 5396 2382
rect 5356 2100 5408 2106
rect 5356 2042 5408 2048
rect 6196 2038 6224 2450
rect 6276 2440 6328 2446
rect 6276 2382 6328 2388
rect 6000 2032 6052 2038
rect 6000 1974 6052 1980
rect 6184 2032 6236 2038
rect 6184 1974 6236 1980
rect 5724 1964 5776 1970
rect 5724 1906 5776 1912
rect 5276 1278 5488 1306
rect 5460 800 5488 1278
rect 5736 800 5764 1906
rect 6012 800 6040 1974
rect 6288 800 6316 2382
rect 6552 2100 6604 2106
rect 6552 2042 6604 2048
rect 6564 800 6592 2042
rect 6840 800 6868 3946
rect 7116 3534 7144 4490
rect 7104 3528 7156 3534
rect 7104 3470 7156 3476
rect 7208 3466 7236 6326
rect 7196 3460 7248 3466
rect 7196 3402 7248 3408
rect 7300 2774 7328 7754
rect 7392 6458 7420 8434
rect 7380 6452 7432 6458
rect 7380 6394 7432 6400
rect 7484 6202 7512 9114
rect 7852 9042 7880 9658
rect 7840 9036 7892 9042
rect 7840 8978 7892 8984
rect 7852 8820 7880 8978
rect 7760 8792 7880 8820
rect 7562 8664 7618 8673
rect 7760 8634 7788 8792
rect 7896 8732 8204 8741
rect 7896 8730 7902 8732
rect 7958 8730 7982 8732
rect 8038 8730 8062 8732
rect 8118 8730 8142 8732
rect 8198 8730 8204 8732
rect 7958 8678 7960 8730
rect 8140 8678 8142 8730
rect 7896 8676 7902 8678
rect 7958 8676 7982 8678
rect 8038 8676 8062 8678
rect 8118 8676 8142 8678
rect 8198 8676 8204 8678
rect 7896 8667 8204 8676
rect 7562 8599 7618 8608
rect 7748 8628 7800 8634
rect 7576 6338 7604 8599
rect 7748 8570 7800 8576
rect 7760 8514 7788 8570
rect 7668 8486 7788 8514
rect 8298 8528 8354 8537
rect 7668 8294 7696 8486
rect 8298 8463 8354 8472
rect 7748 8424 7800 8430
rect 7748 8366 7800 8372
rect 7656 8288 7708 8294
rect 7656 8230 7708 8236
rect 7668 7954 7696 8230
rect 7656 7948 7708 7954
rect 7656 7890 7708 7896
rect 7656 6656 7708 6662
rect 7656 6598 7708 6604
rect 7668 6458 7696 6598
rect 7656 6452 7708 6458
rect 7760 6440 7788 8366
rect 8312 7954 8340 8463
rect 8208 7948 8260 7954
rect 8208 7890 8260 7896
rect 8300 7948 8352 7954
rect 8300 7890 8352 7896
rect 8220 7732 8248 7890
rect 8220 7704 8340 7732
rect 7896 7644 8204 7653
rect 7896 7642 7902 7644
rect 7958 7642 7982 7644
rect 8038 7642 8062 7644
rect 8118 7642 8142 7644
rect 8198 7642 8204 7644
rect 7958 7590 7960 7642
rect 8140 7590 8142 7642
rect 7896 7588 7902 7590
rect 7958 7588 7982 7590
rect 8038 7588 8062 7590
rect 8118 7588 8142 7590
rect 8198 7588 8204 7590
rect 7896 7579 8204 7588
rect 8312 7426 8340 7704
rect 8404 7546 8432 11086
rect 8496 10266 8524 13110
rect 8484 10260 8536 10266
rect 8484 10202 8536 10208
rect 8496 9586 8524 10202
rect 8484 9580 8536 9586
rect 8484 9522 8536 9528
rect 8482 8936 8538 8945
rect 8482 8871 8538 8880
rect 8392 7540 8444 7546
rect 8392 7482 8444 7488
rect 8220 7398 8340 7426
rect 7838 7168 7894 7177
rect 7838 7103 7894 7112
rect 7852 7002 7880 7103
rect 7840 6996 7892 7002
rect 7840 6938 7892 6944
rect 8024 6792 8076 6798
rect 8116 6792 8168 6798
rect 8024 6734 8076 6740
rect 8114 6760 8116 6769
rect 8168 6760 8170 6769
rect 8036 6662 8064 6734
rect 8220 6746 8248 7398
rect 8220 6718 8432 6746
rect 8114 6695 8170 6704
rect 8024 6656 8076 6662
rect 8024 6598 8076 6604
rect 7896 6556 8204 6565
rect 7896 6554 7902 6556
rect 7958 6554 7982 6556
rect 8038 6554 8062 6556
rect 8118 6554 8142 6556
rect 8198 6554 8204 6556
rect 7958 6502 7960 6554
rect 8140 6502 8142 6554
rect 7896 6500 7902 6502
rect 7958 6500 7982 6502
rect 8038 6500 8062 6502
rect 8118 6500 8142 6502
rect 8198 6500 8204 6502
rect 7896 6491 8204 6500
rect 8300 6452 8352 6458
rect 7760 6412 7972 6440
rect 7656 6394 7708 6400
rect 7576 6310 7788 6338
rect 7392 6174 7512 6202
rect 7392 5001 7420 6174
rect 7472 6112 7524 6118
rect 7472 6054 7524 6060
rect 7484 5710 7512 6054
rect 7472 5704 7524 5710
rect 7472 5646 7524 5652
rect 7564 5704 7616 5710
rect 7760 5658 7788 6310
rect 7944 5846 7972 6412
rect 8300 6394 8352 6400
rect 8312 5914 8340 6394
rect 8404 5914 8432 6718
rect 8496 6662 8524 8871
rect 8588 8634 8616 16526
rect 8772 15366 8800 17070
rect 8760 15360 8812 15366
rect 8760 15302 8812 15308
rect 8772 13802 8800 15302
rect 8760 13796 8812 13802
rect 8760 13738 8812 13744
rect 8668 13728 8720 13734
rect 8668 13670 8720 13676
rect 8680 13394 8708 13670
rect 8760 13524 8812 13530
rect 8760 13466 8812 13472
rect 8668 13388 8720 13394
rect 8668 13330 8720 13336
rect 8668 13184 8720 13190
rect 8668 13126 8720 13132
rect 8680 12918 8708 13126
rect 8772 12986 8800 13466
rect 8760 12980 8812 12986
rect 8760 12922 8812 12928
rect 8668 12912 8720 12918
rect 8668 12854 8720 12860
rect 8758 12472 8814 12481
rect 8758 12407 8814 12416
rect 8864 12434 8892 17274
rect 9324 16658 9352 17478
rect 9312 16652 9364 16658
rect 9312 16594 9364 16600
rect 9128 13864 9180 13870
rect 9128 13806 9180 13812
rect 9312 13864 9364 13870
rect 9312 13806 9364 13812
rect 9140 13530 9168 13806
rect 9128 13524 9180 13530
rect 9128 13466 9180 13472
rect 9036 13388 9088 13394
rect 9036 13330 9088 13336
rect 8772 12306 8800 12407
rect 8864 12406 8984 12434
rect 8760 12300 8812 12306
rect 8760 12242 8812 12248
rect 8668 12096 8720 12102
rect 8668 12038 8720 12044
rect 8852 12096 8904 12102
rect 8852 12038 8904 12044
rect 8680 11694 8708 12038
rect 8864 11898 8892 12038
rect 8852 11892 8904 11898
rect 8852 11834 8904 11840
rect 8760 11824 8812 11830
rect 8760 11766 8812 11772
rect 8668 11688 8720 11694
rect 8668 11630 8720 11636
rect 8668 11552 8720 11558
rect 8772 11540 8800 11766
rect 8720 11512 8800 11540
rect 8668 11494 8720 11500
rect 8850 11384 8906 11393
rect 8850 11319 8906 11328
rect 8864 11218 8892 11319
rect 8956 11218 8984 12406
rect 9048 12374 9076 13330
rect 9128 13320 9180 13326
rect 9128 13262 9180 13268
rect 9036 12368 9088 12374
rect 9036 12310 9088 12316
rect 9048 11558 9076 12310
rect 9036 11552 9088 11558
rect 9036 11494 9088 11500
rect 8852 11212 8904 11218
rect 8852 11154 8904 11160
rect 8944 11212 8996 11218
rect 8944 11154 8996 11160
rect 8668 10056 8720 10062
rect 8668 9998 8720 10004
rect 8576 8628 8628 8634
rect 8576 8570 8628 8576
rect 8680 8514 8708 9998
rect 8944 8968 8996 8974
rect 8944 8910 8996 8916
rect 8588 8486 8708 8514
rect 8588 8430 8616 8486
rect 8576 8424 8628 8430
rect 8576 8366 8628 8372
rect 8588 8294 8616 8366
rect 8588 8266 8708 8294
rect 8576 7812 8628 7818
rect 8576 7754 8628 7760
rect 8588 7478 8616 7754
rect 8576 7472 8628 7478
rect 8576 7414 8628 7420
rect 8680 7206 8708 8266
rect 8760 7336 8812 7342
rect 8760 7278 8812 7284
rect 8668 7200 8720 7206
rect 8668 7142 8720 7148
rect 8680 6905 8708 7142
rect 8666 6896 8722 6905
rect 8666 6831 8668 6840
rect 8720 6831 8722 6840
rect 8668 6802 8720 6808
rect 8484 6656 8536 6662
rect 8484 6598 8536 6604
rect 8680 6202 8708 6802
rect 8496 6174 8708 6202
rect 8300 5908 8352 5914
rect 8300 5850 8352 5856
rect 8392 5908 8444 5914
rect 8392 5850 8444 5856
rect 7840 5840 7892 5846
rect 7840 5782 7892 5788
rect 7932 5840 7984 5846
rect 7932 5782 7984 5788
rect 8024 5840 8076 5846
rect 8024 5782 8076 5788
rect 7852 5692 7880 5782
rect 8036 5692 8064 5782
rect 7852 5664 8064 5692
rect 7564 5646 7616 5652
rect 7378 4992 7434 5001
rect 7378 4927 7434 4936
rect 7472 3528 7524 3534
rect 7472 3470 7524 3476
rect 7484 3058 7512 3470
rect 7576 3194 7604 5646
rect 7668 5630 7788 5658
rect 7668 3534 7696 5630
rect 7896 5468 8204 5477
rect 7896 5466 7902 5468
rect 7958 5466 7982 5468
rect 8038 5466 8062 5468
rect 8118 5466 8142 5468
rect 8198 5466 8204 5468
rect 7958 5414 7960 5466
rect 8140 5414 8142 5466
rect 7896 5412 7902 5414
rect 7958 5412 7982 5414
rect 8038 5412 8062 5414
rect 8118 5412 8142 5414
rect 8198 5412 8204 5414
rect 7896 5403 8204 5412
rect 8496 5370 8524 6174
rect 8576 6112 8628 6118
rect 8576 6054 8628 6060
rect 8484 5364 8536 5370
rect 8484 5306 8536 5312
rect 7748 5296 7800 5302
rect 7800 5256 7972 5284
rect 7748 5238 7800 5244
rect 7840 5160 7892 5166
rect 7840 5102 7892 5108
rect 7852 4570 7880 5102
rect 7944 4740 7972 5256
rect 8114 5264 8170 5273
rect 8170 5234 8294 5250
rect 8170 5228 8306 5234
rect 8170 5222 8254 5228
rect 8114 5199 8170 5208
rect 8254 5170 8306 5176
rect 8392 5228 8444 5234
rect 8392 5170 8444 5176
rect 8484 5228 8536 5234
rect 8484 5170 8536 5176
rect 8116 5092 8168 5098
rect 8116 5034 8168 5040
rect 8024 4752 8076 4758
rect 7944 4712 8024 4740
rect 8128 4729 8156 5034
rect 8208 5024 8260 5030
rect 8206 4992 8208 5001
rect 8260 4992 8262 5001
rect 8206 4927 8262 4936
rect 8024 4694 8076 4700
rect 8114 4720 8170 4729
rect 8114 4655 8170 4664
rect 7760 4542 7880 4570
rect 7760 3738 7788 4542
rect 7896 4380 8204 4389
rect 7896 4378 7902 4380
rect 7958 4378 7982 4380
rect 8038 4378 8062 4380
rect 8118 4378 8142 4380
rect 8198 4378 8204 4380
rect 7958 4326 7960 4378
rect 8140 4326 8142 4378
rect 7896 4324 7902 4326
rect 7958 4324 7982 4326
rect 8038 4324 8062 4326
rect 8118 4324 8142 4326
rect 8198 4324 8204 4326
rect 7896 4315 8204 4324
rect 8300 4004 8352 4010
rect 8300 3946 8352 3952
rect 7748 3732 7800 3738
rect 7748 3674 7800 3680
rect 7656 3528 7708 3534
rect 7932 3528 7984 3534
rect 7656 3470 7708 3476
rect 7760 3488 7932 3516
rect 7564 3188 7616 3194
rect 7564 3130 7616 3136
rect 7472 3052 7524 3058
rect 7472 2994 7524 3000
rect 7380 2984 7432 2990
rect 7380 2926 7432 2932
rect 7024 2746 7328 2774
rect 7024 2650 7052 2746
rect 7012 2644 7064 2650
rect 7012 2586 7064 2592
rect 7104 2576 7156 2582
rect 7104 2518 7156 2524
rect 7116 800 7144 2518
rect 7392 800 7420 2926
rect 7656 2372 7708 2378
rect 7656 2314 7708 2320
rect 7668 800 7696 2314
rect 7760 1442 7788 3488
rect 7932 3470 7984 3476
rect 7896 3292 8204 3301
rect 7896 3290 7902 3292
rect 7958 3290 7982 3292
rect 8038 3290 8062 3292
rect 8118 3290 8142 3292
rect 8198 3290 8204 3292
rect 7958 3238 7960 3290
rect 8140 3238 8142 3290
rect 7896 3236 7902 3238
rect 7958 3236 7982 3238
rect 8038 3236 8062 3238
rect 8118 3236 8142 3238
rect 8198 3236 8204 3238
rect 7896 3227 8204 3236
rect 8208 2984 8260 2990
rect 8208 2926 8260 2932
rect 8220 2394 8248 2926
rect 8312 2854 8340 3946
rect 8404 3194 8432 5170
rect 8496 3738 8524 5170
rect 8588 5030 8616 6054
rect 8668 5704 8720 5710
rect 8668 5646 8720 5652
rect 8576 5024 8628 5030
rect 8576 4966 8628 4972
rect 8576 4208 8628 4214
rect 8576 4150 8628 4156
rect 8588 4049 8616 4150
rect 8574 4040 8630 4049
rect 8574 3975 8630 3984
rect 8484 3732 8536 3738
rect 8484 3674 8536 3680
rect 8392 3188 8444 3194
rect 8392 3130 8444 3136
rect 8300 2848 8352 2854
rect 8300 2790 8352 2796
rect 8484 2440 8536 2446
rect 8220 2366 8340 2394
rect 8484 2382 8536 2388
rect 7896 2204 8204 2213
rect 7896 2202 7902 2204
rect 7958 2202 7982 2204
rect 8038 2202 8062 2204
rect 8118 2202 8142 2204
rect 8198 2202 8204 2204
rect 7958 2150 7960 2202
rect 8140 2150 8142 2202
rect 7896 2148 7902 2150
rect 7958 2148 7982 2150
rect 8038 2148 8062 2150
rect 8118 2148 8142 2150
rect 8198 2148 8204 2150
rect 7896 2139 8204 2148
rect 8312 1986 8340 2366
rect 8220 1958 8340 1986
rect 7760 1414 7972 1442
rect 7944 800 7972 1414
rect 8220 800 8248 1958
rect 8496 800 8524 2382
rect 8680 1698 8708 5646
rect 8772 5370 8800 7278
rect 8956 6458 8984 8910
rect 9140 8090 9168 13262
rect 9324 12434 9352 13806
rect 9232 12406 9352 12434
rect 9232 10062 9260 12406
rect 9312 12164 9364 12170
rect 9312 12106 9364 12112
rect 9324 11218 9352 12106
rect 9312 11212 9364 11218
rect 9312 11154 9364 11160
rect 9220 10056 9272 10062
rect 9220 9998 9272 10004
rect 9416 9654 9444 18226
rect 9772 17808 9824 17814
rect 9772 17750 9824 17756
rect 9876 17762 9904 18226
rect 10140 18216 10192 18222
rect 10140 18158 10192 18164
rect 10048 18080 10100 18086
rect 10048 18022 10100 18028
rect 9784 17202 9812 17750
rect 9876 17734 9996 17762
rect 9864 17672 9916 17678
rect 9864 17614 9916 17620
rect 9876 17338 9904 17614
rect 9864 17332 9916 17338
rect 9864 17274 9916 17280
rect 9772 17196 9824 17202
rect 9772 17138 9824 17144
rect 9680 15904 9732 15910
rect 9680 15846 9732 15852
rect 9692 15434 9720 15846
rect 9784 15586 9812 17138
rect 9864 16516 9916 16522
rect 9864 16458 9916 16464
rect 9876 15706 9904 16458
rect 9864 15700 9916 15706
rect 9864 15642 9916 15648
rect 9784 15558 9904 15586
rect 9680 15428 9732 15434
rect 9680 15370 9732 15376
rect 9692 15026 9720 15370
rect 9680 15020 9732 15026
rect 9680 14962 9732 14968
rect 9692 14498 9720 14962
rect 9772 14884 9824 14890
rect 9772 14826 9824 14832
rect 9600 14470 9720 14498
rect 9784 14482 9812 14826
rect 9772 14476 9824 14482
rect 9600 13938 9628 14470
rect 9772 14418 9824 14424
rect 9680 14408 9732 14414
rect 9680 14350 9732 14356
rect 9692 14074 9720 14350
rect 9772 14272 9824 14278
rect 9772 14214 9824 14220
rect 9680 14068 9732 14074
rect 9680 14010 9732 14016
rect 9496 13932 9548 13938
rect 9496 13874 9548 13880
rect 9588 13932 9640 13938
rect 9588 13874 9640 13880
rect 9508 11762 9536 13874
rect 9600 12889 9628 13874
rect 9680 13728 9732 13734
rect 9680 13670 9732 13676
rect 9586 12880 9642 12889
rect 9692 12850 9720 13670
rect 9784 13394 9812 14214
rect 9772 13388 9824 13394
rect 9772 13330 9824 13336
rect 9586 12815 9642 12824
rect 9680 12844 9732 12850
rect 9680 12786 9732 12792
rect 9772 12708 9824 12714
rect 9772 12650 9824 12656
rect 9784 12345 9812 12650
rect 9770 12336 9826 12345
rect 9770 12271 9826 12280
rect 9876 12238 9904 15558
rect 9864 12232 9916 12238
rect 9864 12174 9916 12180
rect 9588 12096 9640 12102
rect 9588 12038 9640 12044
rect 9600 11830 9628 12038
rect 9588 11824 9640 11830
rect 9588 11766 9640 11772
rect 9876 11762 9904 12174
rect 9496 11756 9548 11762
rect 9496 11698 9548 11704
rect 9864 11756 9916 11762
rect 9864 11698 9916 11704
rect 9588 11620 9640 11626
rect 9588 11562 9640 11568
rect 9496 11552 9548 11558
rect 9496 11494 9548 11500
rect 9404 9648 9456 9654
rect 9404 9590 9456 9596
rect 9508 9466 9536 11494
rect 9600 11393 9628 11562
rect 9586 11384 9642 11393
rect 9586 11319 9642 11328
rect 9968 11200 9996 17734
rect 10060 17338 10088 18022
rect 10048 17332 10100 17338
rect 10048 17274 10100 17280
rect 10046 14512 10102 14521
rect 10046 14447 10102 14456
rect 10060 14006 10088 14447
rect 10048 14000 10100 14006
rect 10048 13942 10100 13948
rect 10060 11898 10088 13942
rect 10152 13938 10180 18158
rect 10244 17746 10272 22374
rect 11369 22332 11677 22341
rect 11369 22330 11375 22332
rect 11431 22330 11455 22332
rect 11511 22330 11535 22332
rect 11591 22330 11615 22332
rect 11671 22330 11677 22332
rect 11431 22278 11433 22330
rect 11613 22278 11615 22330
rect 11369 22276 11375 22278
rect 11431 22276 11455 22278
rect 11511 22276 11535 22278
rect 11591 22276 11615 22278
rect 11671 22276 11677 22278
rect 11369 22267 11677 22276
rect 11369 21244 11677 21253
rect 11369 21242 11375 21244
rect 11431 21242 11455 21244
rect 11511 21242 11535 21244
rect 11591 21242 11615 21244
rect 11671 21242 11677 21244
rect 11431 21190 11433 21242
rect 11613 21190 11615 21242
rect 11369 21188 11375 21190
rect 11431 21188 11455 21190
rect 11511 21188 11535 21190
rect 11591 21188 11615 21190
rect 11671 21188 11677 21190
rect 11369 21179 11677 21188
rect 11369 20156 11677 20165
rect 11369 20154 11375 20156
rect 11431 20154 11455 20156
rect 11511 20154 11535 20156
rect 11591 20154 11615 20156
rect 11671 20154 11677 20156
rect 11431 20102 11433 20154
rect 11613 20102 11615 20154
rect 11369 20100 11375 20102
rect 11431 20100 11455 20102
rect 11511 20100 11535 20102
rect 11591 20100 11615 20102
rect 11671 20100 11677 20102
rect 11369 20091 11677 20100
rect 10784 19712 10836 19718
rect 10784 19654 10836 19660
rect 10600 18284 10652 18290
rect 10600 18226 10652 18232
rect 10508 18216 10560 18222
rect 10508 18158 10560 18164
rect 10232 17740 10284 17746
rect 10232 17682 10284 17688
rect 10416 17672 10468 17678
rect 10416 17614 10468 17620
rect 10324 16040 10376 16046
rect 10324 15982 10376 15988
rect 10336 15366 10364 15982
rect 10324 15360 10376 15366
rect 10324 15302 10376 15308
rect 10428 15042 10456 17614
rect 10520 17134 10548 18158
rect 10612 17882 10640 18226
rect 10600 17876 10652 17882
rect 10600 17818 10652 17824
rect 10796 17814 10824 19654
rect 11369 19068 11677 19077
rect 11369 19066 11375 19068
rect 11431 19066 11455 19068
rect 11511 19066 11535 19068
rect 11591 19066 11615 19068
rect 11671 19066 11677 19068
rect 11431 19014 11433 19066
rect 11613 19014 11615 19066
rect 11369 19012 11375 19014
rect 11431 19012 11455 19014
rect 11511 19012 11535 19014
rect 11591 19012 11615 19014
rect 11671 19012 11677 19014
rect 11369 19003 11677 19012
rect 12820 18970 12848 24550
rect 12808 18964 12860 18970
rect 12808 18906 12860 18912
rect 12820 18426 12848 18906
rect 12808 18420 12860 18426
rect 12808 18362 12860 18368
rect 13728 18420 13780 18426
rect 13728 18362 13780 18368
rect 10876 18148 10928 18154
rect 10876 18090 10928 18096
rect 10784 17808 10836 17814
rect 10784 17750 10836 17756
rect 10692 17672 10744 17678
rect 10692 17614 10744 17620
rect 10704 17338 10732 17614
rect 10692 17332 10744 17338
rect 10692 17274 10744 17280
rect 10508 17128 10560 17134
rect 10508 17070 10560 17076
rect 10796 16658 10824 17750
rect 10888 17338 10916 18090
rect 12716 18080 12768 18086
rect 12716 18022 12768 18028
rect 11369 17980 11677 17989
rect 11369 17978 11375 17980
rect 11431 17978 11455 17980
rect 11511 17978 11535 17980
rect 11591 17978 11615 17980
rect 11671 17978 11677 17980
rect 11431 17926 11433 17978
rect 11613 17926 11615 17978
rect 11369 17924 11375 17926
rect 11431 17924 11455 17926
rect 11511 17924 11535 17926
rect 11591 17924 11615 17926
rect 11671 17924 11677 17926
rect 11369 17915 11677 17924
rect 11704 17740 11756 17746
rect 11704 17682 11756 17688
rect 11796 17740 11848 17746
rect 11796 17682 11848 17688
rect 10876 17332 10928 17338
rect 10876 17274 10928 17280
rect 10968 17196 11020 17202
rect 10968 17138 11020 17144
rect 10980 16794 11008 17138
rect 11716 17134 11744 17682
rect 11808 17338 11836 17682
rect 12728 17338 12756 18022
rect 13176 17604 13228 17610
rect 13176 17546 13228 17552
rect 11796 17332 11848 17338
rect 11796 17274 11848 17280
rect 12716 17332 12768 17338
rect 12716 17274 12768 17280
rect 11152 17128 11204 17134
rect 11152 17070 11204 17076
rect 11704 17128 11756 17134
rect 11704 17070 11756 17076
rect 10968 16788 11020 16794
rect 10968 16730 11020 16736
rect 11060 16720 11112 16726
rect 11060 16662 11112 16668
rect 10784 16652 10836 16658
rect 10784 16594 10836 16600
rect 10968 16040 11020 16046
rect 10968 15982 11020 15988
rect 10980 15706 11008 15982
rect 10968 15700 11020 15706
rect 10968 15642 11020 15648
rect 11072 15570 11100 16662
rect 11164 15706 11192 17070
rect 11369 16892 11677 16901
rect 11369 16890 11375 16892
rect 11431 16890 11455 16892
rect 11511 16890 11535 16892
rect 11591 16890 11615 16892
rect 11671 16890 11677 16892
rect 11431 16838 11433 16890
rect 11613 16838 11615 16890
rect 11369 16836 11375 16838
rect 11431 16836 11455 16838
rect 11511 16836 11535 16838
rect 11591 16836 11615 16838
rect 11671 16836 11677 16838
rect 11369 16827 11677 16836
rect 11716 16590 11744 17070
rect 11704 16584 11756 16590
rect 11704 16526 11756 16532
rect 11336 16448 11388 16454
rect 11336 16390 11388 16396
rect 11520 16448 11572 16454
rect 11520 16390 11572 16396
rect 11348 16114 11376 16390
rect 11532 16250 11560 16390
rect 11520 16244 11572 16250
rect 11520 16186 11572 16192
rect 11716 16182 11744 16526
rect 11704 16176 11756 16182
rect 11704 16118 11756 16124
rect 13084 16176 13136 16182
rect 13084 16118 13136 16124
rect 11336 16108 11388 16114
rect 11336 16050 11388 16056
rect 11369 15804 11677 15813
rect 11369 15802 11375 15804
rect 11431 15802 11455 15804
rect 11511 15802 11535 15804
rect 11591 15802 11615 15804
rect 11671 15802 11677 15804
rect 11431 15750 11433 15802
rect 11613 15750 11615 15802
rect 11369 15748 11375 15750
rect 11431 15748 11455 15750
rect 11511 15748 11535 15750
rect 11591 15748 11615 15750
rect 11671 15748 11677 15750
rect 11369 15739 11677 15748
rect 11152 15700 11204 15706
rect 11152 15642 11204 15648
rect 11060 15564 11112 15570
rect 11060 15506 11112 15512
rect 10428 15014 10548 15042
rect 10324 14408 10376 14414
rect 10324 14350 10376 14356
rect 10416 14408 10468 14414
rect 10416 14350 10468 14356
rect 10140 13932 10192 13938
rect 10140 13874 10192 13880
rect 10336 12782 10364 14350
rect 10428 14074 10456 14350
rect 10416 14068 10468 14074
rect 10416 14010 10468 14016
rect 10416 13864 10468 13870
rect 10416 13806 10468 13812
rect 10428 12986 10456 13806
rect 10416 12980 10468 12986
rect 10416 12922 10468 12928
rect 10324 12776 10376 12782
rect 10324 12718 10376 12724
rect 10416 12096 10468 12102
rect 10416 12038 10468 12044
rect 10428 11898 10456 12038
rect 10048 11892 10100 11898
rect 10048 11834 10100 11840
rect 10416 11892 10468 11898
rect 10416 11834 10468 11840
rect 10060 11218 10088 11834
rect 9876 11172 9996 11200
rect 10048 11212 10100 11218
rect 9588 11144 9640 11150
rect 9588 11086 9640 11092
rect 9416 9438 9536 9466
rect 9312 9036 9364 9042
rect 9312 8978 9364 8984
rect 9220 8900 9272 8906
rect 9220 8842 9272 8848
rect 9232 8634 9260 8842
rect 9220 8628 9272 8634
rect 9220 8570 9272 8576
rect 9128 8084 9180 8090
rect 9128 8026 9180 8032
rect 9128 7812 9180 7818
rect 9128 7754 9180 7760
rect 9140 7410 9168 7754
rect 9128 7404 9180 7410
rect 9128 7346 9180 7352
rect 9220 7404 9272 7410
rect 9220 7346 9272 7352
rect 9036 7336 9088 7342
rect 9036 7278 9088 7284
rect 9048 6866 9076 7278
rect 9036 6860 9088 6866
rect 9036 6802 9088 6808
rect 9048 6474 9076 6802
rect 8944 6452 8996 6458
rect 9048 6446 9168 6474
rect 8944 6394 8996 6400
rect 9036 6384 9088 6390
rect 9036 6326 9088 6332
rect 9048 5914 9076 6326
rect 9140 5914 9168 6446
rect 9232 6254 9260 7346
rect 9324 7290 9352 8978
rect 9416 7410 9444 9438
rect 9496 9376 9548 9382
rect 9496 9318 9548 9324
rect 9404 7404 9456 7410
rect 9404 7346 9456 7352
rect 9324 7262 9444 7290
rect 9312 7200 9364 7206
rect 9312 7142 9364 7148
rect 9324 7002 9352 7142
rect 9312 6996 9364 7002
rect 9312 6938 9364 6944
rect 9220 6248 9272 6254
rect 9220 6190 9272 6196
rect 9036 5908 9088 5914
rect 9036 5850 9088 5856
rect 9128 5908 9180 5914
rect 9128 5850 9180 5856
rect 8760 5364 8812 5370
rect 8760 5306 8812 5312
rect 9036 5364 9088 5370
rect 9036 5306 9088 5312
rect 8944 5228 8996 5234
rect 8944 5170 8996 5176
rect 8852 5024 8904 5030
rect 8852 4966 8904 4972
rect 8760 4548 8812 4554
rect 8760 4490 8812 4496
rect 8772 4321 8800 4490
rect 8758 4312 8814 4321
rect 8758 4247 8814 4256
rect 8760 4004 8812 4010
rect 8760 3946 8812 3952
rect 8772 3398 8800 3946
rect 8864 3738 8892 4966
rect 8852 3732 8904 3738
rect 8852 3674 8904 3680
rect 8760 3392 8812 3398
rect 8760 3334 8812 3340
rect 8760 2984 8812 2990
rect 8760 2926 8812 2932
rect 8668 1692 8720 1698
rect 8668 1634 8720 1640
rect 8772 800 8800 2926
rect 8852 2440 8904 2446
rect 8852 2382 8904 2388
rect 8864 1306 8892 2382
rect 8956 2310 8984 5170
rect 9048 4690 9076 5306
rect 9220 5228 9272 5234
rect 9220 5170 9272 5176
rect 9036 4684 9088 4690
rect 9036 4626 9088 4632
rect 9232 4282 9260 5170
rect 9416 4826 9444 7262
rect 9508 6186 9536 9318
rect 9600 6866 9628 11086
rect 9772 11008 9824 11014
rect 9772 10950 9824 10956
rect 9680 10736 9732 10742
rect 9680 10678 9732 10684
rect 9692 10198 9720 10678
rect 9680 10192 9732 10198
rect 9680 10134 9732 10140
rect 9680 9512 9732 9518
rect 9680 9454 9732 9460
rect 9692 9042 9720 9454
rect 9784 9081 9812 10950
rect 9876 10266 9904 11172
rect 10048 11154 10100 11160
rect 10232 11008 10284 11014
rect 10232 10950 10284 10956
rect 9956 10532 10008 10538
rect 9956 10474 10008 10480
rect 9864 10260 9916 10266
rect 9864 10202 9916 10208
rect 9968 10130 9996 10474
rect 10048 10464 10100 10470
rect 10048 10406 10100 10412
rect 10140 10464 10192 10470
rect 10140 10406 10192 10412
rect 10060 10266 10088 10406
rect 10048 10260 10100 10266
rect 10048 10202 10100 10208
rect 9956 10124 10008 10130
rect 9956 10066 10008 10072
rect 9864 10056 9916 10062
rect 9864 9998 9916 10004
rect 9876 9330 9904 9998
rect 10152 9994 10180 10406
rect 10140 9988 10192 9994
rect 10140 9930 10192 9936
rect 10140 9648 10192 9654
rect 10140 9590 10192 9596
rect 10046 9480 10102 9489
rect 10046 9415 10048 9424
rect 10100 9415 10102 9424
rect 10048 9386 10100 9392
rect 9876 9302 9996 9330
rect 9864 9172 9916 9178
rect 9864 9114 9916 9120
rect 9770 9072 9826 9081
rect 9680 9036 9732 9042
rect 9770 9007 9826 9016
rect 9680 8978 9732 8984
rect 9772 8900 9824 8906
rect 9772 8842 9824 8848
rect 9680 7880 9732 7886
rect 9680 7822 9732 7828
rect 9588 6860 9640 6866
rect 9588 6802 9640 6808
rect 9496 6180 9548 6186
rect 9496 6122 9548 6128
rect 9692 5574 9720 7822
rect 9784 7546 9812 8842
rect 9772 7540 9824 7546
rect 9772 7482 9824 7488
rect 9770 7440 9826 7449
rect 9876 7410 9904 9114
rect 9770 7375 9826 7384
rect 9864 7404 9916 7410
rect 9784 7342 9812 7375
rect 9864 7346 9916 7352
rect 9772 7336 9824 7342
rect 9772 7278 9824 7284
rect 9772 6860 9824 6866
rect 9772 6802 9824 6808
rect 9784 6458 9812 6802
rect 9772 6452 9824 6458
rect 9772 6394 9824 6400
rect 9864 6452 9916 6458
rect 9864 6394 9916 6400
rect 9876 5914 9904 6394
rect 9864 5908 9916 5914
rect 9864 5850 9916 5856
rect 9876 5710 9904 5850
rect 9864 5704 9916 5710
rect 9864 5646 9916 5652
rect 9680 5568 9732 5574
rect 9680 5510 9732 5516
rect 9876 5302 9904 5646
rect 9864 5296 9916 5302
rect 9864 5238 9916 5244
rect 9876 4826 9904 5238
rect 9404 4820 9456 4826
rect 9864 4820 9916 4826
rect 9404 4762 9456 4768
rect 9784 4780 9864 4808
rect 9404 4616 9456 4622
rect 9404 4558 9456 4564
rect 9680 4616 9732 4622
rect 9680 4558 9732 4564
rect 9312 4480 9364 4486
rect 9312 4422 9364 4428
rect 9324 4282 9352 4422
rect 9220 4276 9272 4282
rect 9220 4218 9272 4224
rect 9312 4276 9364 4282
rect 9312 4218 9364 4224
rect 9310 4176 9366 4185
rect 9310 4111 9312 4120
rect 9364 4111 9366 4120
rect 9312 4082 9364 4088
rect 9324 3126 9352 4082
rect 9416 3194 9444 4558
rect 9692 4214 9720 4558
rect 9784 4214 9812 4780
rect 9864 4762 9916 4768
rect 9862 4312 9918 4321
rect 9862 4247 9918 4256
rect 9876 4214 9904 4247
rect 9680 4208 9732 4214
rect 9680 4150 9732 4156
rect 9772 4208 9824 4214
rect 9772 4150 9824 4156
rect 9864 4208 9916 4214
rect 9864 4150 9916 4156
rect 9588 3936 9640 3942
rect 9588 3878 9640 3884
rect 9600 3641 9628 3878
rect 9586 3632 9642 3641
rect 9586 3567 9642 3576
rect 9588 3528 9640 3534
rect 9588 3470 9640 3476
rect 9404 3188 9456 3194
rect 9404 3130 9456 3136
rect 9312 3120 9364 3126
rect 9312 3062 9364 3068
rect 9220 2984 9272 2990
rect 9220 2926 9272 2932
rect 9496 2984 9548 2990
rect 9496 2926 9548 2932
rect 9232 2774 9260 2926
rect 9232 2746 9352 2774
rect 8944 2304 8996 2310
rect 8944 2246 8996 2252
rect 8864 1278 9076 1306
rect 9048 800 9076 1278
rect 9324 800 9352 2746
rect 9508 2514 9536 2926
rect 9496 2508 9548 2514
rect 9496 2450 9548 2456
rect 9600 800 9628 3470
rect 9968 3126 9996 9302
rect 10048 7744 10100 7750
rect 10048 7686 10100 7692
rect 10060 7546 10088 7686
rect 10048 7540 10100 7546
rect 10048 7482 10100 7488
rect 10048 4072 10100 4078
rect 10048 4014 10100 4020
rect 10060 3670 10088 4014
rect 10152 3942 10180 9590
rect 10244 9110 10272 10950
rect 10520 10810 10548 15014
rect 10968 14884 11020 14890
rect 10968 14826 11020 14832
rect 10980 14414 11008 14826
rect 11369 14716 11677 14725
rect 11369 14714 11375 14716
rect 11431 14714 11455 14716
rect 11511 14714 11535 14716
rect 11591 14714 11615 14716
rect 11671 14714 11677 14716
rect 11431 14662 11433 14714
rect 11613 14662 11615 14714
rect 11369 14660 11375 14662
rect 11431 14660 11455 14662
rect 11511 14660 11535 14662
rect 11591 14660 11615 14662
rect 11671 14660 11677 14662
rect 11369 14651 11677 14660
rect 10784 14408 10836 14414
rect 10784 14350 10836 14356
rect 10968 14408 11020 14414
rect 10968 14350 11020 14356
rect 11244 14408 11296 14414
rect 11716 14396 11744 16118
rect 11796 16040 11848 16046
rect 11796 15982 11848 15988
rect 11808 15706 11836 15982
rect 13096 15706 13124 16118
rect 13188 15706 13216 17546
rect 13740 17202 13768 18362
rect 13728 17196 13780 17202
rect 13728 17138 13780 17144
rect 13636 16788 13688 16794
rect 13636 16730 13688 16736
rect 13648 16590 13676 16730
rect 13636 16584 13688 16590
rect 13636 16526 13688 16532
rect 13268 16516 13320 16522
rect 13268 16458 13320 16464
rect 13280 16250 13308 16458
rect 13268 16244 13320 16250
rect 13268 16186 13320 16192
rect 13268 15904 13320 15910
rect 13268 15846 13320 15852
rect 11796 15700 11848 15706
rect 11796 15642 11848 15648
rect 13084 15700 13136 15706
rect 13084 15642 13136 15648
rect 13176 15700 13228 15706
rect 13176 15642 13228 15648
rect 13280 15638 13308 15846
rect 13268 15632 13320 15638
rect 13268 15574 13320 15580
rect 12256 15564 12308 15570
rect 12256 15506 12308 15512
rect 11888 15088 11940 15094
rect 11888 15030 11940 15036
rect 11900 14618 11928 15030
rect 12268 14958 12296 15506
rect 13268 15496 13320 15502
rect 13268 15438 13320 15444
rect 12348 15360 12400 15366
rect 12348 15302 12400 15308
rect 12256 14952 12308 14958
rect 12256 14894 12308 14900
rect 11888 14612 11940 14618
rect 11888 14554 11940 14560
rect 11888 14408 11940 14414
rect 11716 14368 11888 14396
rect 11244 14350 11296 14356
rect 11888 14350 11940 14356
rect 10692 13252 10744 13258
rect 10692 13194 10744 13200
rect 10704 12986 10732 13194
rect 10692 12980 10744 12986
rect 10692 12922 10744 12928
rect 10600 12844 10652 12850
rect 10600 12786 10652 12792
rect 10612 12434 10640 12786
rect 10612 12406 10732 12434
rect 10600 12368 10652 12374
rect 10600 12310 10652 12316
rect 10508 10804 10560 10810
rect 10508 10746 10560 10752
rect 10416 10736 10468 10742
rect 10416 10678 10468 10684
rect 10324 10600 10376 10606
rect 10324 10542 10376 10548
rect 10336 9382 10364 10542
rect 10428 9625 10456 10678
rect 10414 9616 10470 9625
rect 10414 9551 10470 9560
rect 10508 9512 10560 9518
rect 10506 9480 10508 9489
rect 10560 9480 10562 9489
rect 10506 9415 10562 9424
rect 10324 9376 10376 9382
rect 10324 9318 10376 9324
rect 10612 9178 10640 12310
rect 10600 9172 10652 9178
rect 10600 9114 10652 9120
rect 10232 9104 10284 9110
rect 10232 9046 10284 9052
rect 10598 9072 10654 9081
rect 10598 9007 10654 9016
rect 10612 8974 10640 9007
rect 10600 8968 10652 8974
rect 10600 8910 10652 8916
rect 10508 8832 10560 8838
rect 10508 8774 10560 8780
rect 10600 8832 10652 8838
rect 10600 8774 10652 8780
rect 10520 8498 10548 8774
rect 10612 8634 10640 8774
rect 10600 8628 10652 8634
rect 10600 8570 10652 8576
rect 10508 8492 10560 8498
rect 10508 8434 10560 8440
rect 10704 7886 10732 12406
rect 10796 8634 10824 14350
rect 11060 14000 11112 14006
rect 11060 13942 11112 13948
rect 10968 13932 11020 13938
rect 10968 13874 11020 13880
rect 10876 10600 10928 10606
rect 10876 10542 10928 10548
rect 10784 8628 10836 8634
rect 10784 8570 10836 8576
rect 10416 7880 10468 7886
rect 10416 7822 10468 7828
rect 10508 7880 10560 7886
rect 10508 7822 10560 7828
rect 10692 7880 10744 7886
rect 10692 7822 10744 7828
rect 10324 7404 10376 7410
rect 10324 7346 10376 7352
rect 10336 6730 10364 7346
rect 10324 6724 10376 6730
rect 10324 6666 10376 6672
rect 10336 6458 10364 6666
rect 10324 6452 10376 6458
rect 10324 6394 10376 6400
rect 10232 6112 10284 6118
rect 10232 6054 10284 6060
rect 10244 5914 10272 6054
rect 10232 5908 10284 5914
rect 10232 5850 10284 5856
rect 10244 5778 10272 5850
rect 10232 5772 10284 5778
rect 10232 5714 10284 5720
rect 10232 4140 10284 4146
rect 10232 4082 10284 4088
rect 10140 3936 10192 3942
rect 10140 3878 10192 3884
rect 10138 3768 10194 3777
rect 10244 3738 10272 4082
rect 10138 3703 10194 3712
rect 10232 3732 10284 3738
rect 10048 3664 10100 3670
rect 10048 3606 10100 3612
rect 10152 3194 10180 3703
rect 10232 3674 10284 3680
rect 10428 3482 10456 7822
rect 10520 7478 10548 7822
rect 10508 7472 10560 7478
rect 10508 7414 10560 7420
rect 10508 7268 10560 7274
rect 10508 7210 10560 7216
rect 10520 4010 10548 7210
rect 10784 7200 10836 7206
rect 10784 7142 10836 7148
rect 10796 6905 10824 7142
rect 10782 6896 10838 6905
rect 10782 6831 10838 6840
rect 10796 6662 10824 6831
rect 10784 6656 10836 6662
rect 10784 6598 10836 6604
rect 10796 5030 10824 6598
rect 10784 5024 10836 5030
rect 10784 4966 10836 4972
rect 10784 4684 10836 4690
rect 10784 4626 10836 4632
rect 10796 4214 10824 4626
rect 10784 4208 10836 4214
rect 10784 4150 10836 4156
rect 10692 4072 10744 4078
rect 10598 4040 10654 4049
rect 10508 4004 10560 4010
rect 10692 4014 10744 4020
rect 10598 3975 10654 3984
rect 10508 3946 10560 3952
rect 10612 3942 10640 3975
rect 10600 3936 10652 3942
rect 10600 3878 10652 3884
rect 10428 3454 10640 3482
rect 10416 3392 10468 3398
rect 10416 3334 10468 3340
rect 10508 3392 10560 3398
rect 10508 3334 10560 3340
rect 10428 3194 10456 3334
rect 10520 3194 10548 3334
rect 10140 3188 10192 3194
rect 10140 3130 10192 3136
rect 10416 3188 10468 3194
rect 10416 3130 10468 3136
rect 10508 3188 10560 3194
rect 10508 3130 10560 3136
rect 9956 3120 10008 3126
rect 10612 3074 10640 3454
rect 9956 3062 10008 3068
rect 10520 3046 10640 3074
rect 10140 2984 10192 2990
rect 10140 2926 10192 2932
rect 9680 2916 9732 2922
rect 9680 2858 9732 2864
rect 9692 2650 9720 2858
rect 9680 2644 9732 2650
rect 9680 2586 9732 2592
rect 9864 2440 9916 2446
rect 9864 2382 9916 2388
rect 9876 800 9904 2382
rect 10152 800 10180 2926
rect 10520 2650 10548 3046
rect 10600 2984 10652 2990
rect 10600 2926 10652 2932
rect 10508 2644 10560 2650
rect 10508 2586 10560 2592
rect 10612 1442 10640 2926
rect 10704 2564 10732 4014
rect 10796 3777 10824 4150
rect 10782 3768 10838 3777
rect 10888 3738 10916 10542
rect 10980 8090 11008 13874
rect 11072 13394 11100 13942
rect 11152 13728 11204 13734
rect 11152 13670 11204 13676
rect 11060 13388 11112 13394
rect 11060 13330 11112 13336
rect 11060 12844 11112 12850
rect 11164 12832 11192 13670
rect 11112 12804 11192 12832
rect 11060 12786 11112 12792
rect 11072 12238 11100 12786
rect 11256 12458 11284 14350
rect 11900 13870 11928 14350
rect 11888 13864 11940 13870
rect 11888 13806 11940 13812
rect 11369 13628 11677 13637
rect 11369 13626 11375 13628
rect 11431 13626 11455 13628
rect 11511 13626 11535 13628
rect 11591 13626 11615 13628
rect 11671 13626 11677 13628
rect 11431 13574 11433 13626
rect 11613 13574 11615 13626
rect 11369 13572 11375 13574
rect 11431 13572 11455 13574
rect 11511 13572 11535 13574
rect 11591 13572 11615 13574
rect 11671 13572 11677 13574
rect 11369 13563 11677 13572
rect 11428 13388 11480 13394
rect 11428 13330 11480 13336
rect 11440 12646 11468 13330
rect 11900 13326 11928 13806
rect 12164 13728 12216 13734
rect 12268 13716 12296 14894
rect 12360 14618 12388 15302
rect 13280 15162 13308 15438
rect 13268 15156 13320 15162
rect 13268 15098 13320 15104
rect 13740 15026 13768 17138
rect 13820 16992 13872 16998
rect 13820 16934 13872 16940
rect 13832 16794 13860 16934
rect 13820 16788 13872 16794
rect 13820 16730 13872 16736
rect 14292 15706 14320 26250
rect 14842 26140 15150 26149
rect 14842 26138 14848 26140
rect 14904 26138 14928 26140
rect 14984 26138 15008 26140
rect 15064 26138 15088 26140
rect 15144 26138 15150 26140
rect 14904 26086 14906 26138
rect 15086 26086 15088 26138
rect 14842 26084 14848 26086
rect 14904 26084 14928 26086
rect 14984 26084 15008 26086
rect 15064 26084 15088 26086
rect 15144 26084 15150 26086
rect 14842 26075 15150 26084
rect 21788 26140 22096 26149
rect 21788 26138 21794 26140
rect 21850 26138 21874 26140
rect 21930 26138 21954 26140
rect 22010 26138 22034 26140
rect 22090 26138 22096 26140
rect 21850 26086 21852 26138
rect 22032 26086 22034 26138
rect 21788 26084 21794 26086
rect 21850 26084 21874 26086
rect 21930 26084 21954 26086
rect 22010 26084 22034 26086
rect 22090 26084 22096 26086
rect 21788 26075 22096 26084
rect 18315 25596 18623 25605
rect 18315 25594 18321 25596
rect 18377 25594 18401 25596
rect 18457 25594 18481 25596
rect 18537 25594 18561 25596
rect 18617 25594 18623 25596
rect 18377 25542 18379 25594
rect 18559 25542 18561 25594
rect 18315 25540 18321 25542
rect 18377 25540 18401 25542
rect 18457 25540 18481 25542
rect 18537 25540 18561 25542
rect 18617 25540 18623 25542
rect 18315 25531 18623 25540
rect 14842 25052 15150 25061
rect 14842 25050 14848 25052
rect 14904 25050 14928 25052
rect 14984 25050 15008 25052
rect 15064 25050 15088 25052
rect 15144 25050 15150 25052
rect 14904 24998 14906 25050
rect 15086 24998 15088 25050
rect 14842 24996 14848 24998
rect 14904 24996 14928 24998
rect 14984 24996 15008 24998
rect 15064 24996 15088 24998
rect 15144 24996 15150 24998
rect 14842 24987 15150 24996
rect 21788 25052 22096 25061
rect 21788 25050 21794 25052
rect 21850 25050 21874 25052
rect 21930 25050 21954 25052
rect 22010 25050 22034 25052
rect 22090 25050 22096 25052
rect 21850 24998 21852 25050
rect 22032 24998 22034 25050
rect 21788 24996 21794 24998
rect 21850 24996 21874 24998
rect 21930 24996 21954 24998
rect 22010 24996 22034 24998
rect 22090 24996 22096 24998
rect 21788 24987 22096 24996
rect 18315 24508 18623 24517
rect 18315 24506 18321 24508
rect 18377 24506 18401 24508
rect 18457 24506 18481 24508
rect 18537 24506 18561 24508
rect 18617 24506 18623 24508
rect 18377 24454 18379 24506
rect 18559 24454 18561 24506
rect 18315 24452 18321 24454
rect 18377 24452 18401 24454
rect 18457 24452 18481 24454
rect 18537 24452 18561 24454
rect 18617 24452 18623 24454
rect 18315 24443 18623 24452
rect 14842 23964 15150 23973
rect 14842 23962 14848 23964
rect 14904 23962 14928 23964
rect 14984 23962 15008 23964
rect 15064 23962 15088 23964
rect 15144 23962 15150 23964
rect 14904 23910 14906 23962
rect 15086 23910 15088 23962
rect 14842 23908 14848 23910
rect 14904 23908 14928 23910
rect 14984 23908 15008 23910
rect 15064 23908 15088 23910
rect 15144 23908 15150 23910
rect 14842 23899 15150 23908
rect 21788 23964 22096 23973
rect 21788 23962 21794 23964
rect 21850 23962 21874 23964
rect 21930 23962 21954 23964
rect 22010 23962 22034 23964
rect 22090 23962 22096 23964
rect 21850 23910 21852 23962
rect 22032 23910 22034 23962
rect 21788 23908 21794 23910
rect 21850 23908 21874 23910
rect 21930 23908 21954 23910
rect 22010 23908 22034 23910
rect 22090 23908 22096 23910
rect 21788 23899 22096 23908
rect 18315 23420 18623 23429
rect 18315 23418 18321 23420
rect 18377 23418 18401 23420
rect 18457 23418 18481 23420
rect 18537 23418 18561 23420
rect 18617 23418 18623 23420
rect 18377 23366 18379 23418
rect 18559 23366 18561 23418
rect 18315 23364 18321 23366
rect 18377 23364 18401 23366
rect 18457 23364 18481 23366
rect 18537 23364 18561 23366
rect 18617 23364 18623 23366
rect 18315 23355 18623 23364
rect 16028 22976 16080 22982
rect 16028 22918 16080 22924
rect 14842 22876 15150 22885
rect 14842 22874 14848 22876
rect 14904 22874 14928 22876
rect 14984 22874 15008 22876
rect 15064 22874 15088 22876
rect 15144 22874 15150 22876
rect 14904 22822 14906 22874
rect 15086 22822 15088 22874
rect 14842 22820 14848 22822
rect 14904 22820 14928 22822
rect 14984 22820 15008 22822
rect 15064 22820 15088 22822
rect 15144 22820 15150 22822
rect 14842 22811 15150 22820
rect 14648 21888 14700 21894
rect 14648 21830 14700 21836
rect 14660 16590 14688 21830
rect 14842 21788 15150 21797
rect 14842 21786 14848 21788
rect 14904 21786 14928 21788
rect 14984 21786 15008 21788
rect 15064 21786 15088 21788
rect 15144 21786 15150 21788
rect 14904 21734 14906 21786
rect 15086 21734 15088 21786
rect 14842 21732 14848 21734
rect 14904 21732 14928 21734
rect 14984 21732 15008 21734
rect 15064 21732 15088 21734
rect 15144 21732 15150 21734
rect 14842 21723 15150 21732
rect 15752 21548 15804 21554
rect 15752 21490 15804 21496
rect 14842 20700 15150 20709
rect 14842 20698 14848 20700
rect 14904 20698 14928 20700
rect 14984 20698 15008 20700
rect 15064 20698 15088 20700
rect 15144 20698 15150 20700
rect 14904 20646 14906 20698
rect 15086 20646 15088 20698
rect 14842 20644 14848 20646
rect 14904 20644 14928 20646
rect 14984 20644 15008 20646
rect 15064 20644 15088 20646
rect 15144 20644 15150 20646
rect 14842 20635 15150 20644
rect 14842 19612 15150 19621
rect 14842 19610 14848 19612
rect 14904 19610 14928 19612
rect 14984 19610 15008 19612
rect 15064 19610 15088 19612
rect 15144 19610 15150 19612
rect 14904 19558 14906 19610
rect 15086 19558 15088 19610
rect 14842 19556 14848 19558
rect 14904 19556 14928 19558
rect 14984 19556 15008 19558
rect 15064 19556 15088 19558
rect 15144 19556 15150 19558
rect 14842 19547 15150 19556
rect 14842 18524 15150 18533
rect 14842 18522 14848 18524
rect 14904 18522 14928 18524
rect 14984 18522 15008 18524
rect 15064 18522 15088 18524
rect 15144 18522 15150 18524
rect 14904 18470 14906 18522
rect 15086 18470 15088 18522
rect 14842 18468 14848 18470
rect 14904 18468 14928 18470
rect 14984 18468 15008 18470
rect 15064 18468 15088 18470
rect 15144 18468 15150 18470
rect 14842 18459 15150 18468
rect 14842 17436 15150 17445
rect 14842 17434 14848 17436
rect 14904 17434 14928 17436
rect 14984 17434 15008 17436
rect 15064 17434 15088 17436
rect 15144 17434 15150 17436
rect 14904 17382 14906 17434
rect 15086 17382 15088 17434
rect 14842 17380 14848 17382
rect 14904 17380 14928 17382
rect 14984 17380 15008 17382
rect 15064 17380 15088 17382
rect 15144 17380 15150 17382
rect 14842 17371 15150 17380
rect 14740 17196 14792 17202
rect 14740 17138 14792 17144
rect 14648 16584 14700 16590
rect 14648 16526 14700 16532
rect 14280 15700 14332 15706
rect 14280 15642 14332 15648
rect 14292 15162 14320 15642
rect 14280 15156 14332 15162
rect 14280 15098 14332 15104
rect 13728 15020 13780 15026
rect 13728 14962 13780 14968
rect 13544 14884 13596 14890
rect 13544 14826 13596 14832
rect 12348 14612 12400 14618
rect 12348 14554 12400 14560
rect 13176 14408 13228 14414
rect 13176 14350 13228 14356
rect 12348 14272 12400 14278
rect 12348 14214 12400 14220
rect 12440 14272 12492 14278
rect 12440 14214 12492 14220
rect 12360 13870 12388 14214
rect 12452 14006 12480 14214
rect 13188 14074 13216 14350
rect 13556 14346 13584 14826
rect 13728 14816 13780 14822
rect 13728 14758 13780 14764
rect 14188 14816 14240 14822
rect 14188 14758 14240 14764
rect 13740 14618 13768 14758
rect 13728 14612 13780 14618
rect 13728 14554 13780 14560
rect 14200 14550 14228 14758
rect 14188 14544 14240 14550
rect 14188 14486 14240 14492
rect 13726 14376 13782 14385
rect 13544 14340 13596 14346
rect 13726 14311 13782 14320
rect 13544 14282 13596 14288
rect 12532 14068 12584 14074
rect 12532 14010 12584 14016
rect 13176 14068 13228 14074
rect 13176 14010 13228 14016
rect 12440 14000 12492 14006
rect 12440 13942 12492 13948
rect 12348 13864 12400 13870
rect 12348 13806 12400 13812
rect 12216 13688 12296 13716
rect 12440 13728 12492 13734
rect 12164 13670 12216 13676
rect 12440 13670 12492 13676
rect 11888 13320 11940 13326
rect 11888 13262 11940 13268
rect 11428 12640 11480 12646
rect 11428 12582 11480 12588
rect 11369 12540 11677 12549
rect 11369 12538 11375 12540
rect 11431 12538 11455 12540
rect 11511 12538 11535 12540
rect 11591 12538 11615 12540
rect 11671 12538 11677 12540
rect 11431 12486 11433 12538
rect 11613 12486 11615 12538
rect 11369 12484 11375 12486
rect 11431 12484 11455 12486
rect 11511 12484 11535 12486
rect 11591 12484 11615 12486
rect 11671 12484 11677 12486
rect 11369 12475 11677 12484
rect 11164 12430 11284 12458
rect 11060 12232 11112 12238
rect 11060 12174 11112 12180
rect 11072 11762 11100 12174
rect 11060 11756 11112 11762
rect 11060 11698 11112 11704
rect 11060 9920 11112 9926
rect 11060 9862 11112 9868
rect 11072 8974 11100 9862
rect 11060 8968 11112 8974
rect 11060 8910 11112 8916
rect 11164 8634 11192 12430
rect 11796 12368 11848 12374
rect 11796 12310 11848 12316
rect 11520 12300 11572 12306
rect 11520 12242 11572 12248
rect 11428 12232 11480 12238
rect 11428 12174 11480 12180
rect 11244 12096 11296 12102
rect 11244 12038 11296 12044
rect 11256 11150 11284 12038
rect 11440 11694 11468 12174
rect 11532 11898 11560 12242
rect 11520 11892 11572 11898
rect 11520 11834 11572 11840
rect 11428 11688 11480 11694
rect 11428 11630 11480 11636
rect 11704 11552 11756 11558
rect 11808 11540 11836 12310
rect 11900 11744 11928 13262
rect 12164 13252 12216 13258
rect 12164 13194 12216 13200
rect 12176 12986 12204 13194
rect 12164 12980 12216 12986
rect 12164 12922 12216 12928
rect 12452 12782 12480 13670
rect 12544 12782 12572 14010
rect 13740 13394 13768 14311
rect 14188 14272 14240 14278
rect 14188 14214 14240 14220
rect 14200 14006 14228 14214
rect 14188 14000 14240 14006
rect 14188 13942 14240 13948
rect 14292 13870 14320 15098
rect 14280 13864 14332 13870
rect 14280 13806 14332 13812
rect 13728 13388 13780 13394
rect 13728 13330 13780 13336
rect 13452 13252 13504 13258
rect 13452 13194 13504 13200
rect 12900 13184 12952 13190
rect 12900 13126 12952 13132
rect 12912 12782 12940 13126
rect 13464 12986 13492 13194
rect 13452 12980 13504 12986
rect 13452 12922 13504 12928
rect 14660 12918 14688 16526
rect 14752 15162 14780 17138
rect 14842 16348 15150 16357
rect 14842 16346 14848 16348
rect 14904 16346 14928 16348
rect 14984 16346 15008 16348
rect 15064 16346 15088 16348
rect 15144 16346 15150 16348
rect 14904 16294 14906 16346
rect 15086 16294 15088 16346
rect 14842 16292 14848 16294
rect 14904 16292 14928 16294
rect 14984 16292 15008 16294
rect 15064 16292 15088 16294
rect 15144 16292 15150 16294
rect 14842 16283 15150 16292
rect 15764 16182 15792 21490
rect 16040 17746 16068 22918
rect 21788 22876 22096 22885
rect 21788 22874 21794 22876
rect 21850 22874 21874 22876
rect 21930 22874 21954 22876
rect 22010 22874 22034 22876
rect 22090 22874 22096 22876
rect 21850 22822 21852 22874
rect 22032 22822 22034 22874
rect 21788 22820 21794 22822
rect 21850 22820 21874 22822
rect 21930 22820 21954 22822
rect 22010 22820 22034 22822
rect 22090 22820 22096 22822
rect 21788 22811 22096 22820
rect 18315 22332 18623 22341
rect 18315 22330 18321 22332
rect 18377 22330 18401 22332
rect 18457 22330 18481 22332
rect 18537 22330 18561 22332
rect 18617 22330 18623 22332
rect 18377 22278 18379 22330
rect 18559 22278 18561 22330
rect 18315 22276 18321 22278
rect 18377 22276 18401 22278
rect 18457 22276 18481 22278
rect 18537 22276 18561 22278
rect 18617 22276 18623 22278
rect 18315 22267 18623 22276
rect 21788 21788 22096 21797
rect 21788 21786 21794 21788
rect 21850 21786 21874 21788
rect 21930 21786 21954 21788
rect 22010 21786 22034 21788
rect 22090 21786 22096 21788
rect 21850 21734 21852 21786
rect 22032 21734 22034 21786
rect 21788 21732 21794 21734
rect 21850 21732 21874 21734
rect 21930 21732 21954 21734
rect 22010 21732 22034 21734
rect 22090 21732 22096 21734
rect 21788 21723 22096 21732
rect 18315 21244 18623 21253
rect 18315 21242 18321 21244
rect 18377 21242 18401 21244
rect 18457 21242 18481 21244
rect 18537 21242 18561 21244
rect 18617 21242 18623 21244
rect 18377 21190 18379 21242
rect 18559 21190 18561 21242
rect 18315 21188 18321 21190
rect 18377 21188 18401 21190
rect 18457 21188 18481 21190
rect 18537 21188 18561 21190
rect 18617 21188 18623 21190
rect 18315 21179 18623 21188
rect 21788 20700 22096 20709
rect 21788 20698 21794 20700
rect 21850 20698 21874 20700
rect 21930 20698 21954 20700
rect 22010 20698 22034 20700
rect 22090 20698 22096 20700
rect 21850 20646 21852 20698
rect 22032 20646 22034 20698
rect 21788 20644 21794 20646
rect 21850 20644 21874 20646
rect 21930 20644 21954 20646
rect 22010 20644 22034 20646
rect 22090 20644 22096 20646
rect 21788 20635 22096 20644
rect 16212 20256 16264 20262
rect 16212 20198 16264 20204
rect 16028 17740 16080 17746
rect 16028 17682 16080 17688
rect 15200 16176 15252 16182
rect 15200 16118 15252 16124
rect 15752 16176 15804 16182
rect 15752 16118 15804 16124
rect 14842 15260 15150 15269
rect 14842 15258 14848 15260
rect 14904 15258 14928 15260
rect 14984 15258 15008 15260
rect 15064 15258 15088 15260
rect 15144 15258 15150 15260
rect 14904 15206 14906 15258
rect 15086 15206 15088 15258
rect 14842 15204 14848 15206
rect 14904 15204 14928 15206
rect 14984 15204 15008 15206
rect 15064 15204 15088 15206
rect 15144 15204 15150 15206
rect 14842 15195 15150 15204
rect 14740 15156 14792 15162
rect 14740 15098 14792 15104
rect 14752 15026 14780 15098
rect 14740 15020 14792 15026
rect 14740 14962 14792 14968
rect 14752 14482 14780 14962
rect 14740 14476 14792 14482
rect 14740 14418 14792 14424
rect 14752 14006 14780 14418
rect 14842 14172 15150 14181
rect 14842 14170 14848 14172
rect 14904 14170 14928 14172
rect 14984 14170 15008 14172
rect 15064 14170 15088 14172
rect 15144 14170 15150 14172
rect 14904 14118 14906 14170
rect 15086 14118 15088 14170
rect 14842 14116 14848 14118
rect 14904 14116 14928 14118
rect 14984 14116 15008 14118
rect 15064 14116 15088 14118
rect 15144 14116 15150 14118
rect 14842 14107 15150 14116
rect 14740 14000 14792 14006
rect 14740 13942 14792 13948
rect 14752 12986 14780 13942
rect 14842 13084 15150 13093
rect 14842 13082 14848 13084
rect 14904 13082 14928 13084
rect 14984 13082 15008 13084
rect 15064 13082 15088 13084
rect 15144 13082 15150 13084
rect 14904 13030 14906 13082
rect 15086 13030 15088 13082
rect 14842 13028 14848 13030
rect 14904 13028 14928 13030
rect 14984 13028 15008 13030
rect 15064 13028 15088 13030
rect 15144 13028 15150 13030
rect 14842 13019 15150 13028
rect 14740 12980 14792 12986
rect 14740 12922 14792 12928
rect 14648 12912 14700 12918
rect 14648 12854 14700 12860
rect 13820 12844 13872 12850
rect 13820 12786 13872 12792
rect 12440 12776 12492 12782
rect 12440 12718 12492 12724
rect 12532 12776 12584 12782
rect 12532 12718 12584 12724
rect 12900 12776 12952 12782
rect 12900 12718 12952 12724
rect 13726 12744 13782 12753
rect 12452 12306 12480 12718
rect 13726 12679 13782 12688
rect 12348 12300 12400 12306
rect 12348 12242 12400 12248
rect 12440 12300 12492 12306
rect 12440 12242 12492 12248
rect 11980 11756 12032 11762
rect 11900 11716 11980 11744
rect 11980 11698 12032 11704
rect 11888 11620 11940 11626
rect 11888 11562 11940 11568
rect 11756 11512 11836 11540
rect 11704 11494 11756 11500
rect 11369 11452 11677 11461
rect 11369 11450 11375 11452
rect 11431 11450 11455 11452
rect 11511 11450 11535 11452
rect 11591 11450 11615 11452
rect 11671 11450 11677 11452
rect 11431 11398 11433 11450
rect 11613 11398 11615 11450
rect 11369 11396 11375 11398
rect 11431 11396 11455 11398
rect 11511 11396 11535 11398
rect 11591 11396 11615 11398
rect 11671 11396 11677 11398
rect 11369 11387 11677 11396
rect 11518 11248 11574 11257
rect 11518 11183 11574 11192
rect 11532 11150 11560 11183
rect 11244 11144 11296 11150
rect 11244 11086 11296 11092
rect 11520 11144 11572 11150
rect 11520 11086 11572 11092
rect 11532 10606 11560 11086
rect 11520 10600 11572 10606
rect 11520 10542 11572 10548
rect 11369 10364 11677 10373
rect 11369 10362 11375 10364
rect 11431 10362 11455 10364
rect 11511 10362 11535 10364
rect 11591 10362 11615 10364
rect 11671 10362 11677 10364
rect 11431 10310 11433 10362
rect 11613 10310 11615 10362
rect 11369 10308 11375 10310
rect 11431 10308 11455 10310
rect 11511 10308 11535 10310
rect 11591 10308 11615 10310
rect 11671 10308 11677 10310
rect 11369 10299 11677 10308
rect 11520 9988 11572 9994
rect 11520 9930 11572 9936
rect 11532 9674 11560 9930
rect 11440 9646 11560 9674
rect 11440 9450 11468 9646
rect 11716 9586 11744 11494
rect 11900 11082 11928 11562
rect 11992 11257 12020 11698
rect 12360 11694 12388 12242
rect 12452 12102 12480 12242
rect 13740 12170 13768 12679
rect 13728 12164 13780 12170
rect 13728 12106 13780 12112
rect 12440 12096 12492 12102
rect 12440 12038 12492 12044
rect 12992 12096 13044 12102
rect 12992 12038 13044 12044
rect 13084 12096 13136 12102
rect 13084 12038 13136 12044
rect 13636 12096 13688 12102
rect 13688 12044 13768 12050
rect 13636 12038 13768 12044
rect 13004 11778 13032 12038
rect 13096 11898 13124 12038
rect 13648 12022 13768 12038
rect 13084 11892 13136 11898
rect 13084 11834 13136 11840
rect 13004 11750 13124 11778
rect 13740 11762 13768 12022
rect 12348 11688 12400 11694
rect 12348 11630 12400 11636
rect 12256 11552 12308 11558
rect 12256 11494 12308 11500
rect 11978 11248 12034 11257
rect 11978 11183 12034 11192
rect 12268 11082 12296 11494
rect 11888 11076 11940 11082
rect 11888 11018 11940 11024
rect 12256 11076 12308 11082
rect 12256 11018 12308 11024
rect 11796 10600 11848 10606
rect 11796 10542 11848 10548
rect 11808 10266 11836 10542
rect 11796 10260 11848 10266
rect 11796 10202 11848 10208
rect 12072 10192 12124 10198
rect 12072 10134 12124 10140
rect 12084 9654 12112 10134
rect 12360 10062 12388 11630
rect 12440 11348 12492 11354
rect 12440 11290 12492 11296
rect 12452 10130 12480 11290
rect 13096 11150 13124 11750
rect 13728 11756 13780 11762
rect 13728 11698 13780 11704
rect 13544 11688 13596 11694
rect 13544 11630 13596 11636
rect 13084 11144 13136 11150
rect 13084 11086 13136 11092
rect 13556 11014 13584 11630
rect 13544 11008 13596 11014
rect 13544 10950 13596 10956
rect 13556 10742 13584 10950
rect 12808 10736 12860 10742
rect 12808 10678 12860 10684
rect 13544 10736 13596 10742
rect 13544 10678 13596 10684
rect 12820 10266 12848 10678
rect 12808 10260 12860 10266
rect 12808 10202 12860 10208
rect 12440 10124 12492 10130
rect 12440 10066 12492 10072
rect 12348 10056 12400 10062
rect 12348 9998 12400 10004
rect 12072 9648 12124 9654
rect 12072 9590 12124 9596
rect 11704 9580 11756 9586
rect 11704 9522 11756 9528
rect 11428 9444 11480 9450
rect 11428 9386 11480 9392
rect 11244 9376 11296 9382
rect 11244 9318 11296 9324
rect 11256 9160 11284 9318
rect 11369 9276 11677 9285
rect 11369 9274 11375 9276
rect 11431 9274 11455 9276
rect 11511 9274 11535 9276
rect 11591 9274 11615 9276
rect 11671 9274 11677 9276
rect 11431 9222 11433 9274
rect 11613 9222 11615 9274
rect 11369 9220 11375 9222
rect 11431 9220 11455 9222
rect 11511 9220 11535 9222
rect 11591 9220 11615 9222
rect 11671 9220 11677 9222
rect 11369 9211 11677 9220
rect 11716 9160 11744 9522
rect 11796 9376 11848 9382
rect 11796 9318 11848 9324
rect 11256 9132 11744 9160
rect 11152 8628 11204 8634
rect 11152 8570 11204 8576
rect 11256 8514 11284 9132
rect 11164 8486 11284 8514
rect 11060 8424 11112 8430
rect 11060 8366 11112 8372
rect 10968 8084 11020 8090
rect 10968 8026 11020 8032
rect 10968 5160 11020 5166
rect 10968 5102 11020 5108
rect 10980 3738 11008 5102
rect 10782 3703 10838 3712
rect 10876 3732 10928 3738
rect 10876 3674 10928 3680
rect 10968 3732 11020 3738
rect 10968 3674 11020 3680
rect 10968 3528 11020 3534
rect 10968 3470 11020 3476
rect 10784 3392 10836 3398
rect 10784 3334 10836 3340
rect 10796 3058 10824 3334
rect 10784 3052 10836 3058
rect 10784 2994 10836 3000
rect 10980 2666 11008 3470
rect 11072 3398 11100 8366
rect 11164 7206 11192 8486
rect 11244 8424 11296 8430
rect 11244 8366 11296 8372
rect 11152 7200 11204 7206
rect 11152 7142 11204 7148
rect 11152 5024 11204 5030
rect 11152 4966 11204 4972
rect 11164 4486 11192 4966
rect 11152 4480 11204 4486
rect 11152 4422 11204 4428
rect 11152 3460 11204 3466
rect 11152 3402 11204 3408
rect 11060 3392 11112 3398
rect 11060 3334 11112 3340
rect 10980 2638 11100 2666
rect 10968 2576 11020 2582
rect 10704 2536 10916 2564
rect 10692 2440 10744 2446
rect 10692 2382 10744 2388
rect 10784 2440 10836 2446
rect 10784 2382 10836 2388
rect 10428 1414 10640 1442
rect 10428 800 10456 1414
rect 10704 800 10732 2382
rect 10796 1306 10824 2382
rect 10888 2038 10916 2536
rect 10968 2518 11020 2524
rect 10876 2032 10928 2038
rect 10876 1974 10928 1980
rect 10980 1766 11008 2518
rect 11072 2446 11100 2638
rect 11060 2440 11112 2446
rect 11060 2382 11112 2388
rect 10968 1760 11020 1766
rect 10968 1702 11020 1708
rect 11164 1562 11192 3402
rect 11256 3194 11284 8366
rect 11369 8188 11677 8197
rect 11369 8186 11375 8188
rect 11431 8186 11455 8188
rect 11511 8186 11535 8188
rect 11591 8186 11615 8188
rect 11671 8186 11677 8188
rect 11431 8134 11433 8186
rect 11613 8134 11615 8186
rect 11369 8132 11375 8134
rect 11431 8132 11455 8134
rect 11511 8132 11535 8134
rect 11591 8132 11615 8134
rect 11671 8132 11677 8134
rect 11369 8123 11677 8132
rect 11808 7410 11836 9318
rect 12084 9042 12112 9590
rect 13556 9450 13584 10678
rect 13740 10674 13768 11698
rect 13728 10668 13780 10674
rect 13728 10610 13780 10616
rect 13544 9444 13596 9450
rect 13544 9386 13596 9392
rect 13832 9382 13860 12786
rect 15212 12442 15240 16118
rect 15292 14952 15344 14958
rect 15292 14894 15344 14900
rect 15304 13870 15332 14894
rect 15476 14816 15528 14822
rect 15476 14758 15528 14764
rect 15752 14816 15804 14822
rect 15752 14758 15804 14764
rect 15936 14816 15988 14822
rect 15936 14758 15988 14764
rect 15488 13938 15516 14758
rect 15764 14414 15792 14758
rect 15752 14408 15804 14414
rect 15752 14350 15804 14356
rect 15476 13932 15528 13938
rect 15476 13874 15528 13880
rect 15292 13864 15344 13870
rect 15292 13806 15344 13812
rect 15290 13424 15346 13433
rect 15290 13359 15346 13368
rect 15304 12850 15332 13359
rect 15752 13320 15804 13326
rect 15750 13288 15752 13297
rect 15804 13288 15806 13297
rect 15750 13223 15806 13232
rect 15844 13184 15896 13190
rect 15844 13126 15896 13132
rect 15292 12844 15344 12850
rect 15292 12786 15344 12792
rect 15476 12640 15528 12646
rect 15476 12582 15528 12588
rect 15200 12436 15252 12442
rect 15200 12378 15252 12384
rect 14188 12096 14240 12102
rect 14188 12038 14240 12044
rect 14200 11830 14228 12038
rect 14842 11996 15150 12005
rect 14842 11994 14848 11996
rect 14904 11994 14928 11996
rect 14984 11994 15008 11996
rect 15064 11994 15088 11996
rect 15144 11994 15150 11996
rect 14904 11942 14906 11994
rect 15086 11942 15088 11994
rect 14842 11940 14848 11942
rect 14904 11940 14928 11942
rect 14984 11940 15008 11942
rect 15064 11940 15088 11942
rect 15144 11940 15150 11942
rect 14842 11931 15150 11940
rect 14188 11824 14240 11830
rect 14188 11766 14240 11772
rect 14464 11076 14516 11082
rect 14464 11018 14516 11024
rect 14004 10464 14056 10470
rect 14004 10406 14056 10412
rect 13820 9376 13872 9382
rect 13820 9318 13872 9324
rect 12072 9036 12124 9042
rect 12072 8978 12124 8984
rect 12440 8832 12492 8838
rect 12440 8774 12492 8780
rect 12164 8424 12216 8430
rect 12164 8366 12216 8372
rect 11796 7404 11848 7410
rect 11796 7346 11848 7352
rect 11369 7100 11677 7109
rect 11369 7098 11375 7100
rect 11431 7098 11455 7100
rect 11511 7098 11535 7100
rect 11591 7098 11615 7100
rect 11671 7098 11677 7100
rect 11431 7046 11433 7098
rect 11613 7046 11615 7098
rect 11369 7044 11375 7046
rect 11431 7044 11455 7046
rect 11511 7044 11535 7046
rect 11591 7044 11615 7046
rect 11671 7044 11677 7046
rect 11369 7035 11677 7044
rect 11980 6928 12032 6934
rect 11980 6870 12032 6876
rect 11369 6012 11677 6021
rect 11369 6010 11375 6012
rect 11431 6010 11455 6012
rect 11511 6010 11535 6012
rect 11591 6010 11615 6012
rect 11671 6010 11677 6012
rect 11431 5958 11433 6010
rect 11613 5958 11615 6010
rect 11369 5956 11375 5958
rect 11431 5956 11455 5958
rect 11511 5956 11535 5958
rect 11591 5956 11615 5958
rect 11671 5956 11677 5958
rect 11369 5947 11677 5956
rect 11704 5840 11756 5846
rect 11704 5782 11756 5788
rect 11369 4924 11677 4933
rect 11369 4922 11375 4924
rect 11431 4922 11455 4924
rect 11511 4922 11535 4924
rect 11591 4922 11615 4924
rect 11671 4922 11677 4924
rect 11431 4870 11433 4922
rect 11613 4870 11615 4922
rect 11369 4868 11375 4870
rect 11431 4868 11455 4870
rect 11511 4868 11535 4870
rect 11591 4868 11615 4870
rect 11671 4868 11677 4870
rect 11369 4859 11677 4868
rect 11334 4176 11390 4185
rect 11334 4111 11336 4120
rect 11388 4111 11390 4120
rect 11336 4082 11388 4088
rect 11369 3836 11677 3845
rect 11369 3834 11375 3836
rect 11431 3834 11455 3836
rect 11511 3834 11535 3836
rect 11591 3834 11615 3836
rect 11671 3834 11677 3836
rect 11431 3782 11433 3834
rect 11613 3782 11615 3834
rect 11369 3780 11375 3782
rect 11431 3780 11455 3782
rect 11511 3780 11535 3782
rect 11591 3780 11615 3782
rect 11671 3780 11677 3782
rect 11369 3771 11677 3780
rect 11336 3528 11388 3534
rect 11336 3470 11388 3476
rect 11244 3188 11296 3194
rect 11244 3130 11296 3136
rect 11348 2854 11376 3470
rect 11716 3176 11744 5782
rect 11796 5568 11848 5574
rect 11796 5510 11848 5516
rect 11808 3346 11836 5510
rect 11888 3936 11940 3942
rect 11888 3878 11940 3884
rect 11900 3738 11928 3878
rect 11888 3732 11940 3738
rect 11888 3674 11940 3680
rect 11808 3318 11928 3346
rect 11900 3194 11928 3318
rect 11992 3194 12020 6870
rect 12072 4480 12124 4486
rect 12072 4422 12124 4428
rect 12084 4010 12112 4422
rect 12072 4004 12124 4010
rect 12072 3946 12124 3952
rect 12084 3738 12112 3946
rect 12072 3732 12124 3738
rect 12072 3674 12124 3680
rect 11888 3188 11940 3194
rect 11716 3148 11836 3176
rect 11704 3052 11756 3058
rect 11704 2994 11756 3000
rect 11336 2848 11388 2854
rect 11336 2790 11388 2796
rect 11369 2748 11677 2757
rect 11369 2746 11375 2748
rect 11431 2746 11455 2748
rect 11511 2746 11535 2748
rect 11591 2746 11615 2748
rect 11671 2746 11677 2748
rect 11431 2694 11433 2746
rect 11613 2694 11615 2746
rect 11369 2692 11375 2694
rect 11431 2692 11455 2694
rect 11511 2692 11535 2694
rect 11591 2692 11615 2694
rect 11671 2692 11677 2694
rect 11369 2683 11677 2692
rect 11716 2650 11744 2994
rect 11808 2774 11836 3148
rect 11888 3130 11940 3136
rect 11980 3188 12032 3194
rect 11980 3130 12032 3136
rect 11808 2746 12020 2774
rect 11704 2644 11756 2650
rect 11704 2586 11756 2592
rect 11244 2440 11296 2446
rect 11244 2382 11296 2388
rect 11152 1556 11204 1562
rect 11152 1498 11204 1504
rect 10796 1278 11008 1306
rect 10980 800 11008 1278
rect 11256 800 11284 2382
rect 11992 2310 12020 2746
rect 12176 2650 12204 8366
rect 12256 8016 12308 8022
rect 12256 7958 12308 7964
rect 12268 7478 12296 7958
rect 12256 7472 12308 7478
rect 12256 7414 12308 7420
rect 12452 4826 12480 8774
rect 13176 8084 13228 8090
rect 13176 8026 13228 8032
rect 12532 7880 12584 7886
rect 12532 7822 12584 7828
rect 12440 4820 12492 4826
rect 12440 4762 12492 4768
rect 12348 4752 12400 4758
rect 12348 4694 12400 4700
rect 12254 3632 12310 3641
rect 12254 3567 12310 3576
rect 12268 3058 12296 3567
rect 12360 3194 12388 4694
rect 12348 3188 12400 3194
rect 12348 3130 12400 3136
rect 12256 3052 12308 3058
rect 12256 2994 12308 3000
rect 12544 2650 12572 7822
rect 13188 7449 13216 8026
rect 13174 7440 13230 7449
rect 13174 7375 13230 7384
rect 13266 7304 13322 7313
rect 13266 7239 13322 7248
rect 12624 6724 12676 6730
rect 12624 6666 12676 6672
rect 12636 4758 12664 6666
rect 13084 5568 13136 5574
rect 13084 5510 13136 5516
rect 12624 4752 12676 4758
rect 12624 4694 12676 4700
rect 12164 2644 12216 2650
rect 12164 2586 12216 2592
rect 12532 2644 12584 2650
rect 12532 2586 12584 2592
rect 13096 2582 13124 5510
rect 13084 2576 13136 2582
rect 13084 2518 13136 2524
rect 13280 2446 13308 7239
rect 14016 5778 14044 10406
rect 14186 9616 14242 9625
rect 14186 9551 14188 9560
rect 14240 9551 14242 9560
rect 14188 9522 14240 9528
rect 14004 5772 14056 5778
rect 14004 5714 14056 5720
rect 14476 5302 14504 11018
rect 14842 10908 15150 10917
rect 14842 10906 14848 10908
rect 14904 10906 14928 10908
rect 14984 10906 15008 10908
rect 15064 10906 15088 10908
rect 15144 10906 15150 10908
rect 14904 10854 14906 10906
rect 15086 10854 15088 10906
rect 14842 10852 14848 10854
rect 14904 10852 14928 10854
rect 14984 10852 15008 10854
rect 15064 10852 15088 10854
rect 15144 10852 15150 10854
rect 14842 10843 15150 10852
rect 14842 9820 15150 9829
rect 14842 9818 14848 9820
rect 14904 9818 14928 9820
rect 14984 9818 15008 9820
rect 15064 9818 15088 9820
rect 15144 9818 15150 9820
rect 14904 9766 14906 9818
rect 15086 9766 15088 9818
rect 14842 9764 14848 9766
rect 14904 9764 14928 9766
rect 14984 9764 15008 9766
rect 15064 9764 15088 9766
rect 15144 9764 15150 9766
rect 14842 9755 15150 9764
rect 14842 8732 15150 8741
rect 14842 8730 14848 8732
rect 14904 8730 14928 8732
rect 14984 8730 15008 8732
rect 15064 8730 15088 8732
rect 15144 8730 15150 8732
rect 14904 8678 14906 8730
rect 15086 8678 15088 8730
rect 14842 8676 14848 8678
rect 14904 8676 14928 8678
rect 14984 8676 15008 8678
rect 15064 8676 15088 8678
rect 15144 8676 15150 8678
rect 14842 8667 15150 8676
rect 15488 7886 15516 12582
rect 15566 12336 15622 12345
rect 15566 12271 15622 12280
rect 15580 12238 15608 12271
rect 15568 12232 15620 12238
rect 15568 12174 15620 12180
rect 15476 7880 15528 7886
rect 15476 7822 15528 7828
rect 14648 7812 14700 7818
rect 14648 7754 14700 7760
rect 14464 5296 14516 5302
rect 14464 5238 14516 5244
rect 13268 2440 13320 2446
rect 13268 2382 13320 2388
rect 11980 2304 12032 2310
rect 11980 2246 12032 2252
rect 13084 2304 13136 2310
rect 13084 2246 13136 2252
rect 13096 2106 13124 2246
rect 13084 2100 13136 2106
rect 13084 2042 13136 2048
rect 14660 1970 14688 7754
rect 14842 7644 15150 7653
rect 14842 7642 14848 7644
rect 14904 7642 14928 7644
rect 14984 7642 15008 7644
rect 15064 7642 15088 7644
rect 15144 7642 15150 7644
rect 14904 7590 14906 7642
rect 15086 7590 15088 7642
rect 14842 7588 14848 7590
rect 14904 7588 14928 7590
rect 14984 7588 15008 7590
rect 15064 7588 15088 7590
rect 15144 7588 15150 7590
rect 14842 7579 15150 7588
rect 14842 6556 15150 6565
rect 14842 6554 14848 6556
rect 14904 6554 14928 6556
rect 14984 6554 15008 6556
rect 15064 6554 15088 6556
rect 15144 6554 15150 6556
rect 14904 6502 14906 6554
rect 15086 6502 15088 6554
rect 14842 6500 14848 6502
rect 14904 6500 14928 6502
rect 14984 6500 15008 6502
rect 15064 6500 15088 6502
rect 15144 6500 15150 6502
rect 14842 6491 15150 6500
rect 14842 5468 15150 5477
rect 14842 5466 14848 5468
rect 14904 5466 14928 5468
rect 14984 5466 15008 5468
rect 15064 5466 15088 5468
rect 15144 5466 15150 5468
rect 14904 5414 14906 5466
rect 15086 5414 15088 5466
rect 14842 5412 14848 5414
rect 14904 5412 14928 5414
rect 14984 5412 15008 5414
rect 15064 5412 15088 5414
rect 15144 5412 15150 5414
rect 14842 5403 15150 5412
rect 14842 4380 15150 4389
rect 14842 4378 14848 4380
rect 14904 4378 14928 4380
rect 14984 4378 15008 4380
rect 15064 4378 15088 4380
rect 15144 4378 15150 4380
rect 14904 4326 14906 4378
rect 15086 4326 15088 4378
rect 14842 4324 14848 4326
rect 14904 4324 14928 4326
rect 14984 4324 15008 4326
rect 15064 4324 15088 4326
rect 15144 4324 15150 4326
rect 14842 4315 15150 4324
rect 15198 3496 15254 3505
rect 15198 3431 15254 3440
rect 14842 3292 15150 3301
rect 14842 3290 14848 3292
rect 14904 3290 14928 3292
rect 14984 3290 15008 3292
rect 15064 3290 15088 3292
rect 15144 3290 15150 3292
rect 14904 3238 14906 3290
rect 15086 3238 15088 3290
rect 14842 3236 14848 3238
rect 14904 3236 14928 3238
rect 14984 3236 15008 3238
rect 15064 3236 15088 3238
rect 15144 3236 15150 3238
rect 14842 3227 15150 3236
rect 15212 2310 15240 3431
rect 15856 3058 15884 13126
rect 15948 11801 15976 14758
rect 16040 13394 16068 17682
rect 16224 15434 16252 20198
rect 18315 20156 18623 20165
rect 18315 20154 18321 20156
rect 18377 20154 18401 20156
rect 18457 20154 18481 20156
rect 18537 20154 18561 20156
rect 18617 20154 18623 20156
rect 18377 20102 18379 20154
rect 18559 20102 18561 20154
rect 18315 20100 18321 20102
rect 18377 20100 18401 20102
rect 18457 20100 18481 20102
rect 18537 20100 18561 20102
rect 18617 20100 18623 20102
rect 18315 20091 18623 20100
rect 21788 19612 22096 19621
rect 21788 19610 21794 19612
rect 21850 19610 21874 19612
rect 21930 19610 21954 19612
rect 22010 19610 22034 19612
rect 22090 19610 22096 19612
rect 21850 19558 21852 19610
rect 22032 19558 22034 19610
rect 21788 19556 21794 19558
rect 21850 19556 21874 19558
rect 21930 19556 21954 19558
rect 22010 19556 22034 19558
rect 22090 19556 22096 19558
rect 21788 19547 22096 19556
rect 18315 19068 18623 19077
rect 18315 19066 18321 19068
rect 18377 19066 18401 19068
rect 18457 19066 18481 19068
rect 18537 19066 18561 19068
rect 18617 19066 18623 19068
rect 18377 19014 18379 19066
rect 18559 19014 18561 19066
rect 18315 19012 18321 19014
rect 18377 19012 18401 19014
rect 18457 19012 18481 19014
rect 18537 19012 18561 19014
rect 18617 19012 18623 19014
rect 18315 19003 18623 19012
rect 17776 18624 17828 18630
rect 17776 18566 17828 18572
rect 16580 17196 16632 17202
rect 16580 17138 16632 17144
rect 16212 15428 16264 15434
rect 16212 15370 16264 15376
rect 16118 13832 16174 13841
rect 16118 13767 16174 13776
rect 16028 13388 16080 13394
rect 16028 13330 16080 13336
rect 16132 12850 16160 13767
rect 16120 12844 16172 12850
rect 16120 12786 16172 12792
rect 16224 12442 16252 15370
rect 16304 14272 16356 14278
rect 16304 14214 16356 14220
rect 16212 12436 16264 12442
rect 16212 12378 16264 12384
rect 15934 11792 15990 11801
rect 15990 11750 16068 11778
rect 15934 11727 15990 11736
rect 16040 10742 16068 11750
rect 16028 10736 16080 10742
rect 16028 10678 16080 10684
rect 15936 10668 15988 10674
rect 15936 10610 15988 10616
rect 15948 10577 15976 10610
rect 15934 10568 15990 10577
rect 15934 10503 15990 10512
rect 16120 10464 16172 10470
rect 16120 10406 16172 10412
rect 16132 4690 16160 10406
rect 16316 7410 16344 14214
rect 16488 13864 16540 13870
rect 16488 13806 16540 13812
rect 16396 13184 16448 13190
rect 16396 13126 16448 13132
rect 16408 12986 16436 13126
rect 16396 12980 16448 12986
rect 16396 12922 16448 12928
rect 16304 7404 16356 7410
rect 16304 7346 16356 7352
rect 16120 4684 16172 4690
rect 16120 4626 16172 4632
rect 16500 4622 16528 13806
rect 16592 11218 16620 17138
rect 17684 14000 17736 14006
rect 17684 13942 17736 13948
rect 17224 12640 17276 12646
rect 17224 12582 17276 12588
rect 16672 12436 16724 12442
rect 17236 12434 17264 12582
rect 17236 12406 17448 12434
rect 16672 12378 16724 12384
rect 16684 11898 16712 12378
rect 17130 12200 17186 12209
rect 17130 12135 17186 12144
rect 16672 11892 16724 11898
rect 16672 11834 16724 11840
rect 17144 11762 17172 12135
rect 17132 11756 17184 11762
rect 17132 11698 17184 11704
rect 16580 11212 16632 11218
rect 16580 11154 16632 11160
rect 17132 10668 17184 10674
rect 17132 10610 17184 10616
rect 17144 10266 17172 10610
rect 17132 10260 17184 10266
rect 17132 10202 17184 10208
rect 17224 10260 17276 10266
rect 17224 10202 17276 10208
rect 17236 9722 17264 10202
rect 17224 9716 17276 9722
rect 17224 9658 17276 9664
rect 17224 9444 17276 9450
rect 17224 9386 17276 9392
rect 17236 8566 17264 9386
rect 17224 8560 17276 8566
rect 17224 8502 17276 8508
rect 17224 6112 17276 6118
rect 17224 6054 17276 6060
rect 17236 5914 17264 6054
rect 17224 5908 17276 5914
rect 17224 5850 17276 5856
rect 17420 5234 17448 12406
rect 17408 5228 17460 5234
rect 17408 5170 17460 5176
rect 16488 4616 16540 4622
rect 16488 4558 16540 4564
rect 15844 3052 15896 3058
rect 15844 2994 15896 3000
rect 17696 2446 17724 13942
rect 17788 12918 17816 18566
rect 21788 18524 22096 18533
rect 21788 18522 21794 18524
rect 21850 18522 21874 18524
rect 21930 18522 21954 18524
rect 22010 18522 22034 18524
rect 22090 18522 22096 18524
rect 21850 18470 21852 18522
rect 22032 18470 22034 18522
rect 21788 18468 21794 18470
rect 21850 18468 21874 18470
rect 21930 18468 21954 18470
rect 22010 18468 22034 18470
rect 22090 18468 22096 18470
rect 21788 18459 22096 18468
rect 18315 17980 18623 17989
rect 18315 17978 18321 17980
rect 18377 17978 18401 17980
rect 18457 17978 18481 17980
rect 18537 17978 18561 17980
rect 18617 17978 18623 17980
rect 18377 17926 18379 17978
rect 18559 17926 18561 17978
rect 18315 17924 18321 17926
rect 18377 17924 18401 17926
rect 18457 17924 18481 17926
rect 18537 17924 18561 17926
rect 18617 17924 18623 17926
rect 18315 17915 18623 17924
rect 21788 17436 22096 17445
rect 21788 17434 21794 17436
rect 21850 17434 21874 17436
rect 21930 17434 21954 17436
rect 22010 17434 22034 17436
rect 22090 17434 22096 17436
rect 21850 17382 21852 17434
rect 22032 17382 22034 17434
rect 21788 17380 21794 17382
rect 21850 17380 21874 17382
rect 21930 17380 21954 17382
rect 22010 17380 22034 17382
rect 22090 17380 22096 17382
rect 21788 17371 22096 17380
rect 18315 16892 18623 16901
rect 18315 16890 18321 16892
rect 18377 16890 18401 16892
rect 18457 16890 18481 16892
rect 18537 16890 18561 16892
rect 18617 16890 18623 16892
rect 18377 16838 18379 16890
rect 18559 16838 18561 16890
rect 18315 16836 18321 16838
rect 18377 16836 18401 16838
rect 18457 16836 18481 16838
rect 18537 16836 18561 16838
rect 18617 16836 18623 16838
rect 18315 16827 18623 16836
rect 21788 16348 22096 16357
rect 21788 16346 21794 16348
rect 21850 16346 21874 16348
rect 21930 16346 21954 16348
rect 22010 16346 22034 16348
rect 22090 16346 22096 16348
rect 21850 16294 21852 16346
rect 22032 16294 22034 16346
rect 21788 16292 21794 16294
rect 21850 16292 21874 16294
rect 21930 16292 21954 16294
rect 22010 16292 22034 16294
rect 22090 16292 22096 16294
rect 21788 16283 22096 16292
rect 18315 15804 18623 15813
rect 18315 15802 18321 15804
rect 18377 15802 18401 15804
rect 18457 15802 18481 15804
rect 18537 15802 18561 15804
rect 18617 15802 18623 15804
rect 18377 15750 18379 15802
rect 18559 15750 18561 15802
rect 18315 15748 18321 15750
rect 18377 15748 18401 15750
rect 18457 15748 18481 15750
rect 18537 15748 18561 15750
rect 18617 15748 18623 15750
rect 18315 15739 18623 15748
rect 21788 15260 22096 15269
rect 21788 15258 21794 15260
rect 21850 15258 21874 15260
rect 21930 15258 21954 15260
rect 22010 15258 22034 15260
rect 22090 15258 22096 15260
rect 21850 15206 21852 15258
rect 22032 15206 22034 15258
rect 21788 15204 21794 15206
rect 21850 15204 21874 15206
rect 21930 15204 21954 15206
rect 22010 15204 22034 15206
rect 22090 15204 22096 15206
rect 21788 15195 22096 15204
rect 18315 14716 18623 14725
rect 18315 14714 18321 14716
rect 18377 14714 18401 14716
rect 18457 14714 18481 14716
rect 18537 14714 18561 14716
rect 18617 14714 18623 14716
rect 18377 14662 18379 14714
rect 18559 14662 18561 14714
rect 18315 14660 18321 14662
rect 18377 14660 18401 14662
rect 18457 14660 18481 14662
rect 18537 14660 18561 14662
rect 18617 14660 18623 14662
rect 18315 14651 18623 14660
rect 22756 14482 22784 26726
rect 25261 26684 25569 26693
rect 28354 26687 28410 26696
rect 25261 26682 25267 26684
rect 25323 26682 25347 26684
rect 25403 26682 25427 26684
rect 25483 26682 25507 26684
rect 25563 26682 25569 26684
rect 25323 26630 25325 26682
rect 25505 26630 25507 26682
rect 25261 26628 25267 26630
rect 25323 26628 25347 26630
rect 25403 26628 25427 26630
rect 25483 26628 25507 26630
rect 25563 26628 25569 26630
rect 25261 26619 25569 26628
rect 28356 26308 28408 26314
rect 28356 26250 28408 26256
rect 28368 25945 28396 26250
rect 28734 26140 29042 26149
rect 28734 26138 28740 26140
rect 28796 26138 28820 26140
rect 28876 26138 28900 26140
rect 28956 26138 28980 26140
rect 29036 26138 29042 26140
rect 28796 26086 28798 26138
rect 28978 26086 28980 26138
rect 28734 26084 28740 26086
rect 28796 26084 28820 26086
rect 28876 26084 28900 26086
rect 28956 26084 28980 26086
rect 29036 26084 29042 26086
rect 28734 26075 29042 26084
rect 28354 25936 28410 25945
rect 28354 25871 28410 25880
rect 25261 25596 25569 25605
rect 25261 25594 25267 25596
rect 25323 25594 25347 25596
rect 25403 25594 25427 25596
rect 25483 25594 25507 25596
rect 25563 25594 25569 25596
rect 25323 25542 25325 25594
rect 25505 25542 25507 25594
rect 25261 25540 25267 25542
rect 25323 25540 25347 25542
rect 25403 25540 25427 25542
rect 25483 25540 25507 25542
rect 25563 25540 25569 25542
rect 25261 25531 25569 25540
rect 28356 25220 28408 25226
rect 28356 25162 28408 25168
rect 25688 25152 25740 25158
rect 28368 25129 28396 25162
rect 25688 25094 25740 25100
rect 28354 25120 28410 25129
rect 25261 24508 25569 24517
rect 25261 24506 25267 24508
rect 25323 24506 25347 24508
rect 25403 24506 25427 24508
rect 25483 24506 25507 24508
rect 25563 24506 25569 24508
rect 25323 24454 25325 24506
rect 25505 24454 25507 24506
rect 25261 24452 25267 24454
rect 25323 24452 25347 24454
rect 25403 24452 25427 24454
rect 25483 24452 25507 24454
rect 25563 24452 25569 24454
rect 25261 24443 25569 24452
rect 25261 23420 25569 23429
rect 25261 23418 25267 23420
rect 25323 23418 25347 23420
rect 25403 23418 25427 23420
rect 25483 23418 25507 23420
rect 25563 23418 25569 23420
rect 25323 23366 25325 23418
rect 25505 23366 25507 23418
rect 25261 23364 25267 23366
rect 25323 23364 25347 23366
rect 25403 23364 25427 23366
rect 25483 23364 25507 23366
rect 25563 23364 25569 23366
rect 25261 23355 25569 23364
rect 25261 22332 25569 22341
rect 25261 22330 25267 22332
rect 25323 22330 25347 22332
rect 25403 22330 25427 22332
rect 25483 22330 25507 22332
rect 25563 22330 25569 22332
rect 25323 22278 25325 22330
rect 25505 22278 25507 22330
rect 25261 22276 25267 22278
rect 25323 22276 25347 22278
rect 25403 22276 25427 22278
rect 25483 22276 25507 22278
rect 25563 22276 25569 22278
rect 25261 22267 25569 22276
rect 25261 21244 25569 21253
rect 25261 21242 25267 21244
rect 25323 21242 25347 21244
rect 25403 21242 25427 21244
rect 25483 21242 25507 21244
rect 25563 21242 25569 21244
rect 25323 21190 25325 21242
rect 25505 21190 25507 21242
rect 25261 21188 25267 21190
rect 25323 21188 25347 21190
rect 25403 21188 25427 21190
rect 25483 21188 25507 21190
rect 25563 21188 25569 21190
rect 25261 21179 25569 21188
rect 25261 20156 25569 20165
rect 25261 20154 25267 20156
rect 25323 20154 25347 20156
rect 25403 20154 25427 20156
rect 25483 20154 25507 20156
rect 25563 20154 25569 20156
rect 25323 20102 25325 20154
rect 25505 20102 25507 20154
rect 25261 20100 25267 20102
rect 25323 20100 25347 20102
rect 25403 20100 25427 20102
rect 25483 20100 25507 20102
rect 25563 20100 25569 20102
rect 25261 20091 25569 20100
rect 25261 19068 25569 19077
rect 25261 19066 25267 19068
rect 25323 19066 25347 19068
rect 25403 19066 25427 19068
rect 25483 19066 25507 19068
rect 25563 19066 25569 19068
rect 25323 19014 25325 19066
rect 25505 19014 25507 19066
rect 25261 19012 25267 19014
rect 25323 19012 25347 19014
rect 25403 19012 25427 19014
rect 25483 19012 25507 19014
rect 25563 19012 25569 19014
rect 25261 19003 25569 19012
rect 25261 17980 25569 17989
rect 25261 17978 25267 17980
rect 25323 17978 25347 17980
rect 25403 17978 25427 17980
rect 25483 17978 25507 17980
rect 25563 17978 25569 17980
rect 25323 17926 25325 17978
rect 25505 17926 25507 17978
rect 25261 17924 25267 17926
rect 25323 17924 25347 17926
rect 25403 17924 25427 17926
rect 25483 17924 25507 17926
rect 25563 17924 25569 17926
rect 25261 17915 25569 17924
rect 25261 16892 25569 16901
rect 25261 16890 25267 16892
rect 25323 16890 25347 16892
rect 25403 16890 25427 16892
rect 25483 16890 25507 16892
rect 25563 16890 25569 16892
rect 25323 16838 25325 16890
rect 25505 16838 25507 16890
rect 25261 16836 25267 16838
rect 25323 16836 25347 16838
rect 25403 16836 25427 16838
rect 25483 16836 25507 16838
rect 25563 16836 25569 16838
rect 25261 16827 25569 16836
rect 23480 16584 23532 16590
rect 23480 16526 23532 16532
rect 22744 14476 22796 14482
rect 22744 14418 22796 14424
rect 21788 14172 22096 14181
rect 21788 14170 21794 14172
rect 21850 14170 21874 14172
rect 21930 14170 21954 14172
rect 22010 14170 22034 14172
rect 22090 14170 22096 14172
rect 21850 14118 21852 14170
rect 22032 14118 22034 14170
rect 21788 14116 21794 14118
rect 21850 14116 21874 14118
rect 21930 14116 21954 14118
rect 22010 14116 22034 14118
rect 22090 14116 22096 14118
rect 21788 14107 22096 14116
rect 18315 13628 18623 13637
rect 18315 13626 18321 13628
rect 18377 13626 18401 13628
rect 18457 13626 18481 13628
rect 18537 13626 18561 13628
rect 18617 13626 18623 13628
rect 18377 13574 18379 13626
rect 18559 13574 18561 13626
rect 18315 13572 18321 13574
rect 18377 13572 18401 13574
rect 18457 13572 18481 13574
rect 18537 13572 18561 13574
rect 18617 13572 18623 13574
rect 18315 13563 18623 13572
rect 21788 13084 22096 13093
rect 21788 13082 21794 13084
rect 21850 13082 21874 13084
rect 21930 13082 21954 13084
rect 22010 13082 22034 13084
rect 22090 13082 22096 13084
rect 21850 13030 21852 13082
rect 22032 13030 22034 13082
rect 21788 13028 21794 13030
rect 21850 13028 21874 13030
rect 21930 13028 21954 13030
rect 22010 13028 22034 13030
rect 22090 13028 22096 13030
rect 21788 13019 22096 13028
rect 22836 12980 22888 12986
rect 22836 12922 22888 12928
rect 17776 12912 17828 12918
rect 17776 12854 17828 12860
rect 17788 11898 17816 12854
rect 18315 12540 18623 12549
rect 18315 12538 18321 12540
rect 18377 12538 18401 12540
rect 18457 12538 18481 12540
rect 18537 12538 18561 12540
rect 18617 12538 18623 12540
rect 18377 12486 18379 12538
rect 18559 12486 18561 12538
rect 18315 12484 18321 12486
rect 18377 12484 18401 12486
rect 18457 12484 18481 12486
rect 18537 12484 18561 12486
rect 18617 12484 18623 12486
rect 18315 12475 18623 12484
rect 20076 12164 20128 12170
rect 20076 12106 20128 12112
rect 20168 12164 20220 12170
rect 20168 12106 20220 12112
rect 18880 12096 18932 12102
rect 18880 12038 18932 12044
rect 17776 11892 17828 11898
rect 17776 11834 17828 11840
rect 18315 11452 18623 11461
rect 18315 11450 18321 11452
rect 18377 11450 18401 11452
rect 18457 11450 18481 11452
rect 18537 11450 18561 11452
rect 18617 11450 18623 11452
rect 18377 11398 18379 11450
rect 18559 11398 18561 11450
rect 18315 11396 18321 11398
rect 18377 11396 18401 11398
rect 18457 11396 18481 11398
rect 18537 11396 18561 11398
rect 18617 11396 18623 11398
rect 18315 11387 18623 11396
rect 18315 10364 18623 10373
rect 18315 10362 18321 10364
rect 18377 10362 18401 10364
rect 18457 10362 18481 10364
rect 18537 10362 18561 10364
rect 18617 10362 18623 10364
rect 18377 10310 18379 10362
rect 18559 10310 18561 10362
rect 18315 10308 18321 10310
rect 18377 10308 18401 10310
rect 18457 10308 18481 10310
rect 18537 10308 18561 10310
rect 18617 10308 18623 10310
rect 18315 10299 18623 10308
rect 18315 9276 18623 9285
rect 18315 9274 18321 9276
rect 18377 9274 18401 9276
rect 18457 9274 18481 9276
rect 18537 9274 18561 9276
rect 18617 9274 18623 9276
rect 18377 9222 18379 9274
rect 18559 9222 18561 9274
rect 18315 9220 18321 9222
rect 18377 9220 18401 9222
rect 18457 9220 18481 9222
rect 18537 9220 18561 9222
rect 18617 9220 18623 9222
rect 18315 9211 18623 9220
rect 18315 8188 18623 8197
rect 18315 8186 18321 8188
rect 18377 8186 18401 8188
rect 18457 8186 18481 8188
rect 18537 8186 18561 8188
rect 18617 8186 18623 8188
rect 18377 8134 18379 8186
rect 18559 8134 18561 8186
rect 18315 8132 18321 8134
rect 18377 8132 18401 8134
rect 18457 8132 18481 8134
rect 18537 8132 18561 8134
rect 18617 8132 18623 8134
rect 18315 8123 18623 8132
rect 18315 7100 18623 7109
rect 18315 7098 18321 7100
rect 18377 7098 18401 7100
rect 18457 7098 18481 7100
rect 18537 7098 18561 7100
rect 18617 7098 18623 7100
rect 18377 7046 18379 7098
rect 18559 7046 18561 7098
rect 18315 7044 18321 7046
rect 18377 7044 18401 7046
rect 18457 7044 18481 7046
rect 18537 7044 18561 7046
rect 18617 7044 18623 7046
rect 18315 7035 18623 7044
rect 18315 6012 18623 6021
rect 18315 6010 18321 6012
rect 18377 6010 18401 6012
rect 18457 6010 18481 6012
rect 18537 6010 18561 6012
rect 18617 6010 18623 6012
rect 18377 5958 18379 6010
rect 18559 5958 18561 6010
rect 18315 5956 18321 5958
rect 18377 5956 18401 5958
rect 18457 5956 18481 5958
rect 18537 5956 18561 5958
rect 18617 5956 18623 5958
rect 18315 5947 18623 5956
rect 18315 4924 18623 4933
rect 18315 4922 18321 4924
rect 18377 4922 18401 4924
rect 18457 4922 18481 4924
rect 18537 4922 18561 4924
rect 18617 4922 18623 4924
rect 18377 4870 18379 4922
rect 18559 4870 18561 4922
rect 18315 4868 18321 4870
rect 18377 4868 18401 4870
rect 18457 4868 18481 4870
rect 18537 4868 18561 4870
rect 18617 4868 18623 4870
rect 18315 4859 18623 4868
rect 18315 3836 18623 3845
rect 18315 3834 18321 3836
rect 18377 3834 18401 3836
rect 18457 3834 18481 3836
rect 18537 3834 18561 3836
rect 18617 3834 18623 3836
rect 18377 3782 18379 3834
rect 18559 3782 18561 3834
rect 18315 3780 18321 3782
rect 18377 3780 18401 3782
rect 18457 3780 18481 3782
rect 18537 3780 18561 3782
rect 18617 3780 18623 3782
rect 18315 3771 18623 3780
rect 18892 3058 18920 12038
rect 19248 11552 19300 11558
rect 19248 11494 19300 11500
rect 19260 4758 19288 11494
rect 19248 4752 19300 4758
rect 19248 4694 19300 4700
rect 20088 3534 20116 12106
rect 20180 11898 20208 12106
rect 21788 11996 22096 12005
rect 21788 11994 21794 11996
rect 21850 11994 21874 11996
rect 21930 11994 21954 11996
rect 22010 11994 22034 11996
rect 22090 11994 22096 11996
rect 21850 11942 21852 11994
rect 22032 11942 22034 11994
rect 21788 11940 21794 11942
rect 21850 11940 21874 11942
rect 21930 11940 21954 11942
rect 22010 11940 22034 11942
rect 22090 11940 22096 11942
rect 21788 11931 22096 11940
rect 20168 11892 20220 11898
rect 20168 11834 20220 11840
rect 21788 10908 22096 10917
rect 21788 10906 21794 10908
rect 21850 10906 21874 10908
rect 21930 10906 21954 10908
rect 22010 10906 22034 10908
rect 22090 10906 22096 10908
rect 21850 10854 21852 10906
rect 22032 10854 22034 10906
rect 21788 10852 21794 10854
rect 21850 10852 21874 10854
rect 21930 10852 21954 10854
rect 22010 10852 22034 10854
rect 22090 10852 22096 10854
rect 21788 10843 22096 10852
rect 21788 9820 22096 9829
rect 21788 9818 21794 9820
rect 21850 9818 21874 9820
rect 21930 9818 21954 9820
rect 22010 9818 22034 9820
rect 22090 9818 22096 9820
rect 21850 9766 21852 9818
rect 22032 9766 22034 9818
rect 21788 9764 21794 9766
rect 21850 9764 21874 9766
rect 21930 9764 21954 9766
rect 22010 9764 22034 9766
rect 22090 9764 22096 9766
rect 21788 9755 22096 9764
rect 21788 8732 22096 8741
rect 21788 8730 21794 8732
rect 21850 8730 21874 8732
rect 21930 8730 21954 8732
rect 22010 8730 22034 8732
rect 22090 8730 22096 8732
rect 21850 8678 21852 8730
rect 22032 8678 22034 8730
rect 21788 8676 21794 8678
rect 21850 8676 21874 8678
rect 21930 8676 21954 8678
rect 22010 8676 22034 8678
rect 22090 8676 22096 8678
rect 21788 8667 22096 8676
rect 21788 7644 22096 7653
rect 21788 7642 21794 7644
rect 21850 7642 21874 7644
rect 21930 7642 21954 7644
rect 22010 7642 22034 7644
rect 22090 7642 22096 7644
rect 21850 7590 21852 7642
rect 22032 7590 22034 7642
rect 21788 7588 21794 7590
rect 21850 7588 21874 7590
rect 21930 7588 21954 7590
rect 22010 7588 22034 7590
rect 22090 7588 22096 7590
rect 21788 7579 22096 7588
rect 22376 6656 22428 6662
rect 22376 6598 22428 6604
rect 21788 6556 22096 6565
rect 21788 6554 21794 6556
rect 21850 6554 21874 6556
rect 21930 6554 21954 6556
rect 22010 6554 22034 6556
rect 22090 6554 22096 6556
rect 21850 6502 21852 6554
rect 22032 6502 22034 6554
rect 21788 6500 21794 6502
rect 21850 6500 21874 6502
rect 21930 6500 21954 6502
rect 22010 6500 22034 6502
rect 22090 6500 22096 6502
rect 21788 6491 22096 6500
rect 21788 5468 22096 5477
rect 21788 5466 21794 5468
rect 21850 5466 21874 5468
rect 21930 5466 21954 5468
rect 22010 5466 22034 5468
rect 22090 5466 22096 5468
rect 21850 5414 21852 5466
rect 22032 5414 22034 5466
rect 21788 5412 21794 5414
rect 21850 5412 21874 5414
rect 21930 5412 21954 5414
rect 22010 5412 22034 5414
rect 22090 5412 22096 5414
rect 21788 5403 22096 5412
rect 20902 4720 20958 4729
rect 20902 4655 20904 4664
rect 20956 4655 20958 4664
rect 20904 4626 20956 4632
rect 21788 4380 22096 4389
rect 21788 4378 21794 4380
rect 21850 4378 21874 4380
rect 21930 4378 21954 4380
rect 22010 4378 22034 4380
rect 22090 4378 22096 4380
rect 21850 4326 21852 4378
rect 22032 4326 22034 4378
rect 21788 4324 21794 4326
rect 21850 4324 21874 4326
rect 21930 4324 21954 4326
rect 22010 4324 22034 4326
rect 22090 4324 22096 4326
rect 21788 4315 22096 4324
rect 22388 4146 22416 6598
rect 22848 5710 22876 12922
rect 23492 12442 23520 16526
rect 25261 15804 25569 15813
rect 25261 15802 25267 15804
rect 25323 15802 25347 15804
rect 25403 15802 25427 15804
rect 25483 15802 25507 15804
rect 25563 15802 25569 15804
rect 25323 15750 25325 15802
rect 25505 15750 25507 15802
rect 25261 15748 25267 15750
rect 25323 15748 25347 15750
rect 25403 15748 25427 15750
rect 25483 15748 25507 15750
rect 25563 15748 25569 15750
rect 25261 15739 25569 15748
rect 25261 14716 25569 14725
rect 25261 14714 25267 14716
rect 25323 14714 25347 14716
rect 25403 14714 25427 14716
rect 25483 14714 25507 14716
rect 25563 14714 25569 14716
rect 25323 14662 25325 14714
rect 25505 14662 25507 14714
rect 25261 14660 25267 14662
rect 25323 14660 25347 14662
rect 25403 14660 25427 14662
rect 25483 14660 25507 14662
rect 25563 14660 25569 14662
rect 25261 14651 25569 14660
rect 25261 13628 25569 13637
rect 25261 13626 25267 13628
rect 25323 13626 25347 13628
rect 25403 13626 25427 13628
rect 25483 13626 25507 13628
rect 25563 13626 25569 13628
rect 25323 13574 25325 13626
rect 25505 13574 25507 13626
rect 25261 13572 25267 13574
rect 25323 13572 25347 13574
rect 25403 13572 25427 13574
rect 25483 13572 25507 13574
rect 25563 13572 25569 13574
rect 25261 13563 25569 13572
rect 25700 13258 25728 25094
rect 28354 25055 28410 25064
rect 28734 25052 29042 25061
rect 28734 25050 28740 25052
rect 28796 25050 28820 25052
rect 28876 25050 28900 25052
rect 28956 25050 28980 25052
rect 29036 25050 29042 25052
rect 28796 24998 28798 25050
rect 28978 24998 28980 25050
rect 28734 24996 28740 24998
rect 28796 24996 28820 24998
rect 28876 24996 28900 24998
rect 28956 24996 28980 24998
rect 29036 24996 29042 24998
rect 28734 24987 29042 24996
rect 28356 24744 28408 24750
rect 28356 24686 28408 24692
rect 28368 24313 28396 24686
rect 28354 24304 28410 24313
rect 28354 24239 28410 24248
rect 28734 23964 29042 23973
rect 28734 23962 28740 23964
rect 28796 23962 28820 23964
rect 28876 23962 28900 23964
rect 28956 23962 28980 23964
rect 29036 23962 29042 23964
rect 28796 23910 28798 23962
rect 28978 23910 28980 23962
rect 28734 23908 28740 23910
rect 28796 23908 28820 23910
rect 28876 23908 28900 23910
rect 28956 23908 28980 23910
rect 29036 23908 29042 23910
rect 28734 23899 29042 23908
rect 28724 23656 28776 23662
rect 28724 23598 28776 23604
rect 25780 23520 25832 23526
rect 28736 23497 28764 23598
rect 25780 23462 25832 23468
rect 28722 23488 28778 23497
rect 25688 13252 25740 13258
rect 25688 13194 25740 13200
rect 25792 12782 25820 23462
rect 28722 23423 28778 23432
rect 28356 23044 28408 23050
rect 28356 22986 28408 22992
rect 28368 22681 28396 22986
rect 28734 22876 29042 22885
rect 28734 22874 28740 22876
rect 28796 22874 28820 22876
rect 28876 22874 28900 22876
rect 28956 22874 28980 22876
rect 29036 22874 29042 22876
rect 28796 22822 28798 22874
rect 28978 22822 28980 22874
rect 28734 22820 28740 22822
rect 28796 22820 28820 22822
rect 28876 22820 28900 22822
rect 28956 22820 28980 22822
rect 29036 22820 29042 22822
rect 28734 22811 29042 22820
rect 28354 22672 28410 22681
rect 28354 22607 28410 22616
rect 28814 22128 28870 22137
rect 28814 22063 28816 22072
rect 28868 22063 28870 22072
rect 28816 22034 28868 22040
rect 28734 21788 29042 21797
rect 28734 21786 28740 21788
rect 28796 21786 28820 21788
rect 28876 21786 28900 21788
rect 28956 21786 28980 21788
rect 29036 21786 29042 21788
rect 28796 21734 28798 21786
rect 28978 21734 28980 21786
rect 28734 21732 28740 21734
rect 28796 21732 28820 21734
rect 28876 21732 28900 21734
rect 28956 21732 28980 21734
rect 29036 21732 29042 21734
rect 28734 21723 29042 21732
rect 28356 21480 28408 21486
rect 28356 21422 28408 21428
rect 28368 21049 28396 21422
rect 28354 21040 28410 21049
rect 28354 20975 28410 20984
rect 28734 20700 29042 20709
rect 28734 20698 28740 20700
rect 28796 20698 28820 20700
rect 28876 20698 28900 20700
rect 28956 20698 28980 20700
rect 29036 20698 29042 20700
rect 28796 20646 28798 20698
rect 28978 20646 28980 20698
rect 28734 20644 28740 20646
rect 28796 20644 28820 20646
rect 28876 20644 28900 20646
rect 28956 20644 28980 20646
rect 29036 20644 29042 20646
rect 28734 20635 29042 20644
rect 28356 20392 28408 20398
rect 28356 20334 28408 20340
rect 28368 20233 28396 20334
rect 28354 20224 28410 20233
rect 28354 20159 28410 20168
rect 28356 19780 28408 19786
rect 28356 19722 28408 19728
rect 28368 19417 28396 19722
rect 28734 19612 29042 19621
rect 28734 19610 28740 19612
rect 28796 19610 28820 19612
rect 28876 19610 28900 19612
rect 28956 19610 28980 19612
rect 29036 19610 29042 19612
rect 28796 19558 28798 19610
rect 28978 19558 28980 19610
rect 28734 19556 28740 19558
rect 28796 19556 28820 19558
rect 28876 19556 28900 19558
rect 28956 19556 28980 19558
rect 29036 19556 29042 19558
rect 28734 19547 29042 19556
rect 28354 19408 28410 19417
rect 28354 19343 28410 19352
rect 28814 18864 28870 18873
rect 28814 18799 28816 18808
rect 28868 18799 28870 18808
rect 28816 18770 28868 18776
rect 28734 18524 29042 18533
rect 28734 18522 28740 18524
rect 28796 18522 28820 18524
rect 28876 18522 28900 18524
rect 28956 18522 28980 18524
rect 29036 18522 29042 18524
rect 28796 18470 28798 18522
rect 28978 18470 28980 18522
rect 28734 18468 28740 18470
rect 28796 18468 28820 18470
rect 28876 18468 28900 18470
rect 28956 18468 28980 18470
rect 29036 18468 29042 18470
rect 28734 18459 29042 18468
rect 28356 18216 28408 18222
rect 28356 18158 28408 18164
rect 28368 17785 28396 18158
rect 28354 17776 28410 17785
rect 28354 17711 28410 17720
rect 28734 17436 29042 17445
rect 28734 17434 28740 17436
rect 28796 17434 28820 17436
rect 28876 17434 28900 17436
rect 28956 17434 28980 17436
rect 29036 17434 29042 17436
rect 28796 17382 28798 17434
rect 28978 17382 28980 17434
rect 28734 17380 28740 17382
rect 28796 17380 28820 17382
rect 28876 17380 28900 17382
rect 28956 17380 28980 17382
rect 29036 17380 29042 17382
rect 28734 17371 29042 17380
rect 28356 17128 28408 17134
rect 28356 17070 28408 17076
rect 28368 16969 28396 17070
rect 28354 16960 28410 16969
rect 28354 16895 28410 16904
rect 28356 16516 28408 16522
rect 28356 16458 28408 16464
rect 28368 16153 28396 16458
rect 28734 16348 29042 16357
rect 28734 16346 28740 16348
rect 28796 16346 28820 16348
rect 28876 16346 28900 16348
rect 28956 16346 28980 16348
rect 29036 16346 29042 16348
rect 28796 16294 28798 16346
rect 28978 16294 28980 16346
rect 28734 16292 28740 16294
rect 28796 16292 28820 16294
rect 28876 16292 28900 16294
rect 28956 16292 28980 16294
rect 29036 16292 29042 16294
rect 28734 16283 29042 16292
rect 28354 16144 28410 16153
rect 28354 16079 28410 16088
rect 28356 15428 28408 15434
rect 28356 15370 28408 15376
rect 26976 15360 27028 15366
rect 28368 15337 28396 15370
rect 26976 15302 27028 15308
rect 28354 15328 28410 15337
rect 26988 14521 27016 15302
rect 28354 15263 28410 15272
rect 28734 15260 29042 15269
rect 28734 15258 28740 15260
rect 28796 15258 28820 15260
rect 28876 15258 28900 15260
rect 28956 15258 28980 15260
rect 29036 15258 29042 15260
rect 28796 15206 28798 15258
rect 28978 15206 28980 15258
rect 28734 15204 28740 15206
rect 28796 15204 28820 15206
rect 28876 15204 28900 15206
rect 28956 15204 28980 15206
rect 29036 15204 29042 15206
rect 28734 15195 29042 15204
rect 28356 14952 28408 14958
rect 28356 14894 28408 14900
rect 28368 14521 28396 14894
rect 26974 14512 27030 14521
rect 26974 14447 27030 14456
rect 28354 14512 28410 14521
rect 28354 14447 28410 14456
rect 28734 14172 29042 14181
rect 28734 14170 28740 14172
rect 28796 14170 28820 14172
rect 28876 14170 28900 14172
rect 28956 14170 28980 14172
rect 29036 14170 29042 14172
rect 28796 14118 28798 14170
rect 28978 14118 28980 14170
rect 28734 14116 28740 14118
rect 28796 14116 28820 14118
rect 28876 14116 28900 14118
rect 28956 14116 28980 14118
rect 29036 14116 29042 14118
rect 28734 14107 29042 14116
rect 28356 13864 28408 13870
rect 28356 13806 28408 13812
rect 28368 13705 28396 13806
rect 28354 13696 28410 13705
rect 28354 13631 28410 13640
rect 28356 13252 28408 13258
rect 28356 13194 28408 13200
rect 28368 12889 28396 13194
rect 28734 13084 29042 13093
rect 28734 13082 28740 13084
rect 28796 13082 28820 13084
rect 28876 13082 28900 13084
rect 28956 13082 28980 13084
rect 29036 13082 29042 13084
rect 28796 13030 28798 13082
rect 28978 13030 28980 13082
rect 28734 13028 28740 13030
rect 28796 13028 28820 13030
rect 28876 13028 28900 13030
rect 28956 13028 28980 13030
rect 29036 13028 29042 13030
rect 28734 13019 29042 13028
rect 28354 12880 28410 12889
rect 28354 12815 28410 12824
rect 25780 12776 25832 12782
rect 25780 12718 25832 12724
rect 25261 12540 25569 12549
rect 25261 12538 25267 12540
rect 25323 12538 25347 12540
rect 25403 12538 25427 12540
rect 25483 12538 25507 12540
rect 25563 12538 25569 12540
rect 25323 12486 25325 12538
rect 25505 12486 25507 12538
rect 25261 12484 25267 12486
rect 25323 12484 25347 12486
rect 25403 12484 25427 12486
rect 25483 12484 25507 12486
rect 25563 12484 25569 12486
rect 25261 12475 25569 12484
rect 23480 12436 23532 12442
rect 23480 12378 23532 12384
rect 28356 12164 28408 12170
rect 28356 12106 28408 12112
rect 28368 12073 28396 12106
rect 28354 12064 28410 12073
rect 28354 11999 28410 12008
rect 28734 11996 29042 12005
rect 28734 11994 28740 11996
rect 28796 11994 28820 11996
rect 28876 11994 28900 11996
rect 28956 11994 28980 11996
rect 29036 11994 29042 11996
rect 28796 11942 28798 11994
rect 28978 11942 28980 11994
rect 28734 11940 28740 11942
rect 28796 11940 28820 11942
rect 28876 11940 28900 11942
rect 28956 11940 28980 11942
rect 29036 11940 29042 11942
rect 28734 11931 29042 11940
rect 28356 11688 28408 11694
rect 28356 11630 28408 11636
rect 26700 11552 26752 11558
rect 26700 11494 26752 11500
rect 25261 11452 25569 11461
rect 25261 11450 25267 11452
rect 25323 11450 25347 11452
rect 25403 11450 25427 11452
rect 25483 11450 25507 11452
rect 25563 11450 25569 11452
rect 25323 11398 25325 11450
rect 25505 11398 25507 11450
rect 25261 11396 25267 11398
rect 25323 11396 25347 11398
rect 25403 11396 25427 11398
rect 25483 11396 25507 11398
rect 25563 11396 25569 11398
rect 25261 11387 25569 11396
rect 26712 10810 26740 11494
rect 28368 11257 28396 11630
rect 28354 11248 28410 11257
rect 28354 11183 28410 11192
rect 28734 10908 29042 10917
rect 28734 10906 28740 10908
rect 28796 10906 28820 10908
rect 28876 10906 28900 10908
rect 28956 10906 28980 10908
rect 29036 10906 29042 10908
rect 28796 10854 28798 10906
rect 28978 10854 28980 10906
rect 28734 10852 28740 10854
rect 28796 10852 28820 10854
rect 28876 10852 28900 10854
rect 28956 10852 28980 10854
rect 29036 10852 29042 10854
rect 28734 10843 29042 10852
rect 26700 10804 26752 10810
rect 26700 10746 26752 10752
rect 28356 10600 28408 10606
rect 28356 10542 28408 10548
rect 28368 10441 28396 10542
rect 28354 10432 28410 10441
rect 25261 10364 25569 10373
rect 28354 10367 28410 10376
rect 25261 10362 25267 10364
rect 25323 10362 25347 10364
rect 25403 10362 25427 10364
rect 25483 10362 25507 10364
rect 25563 10362 25569 10364
rect 25323 10310 25325 10362
rect 25505 10310 25507 10362
rect 25261 10308 25267 10310
rect 25323 10308 25347 10310
rect 25403 10308 25427 10310
rect 25483 10308 25507 10310
rect 25563 10308 25569 10310
rect 25261 10299 25569 10308
rect 28356 9988 28408 9994
rect 28356 9930 28408 9936
rect 28368 9625 28396 9930
rect 28734 9820 29042 9829
rect 28734 9818 28740 9820
rect 28796 9818 28820 9820
rect 28876 9818 28900 9820
rect 28956 9818 28980 9820
rect 29036 9818 29042 9820
rect 28796 9766 28798 9818
rect 28978 9766 28980 9818
rect 28734 9764 28740 9766
rect 28796 9764 28820 9766
rect 28876 9764 28900 9766
rect 28956 9764 28980 9766
rect 29036 9764 29042 9766
rect 28734 9755 29042 9764
rect 28354 9616 28410 9625
rect 28354 9551 28410 9560
rect 23848 9444 23900 9450
rect 23848 9386 23900 9392
rect 23480 9172 23532 9178
rect 23480 9114 23532 9120
rect 23388 8288 23440 8294
rect 23388 8230 23440 8236
rect 23400 8022 23428 8230
rect 23388 8016 23440 8022
rect 23388 7958 23440 7964
rect 22836 5704 22888 5710
rect 22836 5646 22888 5652
rect 23492 5234 23520 9114
rect 23756 6316 23808 6322
rect 23756 6258 23808 6264
rect 23768 6118 23796 6258
rect 23756 6112 23808 6118
rect 23756 6054 23808 6060
rect 23480 5228 23532 5234
rect 23480 5170 23532 5176
rect 22928 4820 22980 4826
rect 22928 4762 22980 4768
rect 22940 4622 22968 4762
rect 22928 4616 22980 4622
rect 22928 4558 22980 4564
rect 22560 4548 22612 4554
rect 22560 4490 22612 4496
rect 22572 4282 22600 4490
rect 23664 4480 23716 4486
rect 23664 4422 23716 4428
rect 22560 4276 22612 4282
rect 22560 4218 22612 4224
rect 23296 4208 23348 4214
rect 23296 4150 23348 4156
rect 22376 4140 22428 4146
rect 22376 4082 22428 4088
rect 22284 4072 22336 4078
rect 22284 4014 22336 4020
rect 23112 4072 23164 4078
rect 23112 4014 23164 4020
rect 20352 3664 20404 3670
rect 20352 3606 20404 3612
rect 21456 3664 21508 3670
rect 21456 3606 21508 3612
rect 20076 3528 20128 3534
rect 20076 3470 20128 3476
rect 18880 3052 18932 3058
rect 18880 2994 18932 3000
rect 18315 2748 18623 2757
rect 18315 2746 18321 2748
rect 18377 2746 18401 2748
rect 18457 2746 18481 2748
rect 18537 2746 18561 2748
rect 18617 2746 18623 2748
rect 18377 2694 18379 2746
rect 18559 2694 18561 2746
rect 18315 2692 18321 2694
rect 18377 2692 18401 2694
rect 18457 2692 18481 2694
rect 18537 2692 18561 2694
rect 18617 2692 18623 2694
rect 18315 2683 18623 2692
rect 20364 2446 20392 3606
rect 21364 2916 21416 2922
rect 21364 2858 21416 2864
rect 20720 2508 20772 2514
rect 20720 2450 20772 2456
rect 21180 2508 21232 2514
rect 21180 2450 21232 2456
rect 17684 2440 17736 2446
rect 17684 2382 17736 2388
rect 20352 2440 20404 2446
rect 20352 2382 20404 2388
rect 18880 2372 18932 2378
rect 18880 2314 18932 2320
rect 15200 2304 15252 2310
rect 15200 2246 15252 2252
rect 14842 2204 15150 2213
rect 14842 2202 14848 2204
rect 14904 2202 14928 2204
rect 14984 2202 15008 2204
rect 15064 2202 15088 2204
rect 15144 2202 15150 2204
rect 14904 2150 14906 2202
rect 15086 2150 15088 2202
rect 14842 2148 14848 2150
rect 14904 2148 14928 2150
rect 14984 2148 15008 2150
rect 15064 2148 15088 2150
rect 15144 2148 15150 2150
rect 14842 2139 15150 2148
rect 18892 2106 18920 2314
rect 18880 2100 18932 2106
rect 18880 2042 18932 2048
rect 14648 1964 14700 1970
rect 14648 1906 14700 1912
rect 20732 1442 20760 2450
rect 20640 1414 20760 1442
rect 20640 800 20668 1414
rect 21192 1170 21220 2450
rect 20916 1142 21220 1170
rect 20916 800 20944 1142
rect 21376 1034 21404 2858
rect 21192 1006 21404 1034
rect 21192 800 21220 1006
rect 21468 800 21496 3606
rect 21788 3292 22096 3301
rect 21788 3290 21794 3292
rect 21850 3290 21874 3292
rect 21930 3290 21954 3292
rect 22010 3290 22034 3292
rect 22090 3290 22096 3292
rect 21850 3238 21852 3290
rect 22032 3238 22034 3290
rect 21788 3236 21794 3238
rect 21850 3236 21874 3238
rect 21930 3236 21954 3238
rect 22010 3236 22034 3238
rect 22090 3236 22096 3238
rect 21788 3227 22096 3236
rect 21824 3052 21876 3058
rect 21824 2994 21876 3000
rect 21836 2961 21864 2994
rect 21822 2952 21878 2961
rect 21822 2887 21878 2896
rect 21548 2848 21600 2854
rect 21548 2790 21600 2796
rect 21560 1850 21588 2790
rect 21788 2204 22096 2213
rect 21788 2202 21794 2204
rect 21850 2202 21874 2204
rect 21930 2202 21954 2204
rect 22010 2202 22034 2204
rect 22090 2202 22096 2204
rect 21850 2150 21852 2202
rect 22032 2150 22034 2202
rect 21788 2148 21794 2150
rect 21850 2148 21874 2150
rect 21930 2148 21954 2150
rect 22010 2148 22034 2150
rect 22090 2148 22096 2150
rect 21788 2139 22096 2148
rect 21560 1822 21772 1850
rect 21744 800 21772 1822
rect 22008 1420 22060 1426
rect 22008 1362 22060 1368
rect 22020 800 22048 1362
rect 22296 800 22324 4014
rect 22836 3596 22888 3602
rect 22836 3538 22888 3544
rect 22560 2984 22612 2990
rect 22560 2926 22612 2932
rect 22572 800 22600 2926
rect 22848 800 22876 3538
rect 23124 800 23152 4014
rect 23308 3058 23336 4150
rect 23388 3188 23440 3194
rect 23388 3130 23440 3136
rect 23296 3052 23348 3058
rect 23296 2994 23348 3000
rect 23400 2961 23428 3130
rect 23386 2952 23442 2961
rect 23386 2887 23442 2896
rect 23388 2372 23440 2378
rect 23388 2314 23440 2320
rect 23400 800 23428 2314
rect 23676 800 23704 4422
rect 23768 3942 23796 6054
rect 23860 4146 23888 9386
rect 25780 9376 25832 9382
rect 25780 9318 25832 9324
rect 25261 9276 25569 9285
rect 25261 9274 25267 9276
rect 25323 9274 25347 9276
rect 25403 9274 25427 9276
rect 25483 9274 25507 9276
rect 25563 9274 25569 9276
rect 25323 9222 25325 9274
rect 25505 9222 25507 9274
rect 25261 9220 25267 9222
rect 25323 9220 25347 9222
rect 25403 9220 25427 9222
rect 25483 9220 25507 9222
rect 25563 9220 25569 9222
rect 25261 9211 25569 9220
rect 25261 8188 25569 8197
rect 25261 8186 25267 8188
rect 25323 8186 25347 8188
rect 25403 8186 25427 8188
rect 25483 8186 25507 8188
rect 25563 8186 25569 8188
rect 25323 8134 25325 8186
rect 25505 8134 25507 8186
rect 25261 8132 25267 8134
rect 25323 8132 25347 8134
rect 25403 8132 25427 8134
rect 25483 8132 25507 8134
rect 25563 8132 25569 8134
rect 25261 8123 25569 8132
rect 24400 7540 24452 7546
rect 24400 7482 24452 7488
rect 24122 6216 24178 6225
rect 24122 6151 24178 6160
rect 24136 4146 24164 6151
rect 23848 4140 23900 4146
rect 23848 4082 23900 4088
rect 24124 4140 24176 4146
rect 24124 4082 24176 4088
rect 23940 4004 23992 4010
rect 23940 3946 23992 3952
rect 23756 3936 23808 3942
rect 23756 3878 23808 3884
rect 23952 800 23980 3946
rect 24136 3738 24164 4082
rect 24124 3732 24176 3738
rect 24124 3674 24176 3680
rect 24412 3534 24440 7482
rect 25261 7100 25569 7109
rect 25261 7098 25267 7100
rect 25323 7098 25347 7100
rect 25403 7098 25427 7100
rect 25483 7098 25507 7100
rect 25563 7098 25569 7100
rect 25323 7046 25325 7098
rect 25505 7046 25507 7098
rect 25261 7044 25267 7046
rect 25323 7044 25347 7046
rect 25403 7044 25427 7046
rect 25483 7044 25507 7046
rect 25563 7044 25569 7046
rect 25261 7035 25569 7044
rect 24952 6928 25004 6934
rect 24952 6870 25004 6876
rect 24584 6316 24636 6322
rect 24584 6258 24636 6264
rect 24596 5370 24624 6258
rect 24676 6248 24728 6254
rect 24676 6190 24728 6196
rect 24584 5364 24636 5370
rect 24584 5306 24636 5312
rect 24400 3528 24452 3534
rect 24400 3470 24452 3476
rect 24216 3460 24268 3466
rect 24216 3402 24268 3408
rect 24228 800 24256 3402
rect 24688 3097 24716 6190
rect 24860 6180 24912 6186
rect 24860 6122 24912 6128
rect 24872 5234 24900 6122
rect 24860 5228 24912 5234
rect 24860 5170 24912 5176
rect 24768 5160 24820 5166
rect 24768 5102 24820 5108
rect 24674 3088 24730 3097
rect 24674 3023 24730 3032
rect 24676 2916 24728 2922
rect 24676 2858 24728 2864
rect 24584 2508 24636 2514
rect 24584 2450 24636 2456
rect 24596 1562 24624 2450
rect 24584 1556 24636 1562
rect 24584 1498 24636 1504
rect 24688 1442 24716 2858
rect 24504 1414 24716 1442
rect 24504 800 24532 1414
rect 24780 800 24808 5102
rect 24860 4548 24912 4554
rect 24860 4490 24912 4496
rect 24872 1902 24900 4490
rect 24964 3058 24992 6870
rect 25261 6012 25569 6021
rect 25261 6010 25267 6012
rect 25323 6010 25347 6012
rect 25403 6010 25427 6012
rect 25483 6010 25507 6012
rect 25563 6010 25569 6012
rect 25323 5958 25325 6010
rect 25505 5958 25507 6010
rect 25261 5956 25267 5958
rect 25323 5956 25347 5958
rect 25403 5956 25427 5958
rect 25483 5956 25507 5958
rect 25563 5956 25569 5958
rect 25261 5947 25569 5956
rect 25261 4924 25569 4933
rect 25261 4922 25267 4924
rect 25323 4922 25347 4924
rect 25403 4922 25427 4924
rect 25483 4922 25507 4924
rect 25563 4922 25569 4924
rect 25323 4870 25325 4922
rect 25505 4870 25507 4922
rect 25261 4868 25267 4870
rect 25323 4868 25347 4870
rect 25403 4868 25427 4870
rect 25483 4868 25507 4870
rect 25563 4868 25569 4870
rect 25261 4859 25569 4868
rect 25136 4684 25188 4690
rect 25136 4626 25188 4632
rect 25148 4154 25176 4626
rect 25056 4126 25176 4154
rect 25792 4154 25820 9318
rect 28814 9072 28870 9081
rect 26608 9036 26660 9042
rect 28814 9007 28816 9016
rect 26608 8978 26660 8984
rect 28868 9007 28870 9016
rect 28816 8978 28868 8984
rect 26148 6248 26200 6254
rect 26148 6190 26200 6196
rect 25964 5160 26016 5166
rect 25964 5102 26016 5108
rect 25870 4720 25926 4729
rect 25870 4655 25926 4664
rect 25884 4622 25912 4655
rect 25872 4616 25924 4622
rect 25872 4558 25924 4564
rect 25792 4126 25912 4154
rect 24952 3052 25004 3058
rect 24952 2994 25004 3000
rect 24860 1896 24912 1902
rect 24860 1838 24912 1844
rect 25056 800 25084 4126
rect 25136 4004 25188 4010
rect 25136 3946 25188 3952
rect 25148 2122 25176 3946
rect 25596 3936 25648 3942
rect 25596 3878 25648 3884
rect 25261 3836 25569 3845
rect 25261 3834 25267 3836
rect 25323 3834 25347 3836
rect 25403 3834 25427 3836
rect 25483 3834 25507 3836
rect 25563 3834 25569 3836
rect 25323 3782 25325 3834
rect 25505 3782 25507 3834
rect 25261 3780 25267 3782
rect 25323 3780 25347 3782
rect 25403 3780 25427 3782
rect 25483 3780 25507 3782
rect 25563 3780 25569 3782
rect 25261 3771 25569 3780
rect 25261 2748 25569 2757
rect 25261 2746 25267 2748
rect 25323 2746 25347 2748
rect 25403 2746 25427 2748
rect 25483 2746 25507 2748
rect 25563 2746 25569 2748
rect 25323 2694 25325 2746
rect 25505 2694 25507 2746
rect 25261 2692 25267 2694
rect 25323 2692 25347 2694
rect 25403 2692 25427 2694
rect 25483 2692 25507 2694
rect 25563 2692 25569 2694
rect 25261 2683 25569 2692
rect 25608 2417 25636 3878
rect 25884 3534 25912 4126
rect 25872 3528 25924 3534
rect 25872 3470 25924 3476
rect 25594 2408 25650 2417
rect 25594 2343 25650 2352
rect 25976 2122 26004 5102
rect 25148 2094 25360 2122
rect 25332 800 25360 2094
rect 25596 2100 25648 2106
rect 25596 2042 25648 2048
rect 25884 2094 26004 2122
rect 25608 800 25636 2042
rect 25884 800 25912 2094
rect 26160 800 26188 6190
rect 26424 5772 26476 5778
rect 26424 5714 26476 5720
rect 26240 2304 26292 2310
rect 26240 2246 26292 2252
rect 26252 1970 26280 2246
rect 26436 2106 26464 5714
rect 26516 5092 26568 5098
rect 26516 5034 26568 5040
rect 26528 2122 26556 5034
rect 26620 4146 26648 8978
rect 27160 8968 27212 8974
rect 27160 8910 27212 8916
rect 26884 8900 26936 8906
rect 26884 8842 26936 8848
rect 26896 8294 26924 8842
rect 27172 8634 27200 8910
rect 28734 8732 29042 8741
rect 28734 8730 28740 8732
rect 28796 8730 28820 8732
rect 28876 8730 28900 8732
rect 28956 8730 28980 8732
rect 29036 8730 29042 8732
rect 28796 8678 28798 8730
rect 28978 8678 28980 8730
rect 28734 8676 28740 8678
rect 28796 8676 28820 8678
rect 28876 8676 28900 8678
rect 28956 8676 28980 8678
rect 29036 8676 29042 8678
rect 28734 8667 29042 8676
rect 27160 8628 27212 8634
rect 27160 8570 27212 8576
rect 28356 8424 28408 8430
rect 28356 8366 28408 8372
rect 26896 8266 27016 8294
rect 26884 6724 26936 6730
rect 26884 6666 26936 6672
rect 26700 5908 26752 5914
rect 26700 5850 26752 5856
rect 26712 5370 26740 5850
rect 26700 5364 26752 5370
rect 26700 5306 26752 5312
rect 26608 4140 26660 4146
rect 26608 4082 26660 4088
rect 26896 3913 26924 6666
rect 26882 3904 26938 3913
rect 26882 3839 26938 3848
rect 26792 3120 26844 3126
rect 26792 3062 26844 3068
rect 26424 2100 26476 2106
rect 26528 2094 26740 2122
rect 26424 2042 26476 2048
rect 26240 1964 26292 1970
rect 26240 1906 26292 1912
rect 26424 1896 26476 1902
rect 26424 1838 26476 1844
rect 26436 800 26464 1838
rect 26712 800 26740 2094
rect 26804 1034 26832 3062
rect 26988 3058 27016 8266
rect 27160 8084 27212 8090
rect 27160 8026 27212 8032
rect 27172 7410 27200 8026
rect 28368 7993 28396 8366
rect 28354 7984 28410 7993
rect 27620 7948 27672 7954
rect 28354 7919 28410 7928
rect 27620 7890 27672 7896
rect 27160 7404 27212 7410
rect 27160 7346 27212 7352
rect 27252 5636 27304 5642
rect 27252 5578 27304 5584
rect 27160 4140 27212 4146
rect 27160 4082 27212 4088
rect 27172 3738 27200 4082
rect 27160 3732 27212 3738
rect 27160 3674 27212 3680
rect 27068 3392 27120 3398
rect 27068 3334 27120 3340
rect 26976 3052 27028 3058
rect 26976 2994 27028 3000
rect 27080 1714 27108 3334
rect 27264 2106 27292 5578
rect 27632 4154 27660 7890
rect 28734 7644 29042 7653
rect 28734 7642 28740 7644
rect 28796 7642 28820 7644
rect 28876 7642 28900 7644
rect 28956 7642 28980 7644
rect 29036 7642 29042 7644
rect 28796 7590 28798 7642
rect 28978 7590 28980 7642
rect 28734 7588 28740 7590
rect 28796 7588 28820 7590
rect 28876 7588 28900 7590
rect 28956 7588 28980 7590
rect 29036 7588 29042 7590
rect 28734 7579 29042 7588
rect 29184 7472 29236 7478
rect 29184 7414 29236 7420
rect 28356 7336 28408 7342
rect 28356 7278 28408 7284
rect 28368 7177 28396 7278
rect 28354 7168 28410 7177
rect 28354 7103 28410 7112
rect 28356 6724 28408 6730
rect 28356 6666 28408 6672
rect 28368 6361 28396 6666
rect 28734 6556 29042 6565
rect 28734 6554 28740 6556
rect 28796 6554 28820 6556
rect 28876 6554 28900 6556
rect 28956 6554 28980 6556
rect 29036 6554 29042 6556
rect 28796 6502 28798 6554
rect 28978 6502 28980 6554
rect 28734 6500 28740 6502
rect 28796 6500 28820 6502
rect 28876 6500 28900 6502
rect 28956 6500 28980 6502
rect 29036 6500 29042 6502
rect 28734 6491 29042 6500
rect 28354 6352 28410 6361
rect 28354 6287 28410 6296
rect 28632 6248 28684 6254
rect 28632 6190 28684 6196
rect 28080 5024 28132 5030
rect 28080 4966 28132 4972
rect 27540 4126 27660 4154
rect 27252 2100 27304 2106
rect 27252 2042 27304 2048
rect 27080 1686 27292 1714
rect 26804 1006 27016 1034
rect 26988 800 27016 1006
rect 27264 800 27292 1686
rect 27540 800 27568 4126
rect 27804 2100 27856 2106
rect 27804 2042 27856 2048
rect 27816 800 27844 2042
rect 28092 800 28120 4966
rect 28644 4706 28672 6190
rect 28814 5808 28870 5817
rect 28814 5743 28816 5752
rect 28868 5743 28870 5752
rect 28816 5714 28868 5720
rect 28734 5468 29042 5477
rect 28734 5466 28740 5468
rect 28796 5466 28820 5468
rect 28876 5466 28900 5468
rect 28956 5466 28980 5468
rect 29036 5466 29042 5468
rect 28796 5414 28798 5466
rect 28978 5414 28980 5466
rect 28734 5412 28740 5414
rect 28796 5412 28820 5414
rect 28876 5412 28900 5414
rect 28956 5412 28980 5414
rect 29036 5412 29042 5414
rect 28734 5403 29042 5412
rect 28722 4720 28778 4729
rect 28644 4678 28722 4706
rect 28722 4655 28778 4664
rect 28734 4380 29042 4389
rect 28734 4378 28740 4380
rect 28796 4378 28820 4380
rect 28876 4378 28900 4380
rect 28956 4378 28980 4380
rect 29036 4378 29042 4380
rect 28796 4326 28798 4378
rect 28978 4326 28980 4378
rect 28734 4324 28740 4326
rect 28796 4324 28820 4326
rect 28876 4324 28900 4326
rect 28956 4324 28980 4326
rect 29036 4324 29042 4326
rect 28734 4315 29042 4324
rect 28356 4276 28408 4282
rect 28356 4218 28408 4224
rect 28368 800 28396 4218
rect 28734 3292 29042 3301
rect 28734 3290 28740 3292
rect 28796 3290 28820 3292
rect 28876 3290 28900 3292
rect 28956 3290 28980 3292
rect 29036 3290 29042 3292
rect 28796 3238 28798 3290
rect 28978 3238 28980 3290
rect 28734 3236 28740 3238
rect 28796 3236 28820 3238
rect 28876 3236 28900 3238
rect 28956 3236 28980 3238
rect 29036 3236 29042 3238
rect 28734 3227 29042 3236
rect 28630 2952 28686 2961
rect 28630 2887 28686 2896
rect 28644 800 28672 2887
rect 28734 2204 29042 2213
rect 28734 2202 28740 2204
rect 28796 2202 28820 2204
rect 28876 2202 28900 2204
rect 28956 2202 28980 2204
rect 29036 2202 29042 2204
rect 28796 2150 28798 2202
rect 28978 2150 28980 2202
rect 28734 2148 28740 2150
rect 28796 2148 28820 2150
rect 28876 2148 28900 2150
rect 28956 2148 28980 2150
rect 29036 2148 29042 2150
rect 28734 2139 29042 2148
rect 28908 2032 28960 2038
rect 28908 1974 28960 1980
rect 28920 800 28948 1974
rect 29196 800 29224 7414
rect 29460 3528 29512 3534
rect 29460 3470 29512 3476
rect 29472 800 29500 3470
rect 478 0 534 800
rect 754 0 810 800
rect 1030 0 1086 800
rect 1306 0 1362 800
rect 1582 0 1638 800
rect 1858 0 1914 800
rect 2134 0 2190 800
rect 2410 0 2466 800
rect 2686 0 2742 800
rect 2962 0 3018 800
rect 3238 0 3294 800
rect 3514 0 3570 800
rect 3790 0 3846 800
rect 4066 0 4122 800
rect 4342 0 4398 800
rect 4618 0 4674 800
rect 4894 0 4950 800
rect 5170 0 5226 800
rect 5446 0 5502 800
rect 5722 0 5778 800
rect 5998 0 6054 800
rect 6274 0 6330 800
rect 6550 0 6606 800
rect 6826 0 6882 800
rect 7102 0 7158 800
rect 7378 0 7434 800
rect 7654 0 7710 800
rect 7930 0 7986 800
rect 8206 0 8262 800
rect 8482 0 8538 800
rect 8758 0 8814 800
rect 9034 0 9090 800
rect 9310 0 9366 800
rect 9586 0 9642 800
rect 9862 0 9918 800
rect 10138 0 10194 800
rect 10414 0 10470 800
rect 10690 0 10746 800
rect 10966 0 11022 800
rect 11242 0 11298 800
rect 11518 0 11574 800
rect 11794 0 11850 800
rect 12070 0 12126 800
rect 12346 0 12402 800
rect 12622 0 12678 800
rect 12898 0 12954 800
rect 13174 0 13230 800
rect 13450 0 13506 800
rect 13726 0 13782 800
rect 14002 0 14058 800
rect 14278 0 14334 800
rect 14554 0 14610 800
rect 14830 0 14886 800
rect 15106 0 15162 800
rect 15382 0 15438 800
rect 15658 0 15714 800
rect 15934 0 15990 800
rect 16210 0 16266 800
rect 16486 0 16542 800
rect 16762 0 16818 800
rect 17038 0 17094 800
rect 17314 0 17370 800
rect 17590 0 17646 800
rect 17866 0 17922 800
rect 18142 0 18198 800
rect 18418 0 18474 800
rect 18694 0 18750 800
rect 18970 0 19026 800
rect 19246 0 19302 800
rect 19522 0 19578 800
rect 19798 0 19854 800
rect 20074 0 20130 800
rect 20350 0 20406 800
rect 20626 0 20682 800
rect 20902 0 20958 800
rect 21178 0 21234 800
rect 21454 0 21510 800
rect 21730 0 21786 800
rect 22006 0 22062 800
rect 22282 0 22338 800
rect 22558 0 22614 800
rect 22834 0 22890 800
rect 23110 0 23166 800
rect 23386 0 23442 800
rect 23662 0 23718 800
rect 23938 0 23994 800
rect 24214 0 24270 800
rect 24490 0 24546 800
rect 24766 0 24822 800
rect 25042 0 25098 800
rect 25318 0 25374 800
rect 25594 0 25650 800
rect 25870 0 25926 800
rect 26146 0 26202 800
rect 26422 0 26478 800
rect 26698 0 26754 800
rect 26974 0 27030 800
rect 27250 0 27306 800
rect 27526 0 27582 800
rect 27802 0 27858 800
rect 28078 0 28134 800
rect 28354 0 28410 800
rect 28630 0 28686 800
rect 28906 0 28962 800
rect 29182 0 29238 800
rect 29458 0 29514 800
<< via2 >>
rect 4429 27770 4485 27772
rect 4509 27770 4565 27772
rect 4589 27770 4645 27772
rect 4669 27770 4725 27772
rect 4429 27718 4475 27770
rect 4475 27718 4485 27770
rect 4509 27718 4539 27770
rect 4539 27718 4551 27770
rect 4551 27718 4565 27770
rect 4589 27718 4603 27770
rect 4603 27718 4615 27770
rect 4615 27718 4645 27770
rect 4669 27718 4679 27770
rect 4679 27718 4725 27770
rect 4429 27716 4485 27718
rect 4509 27716 4565 27718
rect 4589 27716 4645 27718
rect 4669 27716 4725 27718
rect 11375 27770 11431 27772
rect 11455 27770 11511 27772
rect 11535 27770 11591 27772
rect 11615 27770 11671 27772
rect 11375 27718 11421 27770
rect 11421 27718 11431 27770
rect 11455 27718 11485 27770
rect 11485 27718 11497 27770
rect 11497 27718 11511 27770
rect 11535 27718 11549 27770
rect 11549 27718 11561 27770
rect 11561 27718 11591 27770
rect 11615 27718 11625 27770
rect 11625 27718 11671 27770
rect 11375 27716 11431 27718
rect 11455 27716 11511 27718
rect 11535 27716 11591 27718
rect 11615 27716 11671 27718
rect 18321 27770 18377 27772
rect 18401 27770 18457 27772
rect 18481 27770 18537 27772
rect 18561 27770 18617 27772
rect 18321 27718 18367 27770
rect 18367 27718 18377 27770
rect 18401 27718 18431 27770
rect 18431 27718 18443 27770
rect 18443 27718 18457 27770
rect 18481 27718 18495 27770
rect 18495 27718 18507 27770
rect 18507 27718 18537 27770
rect 18561 27718 18571 27770
rect 18571 27718 18617 27770
rect 18321 27716 18377 27718
rect 18401 27716 18457 27718
rect 18481 27716 18537 27718
rect 18561 27716 18617 27718
rect 25267 27770 25323 27772
rect 25347 27770 25403 27772
rect 25427 27770 25483 27772
rect 25507 27770 25563 27772
rect 25267 27718 25313 27770
rect 25313 27718 25323 27770
rect 25347 27718 25377 27770
rect 25377 27718 25389 27770
rect 25389 27718 25403 27770
rect 25427 27718 25441 27770
rect 25441 27718 25453 27770
rect 25453 27718 25483 27770
rect 25507 27718 25517 27770
rect 25517 27718 25563 27770
rect 25267 27716 25323 27718
rect 25347 27716 25403 27718
rect 25427 27716 25483 27718
rect 25507 27716 25563 27718
rect 28538 27532 28594 27568
rect 28538 27512 28540 27532
rect 28540 27512 28592 27532
rect 28592 27512 28594 27532
rect 7902 27226 7958 27228
rect 7982 27226 8038 27228
rect 8062 27226 8118 27228
rect 8142 27226 8198 27228
rect 7902 27174 7948 27226
rect 7948 27174 7958 27226
rect 7982 27174 8012 27226
rect 8012 27174 8024 27226
rect 8024 27174 8038 27226
rect 8062 27174 8076 27226
rect 8076 27174 8088 27226
rect 8088 27174 8118 27226
rect 8142 27174 8152 27226
rect 8152 27174 8198 27226
rect 7902 27172 7958 27174
rect 7982 27172 8038 27174
rect 8062 27172 8118 27174
rect 8142 27172 8198 27174
rect 14848 27226 14904 27228
rect 14928 27226 14984 27228
rect 15008 27226 15064 27228
rect 15088 27226 15144 27228
rect 14848 27174 14894 27226
rect 14894 27174 14904 27226
rect 14928 27174 14958 27226
rect 14958 27174 14970 27226
rect 14970 27174 14984 27226
rect 15008 27174 15022 27226
rect 15022 27174 15034 27226
rect 15034 27174 15064 27226
rect 15088 27174 15098 27226
rect 15098 27174 15144 27226
rect 14848 27172 14904 27174
rect 14928 27172 14984 27174
rect 15008 27172 15064 27174
rect 15088 27172 15144 27174
rect 21794 27226 21850 27228
rect 21874 27226 21930 27228
rect 21954 27226 22010 27228
rect 22034 27226 22090 27228
rect 21794 27174 21840 27226
rect 21840 27174 21850 27226
rect 21874 27174 21904 27226
rect 21904 27174 21916 27226
rect 21916 27174 21930 27226
rect 21954 27174 21968 27226
rect 21968 27174 21980 27226
rect 21980 27174 22010 27226
rect 22034 27174 22044 27226
rect 22044 27174 22090 27226
rect 21794 27172 21850 27174
rect 21874 27172 21930 27174
rect 21954 27172 22010 27174
rect 22034 27172 22090 27174
rect 28740 27226 28796 27228
rect 28820 27226 28876 27228
rect 28900 27226 28956 27228
rect 28980 27226 29036 27228
rect 28740 27174 28786 27226
rect 28786 27174 28796 27226
rect 28820 27174 28850 27226
rect 28850 27174 28862 27226
rect 28862 27174 28876 27226
rect 28900 27174 28914 27226
rect 28914 27174 28926 27226
rect 28926 27174 28956 27226
rect 28980 27174 28990 27226
rect 28990 27174 29036 27226
rect 28740 27172 28796 27174
rect 28820 27172 28876 27174
rect 28900 27172 28956 27174
rect 28980 27172 29036 27174
rect 4429 26682 4485 26684
rect 4509 26682 4565 26684
rect 4589 26682 4645 26684
rect 4669 26682 4725 26684
rect 4429 26630 4475 26682
rect 4475 26630 4485 26682
rect 4509 26630 4539 26682
rect 4539 26630 4551 26682
rect 4551 26630 4565 26682
rect 4589 26630 4603 26682
rect 4603 26630 4615 26682
rect 4615 26630 4645 26682
rect 4669 26630 4679 26682
rect 4679 26630 4725 26682
rect 4429 26628 4485 26630
rect 4509 26628 4565 26630
rect 4589 26628 4645 26630
rect 4669 26628 4725 26630
rect 11375 26682 11431 26684
rect 11455 26682 11511 26684
rect 11535 26682 11591 26684
rect 11615 26682 11671 26684
rect 11375 26630 11421 26682
rect 11421 26630 11431 26682
rect 11455 26630 11485 26682
rect 11485 26630 11497 26682
rect 11497 26630 11511 26682
rect 11535 26630 11549 26682
rect 11549 26630 11561 26682
rect 11561 26630 11591 26682
rect 11615 26630 11625 26682
rect 11625 26630 11671 26682
rect 11375 26628 11431 26630
rect 11455 26628 11511 26630
rect 11535 26628 11591 26630
rect 11615 26628 11671 26630
rect 18321 26682 18377 26684
rect 18401 26682 18457 26684
rect 18481 26682 18537 26684
rect 18561 26682 18617 26684
rect 18321 26630 18367 26682
rect 18367 26630 18377 26682
rect 18401 26630 18431 26682
rect 18431 26630 18443 26682
rect 18443 26630 18457 26682
rect 18481 26630 18495 26682
rect 18495 26630 18507 26682
rect 18507 26630 18537 26682
rect 18561 26630 18571 26682
rect 18571 26630 18617 26682
rect 18321 26628 18377 26630
rect 18401 26628 18457 26630
rect 18481 26628 18537 26630
rect 18561 26628 18617 26630
rect 7902 26138 7958 26140
rect 7982 26138 8038 26140
rect 8062 26138 8118 26140
rect 8142 26138 8198 26140
rect 7902 26086 7948 26138
rect 7948 26086 7958 26138
rect 7982 26086 8012 26138
rect 8012 26086 8024 26138
rect 8024 26086 8038 26138
rect 8062 26086 8076 26138
rect 8076 26086 8088 26138
rect 8088 26086 8118 26138
rect 8142 26086 8152 26138
rect 8152 26086 8198 26138
rect 7902 26084 7958 26086
rect 7982 26084 8038 26086
rect 8062 26084 8118 26086
rect 8142 26084 8198 26086
rect 4429 25594 4485 25596
rect 4509 25594 4565 25596
rect 4589 25594 4645 25596
rect 4669 25594 4725 25596
rect 4429 25542 4475 25594
rect 4475 25542 4485 25594
rect 4509 25542 4539 25594
rect 4539 25542 4551 25594
rect 4551 25542 4565 25594
rect 4589 25542 4603 25594
rect 4603 25542 4615 25594
rect 4615 25542 4645 25594
rect 4669 25542 4679 25594
rect 4679 25542 4725 25594
rect 4429 25540 4485 25542
rect 4509 25540 4565 25542
rect 4589 25540 4645 25542
rect 4669 25540 4725 25542
rect 11375 25594 11431 25596
rect 11455 25594 11511 25596
rect 11535 25594 11591 25596
rect 11615 25594 11671 25596
rect 11375 25542 11421 25594
rect 11421 25542 11431 25594
rect 11455 25542 11485 25594
rect 11485 25542 11497 25594
rect 11497 25542 11511 25594
rect 11535 25542 11549 25594
rect 11549 25542 11561 25594
rect 11561 25542 11591 25594
rect 11615 25542 11625 25594
rect 11625 25542 11671 25594
rect 11375 25540 11431 25542
rect 11455 25540 11511 25542
rect 11535 25540 11591 25542
rect 11615 25540 11671 25542
rect 7902 25050 7958 25052
rect 7982 25050 8038 25052
rect 8062 25050 8118 25052
rect 8142 25050 8198 25052
rect 7902 24998 7948 25050
rect 7948 24998 7958 25050
rect 7982 24998 8012 25050
rect 8012 24998 8024 25050
rect 8024 24998 8038 25050
rect 8062 24998 8076 25050
rect 8076 24998 8088 25050
rect 8088 24998 8118 25050
rect 8142 24998 8152 25050
rect 8152 24998 8198 25050
rect 7902 24996 7958 24998
rect 7982 24996 8038 24998
rect 8062 24996 8118 24998
rect 8142 24996 8198 24998
rect 4429 24506 4485 24508
rect 4509 24506 4565 24508
rect 4589 24506 4645 24508
rect 4669 24506 4725 24508
rect 4429 24454 4475 24506
rect 4475 24454 4485 24506
rect 4509 24454 4539 24506
rect 4539 24454 4551 24506
rect 4551 24454 4565 24506
rect 4589 24454 4603 24506
rect 4603 24454 4615 24506
rect 4615 24454 4645 24506
rect 4669 24454 4679 24506
rect 4679 24454 4725 24506
rect 4429 24452 4485 24454
rect 4509 24452 4565 24454
rect 4589 24452 4645 24454
rect 4669 24452 4725 24454
rect 11375 24506 11431 24508
rect 11455 24506 11511 24508
rect 11535 24506 11591 24508
rect 11615 24506 11671 24508
rect 11375 24454 11421 24506
rect 11421 24454 11431 24506
rect 11455 24454 11485 24506
rect 11485 24454 11497 24506
rect 11497 24454 11511 24506
rect 11535 24454 11549 24506
rect 11549 24454 11561 24506
rect 11561 24454 11591 24506
rect 11615 24454 11625 24506
rect 11625 24454 11671 24506
rect 11375 24452 11431 24454
rect 11455 24452 11511 24454
rect 11535 24452 11591 24454
rect 11615 24452 11671 24454
rect 7902 23962 7958 23964
rect 7982 23962 8038 23964
rect 8062 23962 8118 23964
rect 8142 23962 8198 23964
rect 7902 23910 7948 23962
rect 7948 23910 7958 23962
rect 7982 23910 8012 23962
rect 8012 23910 8024 23962
rect 8024 23910 8038 23962
rect 8062 23910 8076 23962
rect 8076 23910 8088 23962
rect 8088 23910 8118 23962
rect 8142 23910 8152 23962
rect 8152 23910 8198 23962
rect 7902 23908 7958 23910
rect 7982 23908 8038 23910
rect 8062 23908 8118 23910
rect 8142 23908 8198 23910
rect 1398 23432 1454 23488
rect 1030 22888 1086 22944
rect 938 22616 994 22672
rect 938 22344 994 22400
rect 1030 22072 1086 22128
rect 1030 21800 1086 21856
rect 938 21528 994 21584
rect 938 21256 994 21312
rect 1030 20984 1086 21040
rect 938 20712 994 20768
rect 1398 20576 1454 20632
rect 4429 23418 4485 23420
rect 4509 23418 4565 23420
rect 4589 23418 4645 23420
rect 4669 23418 4725 23420
rect 4429 23366 4475 23418
rect 4475 23366 4485 23418
rect 4509 23366 4539 23418
rect 4539 23366 4551 23418
rect 4551 23366 4565 23418
rect 4589 23366 4603 23418
rect 4603 23366 4615 23418
rect 4615 23366 4645 23418
rect 4669 23366 4679 23418
rect 4679 23366 4725 23418
rect 4429 23364 4485 23366
rect 4509 23364 4565 23366
rect 4589 23364 4645 23366
rect 4669 23364 4725 23366
rect 11375 23418 11431 23420
rect 11455 23418 11511 23420
rect 11535 23418 11591 23420
rect 11615 23418 11671 23420
rect 11375 23366 11421 23418
rect 11421 23366 11431 23418
rect 11455 23366 11485 23418
rect 11485 23366 11497 23418
rect 11497 23366 11511 23418
rect 11535 23366 11549 23418
rect 11549 23366 11561 23418
rect 11561 23366 11591 23418
rect 11615 23366 11625 23418
rect 11625 23366 11671 23418
rect 11375 23364 11431 23366
rect 11455 23364 11511 23366
rect 11535 23364 11591 23366
rect 11615 23364 11671 23366
rect 1030 20168 1086 20224
rect 938 19896 994 19952
rect 1030 19624 1086 19680
rect 938 19352 994 19408
rect 1398 18944 1454 19000
rect 1030 18536 1086 18592
rect 938 18264 994 18320
rect 938 17992 994 18048
rect 1398 17856 1454 17912
rect 938 17448 994 17504
rect 1030 17176 1086 17232
rect 938 16904 994 16960
rect 1030 16632 1086 16688
rect 938 16360 994 16416
rect 1030 16088 1086 16144
rect 938 15816 994 15872
rect 1030 15544 1086 15600
rect 938 15272 994 15328
rect 938 14456 994 14512
rect 938 14184 994 14240
rect 1030 13912 1086 13968
rect 938 13096 994 13152
rect 1030 12824 1086 12880
rect 938 12552 994 12608
rect 938 12008 994 12064
rect 1030 11736 1086 11792
rect 938 11464 994 11520
rect 1030 11192 1086 11248
rect 938 10376 994 10432
rect 1030 10104 1086 10160
rect 938 9832 994 9888
rect 938 9288 994 9344
rect 1030 9016 1086 9072
rect 938 8744 994 8800
rect 1030 8472 1086 8528
rect 1030 8372 1032 8392
rect 1032 8372 1084 8392
rect 1084 8372 1086 8392
rect 1030 8336 1086 8372
rect 938 7112 994 7168
rect 1674 19216 1730 19272
rect 1674 15272 1730 15328
rect 1858 15136 1914 15192
rect 1858 14320 1914 14376
rect 1858 13776 1914 13832
rect 1398 13640 1454 13696
rect 1674 13640 1730 13696
rect 1858 13404 1860 13424
rect 1860 13404 1912 13424
rect 1912 13404 1914 13424
rect 1858 13368 1914 13404
rect 1582 13232 1638 13288
rect 1858 12708 1914 12744
rect 1858 12688 1860 12708
rect 1860 12688 1912 12708
rect 1912 12688 1914 12708
rect 1674 12280 1730 12336
rect 1858 12144 1914 12200
rect 1398 10920 1454 10976
rect 1674 10920 1730 10976
rect 1582 10532 1638 10568
rect 1582 10512 1584 10532
rect 1584 10512 1636 10532
rect 1636 10512 1638 10532
rect 1674 9560 1730 9616
rect 1582 8744 1638 8800
rect 1398 8200 1454 8256
rect 1306 7112 1362 7168
rect 1306 6296 1362 6352
rect 1582 8472 1638 8528
rect 1674 8200 1730 8256
rect 1766 7656 1822 7712
rect 1490 6840 1546 6896
rect 1766 6840 1822 6896
rect 2134 8880 2190 8936
rect 2042 6568 2098 6624
rect 1950 5480 2006 5536
rect 2410 8608 2466 8664
rect 2502 7268 2558 7304
rect 2502 7248 2504 7268
rect 2504 7248 2556 7268
rect 2556 7248 2558 7268
rect 2410 5208 2466 5264
rect 2778 7656 2834 7712
rect 2778 7384 2834 7440
rect 2042 3440 2098 3496
rect 3054 7112 3110 7168
rect 2962 5480 3018 5536
rect 2870 3304 2926 3360
rect 3330 7656 3386 7712
rect 4066 18808 4122 18864
rect 7902 22874 7958 22876
rect 7982 22874 8038 22876
rect 8062 22874 8118 22876
rect 8142 22874 8198 22876
rect 7902 22822 7948 22874
rect 7948 22822 7958 22874
rect 7982 22822 8012 22874
rect 8012 22822 8024 22874
rect 8024 22822 8038 22874
rect 8062 22822 8076 22874
rect 8076 22822 8088 22874
rect 8088 22822 8118 22874
rect 8142 22822 8152 22874
rect 8152 22822 8198 22874
rect 7902 22820 7958 22822
rect 7982 22820 8038 22822
rect 8062 22820 8118 22822
rect 8142 22820 8198 22822
rect 4429 22330 4485 22332
rect 4509 22330 4565 22332
rect 4589 22330 4645 22332
rect 4669 22330 4725 22332
rect 4429 22278 4475 22330
rect 4475 22278 4485 22330
rect 4509 22278 4539 22330
rect 4539 22278 4551 22330
rect 4551 22278 4565 22330
rect 4589 22278 4603 22330
rect 4603 22278 4615 22330
rect 4615 22278 4645 22330
rect 4669 22278 4679 22330
rect 4679 22278 4725 22330
rect 4429 22276 4485 22278
rect 4509 22276 4565 22278
rect 4589 22276 4645 22278
rect 4669 22276 4725 22278
rect 7902 21786 7958 21788
rect 7982 21786 8038 21788
rect 8062 21786 8118 21788
rect 8142 21786 8198 21788
rect 7902 21734 7948 21786
rect 7948 21734 7958 21786
rect 7982 21734 8012 21786
rect 8012 21734 8024 21786
rect 8024 21734 8038 21786
rect 8062 21734 8076 21786
rect 8076 21734 8088 21786
rect 8088 21734 8118 21786
rect 8142 21734 8152 21786
rect 8152 21734 8198 21786
rect 7902 21732 7958 21734
rect 7982 21732 8038 21734
rect 8062 21732 8118 21734
rect 8142 21732 8198 21734
rect 4429 21242 4485 21244
rect 4509 21242 4565 21244
rect 4589 21242 4645 21244
rect 4669 21242 4725 21244
rect 4429 21190 4475 21242
rect 4475 21190 4485 21242
rect 4509 21190 4539 21242
rect 4539 21190 4551 21242
rect 4551 21190 4565 21242
rect 4589 21190 4603 21242
rect 4603 21190 4615 21242
rect 4615 21190 4645 21242
rect 4669 21190 4679 21242
rect 4679 21190 4725 21242
rect 4429 21188 4485 21190
rect 4509 21188 4565 21190
rect 4589 21188 4645 21190
rect 4669 21188 4725 21190
rect 4429 20154 4485 20156
rect 4509 20154 4565 20156
rect 4589 20154 4645 20156
rect 4669 20154 4725 20156
rect 4429 20102 4475 20154
rect 4475 20102 4485 20154
rect 4509 20102 4539 20154
rect 4539 20102 4551 20154
rect 4551 20102 4565 20154
rect 4589 20102 4603 20154
rect 4603 20102 4615 20154
rect 4615 20102 4645 20154
rect 4669 20102 4679 20154
rect 4679 20102 4725 20154
rect 4429 20100 4485 20102
rect 4509 20100 4565 20102
rect 4589 20100 4645 20102
rect 4669 20100 4725 20102
rect 4429 19066 4485 19068
rect 4509 19066 4565 19068
rect 4589 19066 4645 19068
rect 4669 19066 4725 19068
rect 4429 19014 4475 19066
rect 4475 19014 4485 19066
rect 4509 19014 4539 19066
rect 4539 19014 4551 19066
rect 4551 19014 4565 19066
rect 4589 19014 4603 19066
rect 4603 19014 4615 19066
rect 4615 19014 4645 19066
rect 4669 19014 4679 19066
rect 4679 19014 4725 19066
rect 4429 19012 4485 19014
rect 4509 19012 4565 19014
rect 4589 19012 4645 19014
rect 4669 19012 4725 19014
rect 4429 17978 4485 17980
rect 4509 17978 4565 17980
rect 4589 17978 4645 17980
rect 4669 17978 4725 17980
rect 4429 17926 4475 17978
rect 4475 17926 4485 17978
rect 4509 17926 4539 17978
rect 4539 17926 4551 17978
rect 4551 17926 4565 17978
rect 4589 17926 4603 17978
rect 4603 17926 4615 17978
rect 4615 17926 4645 17978
rect 4669 17926 4679 17978
rect 4679 17926 4725 17978
rect 4429 17924 4485 17926
rect 4509 17924 4565 17926
rect 4589 17924 4645 17926
rect 4669 17924 4725 17926
rect 4429 16890 4485 16892
rect 4509 16890 4565 16892
rect 4589 16890 4645 16892
rect 4669 16890 4725 16892
rect 4429 16838 4475 16890
rect 4475 16838 4485 16890
rect 4509 16838 4539 16890
rect 4539 16838 4551 16890
rect 4551 16838 4565 16890
rect 4589 16838 4603 16890
rect 4603 16838 4615 16890
rect 4615 16838 4645 16890
rect 4669 16838 4679 16890
rect 4679 16838 4725 16890
rect 4429 16836 4485 16838
rect 4509 16836 4565 16838
rect 4589 16836 4645 16838
rect 4669 16836 4725 16838
rect 4429 15802 4485 15804
rect 4509 15802 4565 15804
rect 4589 15802 4645 15804
rect 4669 15802 4725 15804
rect 4429 15750 4475 15802
rect 4475 15750 4485 15802
rect 4509 15750 4539 15802
rect 4539 15750 4551 15802
rect 4551 15750 4565 15802
rect 4589 15750 4603 15802
rect 4603 15750 4615 15802
rect 4615 15750 4645 15802
rect 4669 15750 4679 15802
rect 4679 15750 4725 15802
rect 4429 15748 4485 15750
rect 4509 15748 4565 15750
rect 4589 15748 4645 15750
rect 4669 15748 4725 15750
rect 4429 14714 4485 14716
rect 4509 14714 4565 14716
rect 4589 14714 4645 14716
rect 4669 14714 4725 14716
rect 4429 14662 4475 14714
rect 4475 14662 4485 14714
rect 4509 14662 4539 14714
rect 4539 14662 4551 14714
rect 4551 14662 4565 14714
rect 4589 14662 4603 14714
rect 4603 14662 4615 14714
rect 4615 14662 4645 14714
rect 4669 14662 4679 14714
rect 4679 14662 4725 14714
rect 4429 14660 4485 14662
rect 4509 14660 4565 14662
rect 4589 14660 4645 14662
rect 4669 14660 4725 14662
rect 4429 13626 4485 13628
rect 4509 13626 4565 13628
rect 4589 13626 4645 13628
rect 4669 13626 4725 13628
rect 4429 13574 4475 13626
rect 4475 13574 4485 13626
rect 4509 13574 4539 13626
rect 4539 13574 4551 13626
rect 4551 13574 4565 13626
rect 4589 13574 4603 13626
rect 4603 13574 4615 13626
rect 4615 13574 4645 13626
rect 4669 13574 4679 13626
rect 4679 13574 4725 13626
rect 4429 13572 4485 13574
rect 4509 13572 4565 13574
rect 4589 13572 4645 13574
rect 4669 13572 4725 13574
rect 4429 12538 4485 12540
rect 4509 12538 4565 12540
rect 4589 12538 4645 12540
rect 4669 12538 4725 12540
rect 4429 12486 4475 12538
rect 4475 12486 4485 12538
rect 4509 12486 4539 12538
rect 4539 12486 4551 12538
rect 4551 12486 4565 12538
rect 4589 12486 4603 12538
rect 4603 12486 4615 12538
rect 4615 12486 4645 12538
rect 4669 12486 4679 12538
rect 4679 12486 4725 12538
rect 4429 12484 4485 12486
rect 4509 12484 4565 12486
rect 4589 12484 4645 12486
rect 4669 12484 4725 12486
rect 5170 11736 5226 11792
rect 4429 11450 4485 11452
rect 4509 11450 4565 11452
rect 4589 11450 4645 11452
rect 4669 11450 4725 11452
rect 4429 11398 4475 11450
rect 4475 11398 4485 11450
rect 4509 11398 4539 11450
rect 4539 11398 4551 11450
rect 4551 11398 4565 11450
rect 4589 11398 4603 11450
rect 4603 11398 4615 11450
rect 4615 11398 4645 11450
rect 4669 11398 4679 11450
rect 4679 11398 4725 11450
rect 4429 11396 4485 11398
rect 4509 11396 4565 11398
rect 4589 11396 4645 11398
rect 4669 11396 4725 11398
rect 4066 4664 4122 4720
rect 4429 10362 4485 10364
rect 4509 10362 4565 10364
rect 4589 10362 4645 10364
rect 4669 10362 4725 10364
rect 4429 10310 4475 10362
rect 4475 10310 4485 10362
rect 4509 10310 4539 10362
rect 4539 10310 4551 10362
rect 4551 10310 4565 10362
rect 4589 10310 4603 10362
rect 4603 10310 4615 10362
rect 4615 10310 4645 10362
rect 4669 10310 4679 10362
rect 4679 10310 4725 10362
rect 4429 10308 4485 10310
rect 4509 10308 4565 10310
rect 4589 10308 4645 10310
rect 4669 10308 4725 10310
rect 4802 9968 4858 10024
rect 4618 9596 4620 9616
rect 4620 9596 4672 9616
rect 4672 9596 4674 9616
rect 4618 9560 4674 9596
rect 4429 9274 4485 9276
rect 4509 9274 4565 9276
rect 4589 9274 4645 9276
rect 4669 9274 4725 9276
rect 4429 9222 4475 9274
rect 4475 9222 4485 9274
rect 4509 9222 4539 9274
rect 4539 9222 4551 9274
rect 4551 9222 4565 9274
rect 4589 9222 4603 9274
rect 4603 9222 4615 9274
rect 4615 9222 4645 9274
rect 4669 9222 4679 9274
rect 4679 9222 4725 9274
rect 4429 9220 4485 9222
rect 4509 9220 4565 9222
rect 4589 9220 4645 9222
rect 4669 9220 4725 9222
rect 4429 8186 4485 8188
rect 4509 8186 4565 8188
rect 4589 8186 4645 8188
rect 4669 8186 4725 8188
rect 4429 8134 4475 8186
rect 4475 8134 4485 8186
rect 4509 8134 4539 8186
rect 4539 8134 4551 8186
rect 4551 8134 4565 8186
rect 4589 8134 4603 8186
rect 4603 8134 4615 8186
rect 4615 8134 4645 8186
rect 4669 8134 4679 8186
rect 4679 8134 4725 8186
rect 4429 8132 4485 8134
rect 4509 8132 4565 8134
rect 4589 8132 4645 8134
rect 4669 8132 4725 8134
rect 4429 7098 4485 7100
rect 4509 7098 4565 7100
rect 4589 7098 4645 7100
rect 4669 7098 4725 7100
rect 4429 7046 4475 7098
rect 4475 7046 4485 7098
rect 4509 7046 4539 7098
rect 4539 7046 4551 7098
rect 4551 7046 4565 7098
rect 4589 7046 4603 7098
rect 4603 7046 4615 7098
rect 4615 7046 4645 7098
rect 4669 7046 4679 7098
rect 4679 7046 4725 7098
rect 4429 7044 4485 7046
rect 4509 7044 4565 7046
rect 4589 7044 4645 7046
rect 4669 7044 4725 7046
rect 4429 6010 4485 6012
rect 4509 6010 4565 6012
rect 4589 6010 4645 6012
rect 4669 6010 4725 6012
rect 4429 5958 4475 6010
rect 4475 5958 4485 6010
rect 4509 5958 4539 6010
rect 4539 5958 4551 6010
rect 4551 5958 4565 6010
rect 4589 5958 4603 6010
rect 4603 5958 4615 6010
rect 4615 5958 4645 6010
rect 4669 5958 4679 6010
rect 4679 5958 4725 6010
rect 4429 5956 4485 5958
rect 4509 5956 4565 5958
rect 4589 5956 4645 5958
rect 4669 5956 4725 5958
rect 5078 9580 5134 9616
rect 5078 9560 5080 9580
rect 5080 9560 5132 9580
rect 5132 9560 5134 9580
rect 7902 20698 7958 20700
rect 7982 20698 8038 20700
rect 8062 20698 8118 20700
rect 8142 20698 8198 20700
rect 7902 20646 7948 20698
rect 7948 20646 7958 20698
rect 7982 20646 8012 20698
rect 8012 20646 8024 20698
rect 8024 20646 8038 20698
rect 8062 20646 8076 20698
rect 8076 20646 8088 20698
rect 8088 20646 8118 20698
rect 8142 20646 8152 20698
rect 8152 20646 8198 20698
rect 7902 20644 7958 20646
rect 7982 20644 8038 20646
rect 8062 20644 8118 20646
rect 8142 20644 8198 20646
rect 7902 19610 7958 19612
rect 7982 19610 8038 19612
rect 8062 19610 8118 19612
rect 8142 19610 8198 19612
rect 7902 19558 7948 19610
rect 7948 19558 7958 19610
rect 7982 19558 8012 19610
rect 8012 19558 8024 19610
rect 8024 19558 8038 19610
rect 8062 19558 8076 19610
rect 8076 19558 8088 19610
rect 8088 19558 8118 19610
rect 8142 19558 8152 19610
rect 8152 19558 8198 19610
rect 7902 19556 7958 19558
rect 7982 19556 8038 19558
rect 8062 19556 8118 19558
rect 8142 19556 8198 19558
rect 7902 18522 7958 18524
rect 7982 18522 8038 18524
rect 8062 18522 8118 18524
rect 8142 18522 8198 18524
rect 7902 18470 7948 18522
rect 7948 18470 7958 18522
rect 7982 18470 8012 18522
rect 8012 18470 8024 18522
rect 8024 18470 8038 18522
rect 8062 18470 8076 18522
rect 8076 18470 8088 18522
rect 8088 18470 8118 18522
rect 8142 18470 8152 18522
rect 8152 18470 8198 18522
rect 7902 18468 7958 18470
rect 7982 18468 8038 18470
rect 8062 18468 8118 18470
rect 8142 18468 8198 18470
rect 7902 17434 7958 17436
rect 7982 17434 8038 17436
rect 8062 17434 8118 17436
rect 8142 17434 8198 17436
rect 7902 17382 7948 17434
rect 7948 17382 7958 17434
rect 7982 17382 8012 17434
rect 8012 17382 8024 17434
rect 8024 17382 8038 17434
rect 8062 17382 8076 17434
rect 8076 17382 8088 17434
rect 8088 17382 8118 17434
rect 8142 17382 8152 17434
rect 8152 17382 8198 17434
rect 7902 17380 7958 17382
rect 7982 17380 8038 17382
rect 8062 17380 8118 17382
rect 8142 17380 8198 17382
rect 5722 9988 5778 10024
rect 5722 9968 5724 9988
rect 5724 9968 5776 9988
rect 5776 9968 5778 9988
rect 5354 9152 5410 9208
rect 4429 4922 4485 4924
rect 4509 4922 4565 4924
rect 4589 4922 4645 4924
rect 4669 4922 4725 4924
rect 4429 4870 4475 4922
rect 4475 4870 4485 4922
rect 4509 4870 4539 4922
rect 4539 4870 4551 4922
rect 4551 4870 4565 4922
rect 4589 4870 4603 4922
rect 4603 4870 4615 4922
rect 4615 4870 4645 4922
rect 4669 4870 4679 4922
rect 4679 4870 4725 4922
rect 4429 4868 4485 4870
rect 4509 4868 4565 4870
rect 4589 4868 4645 4870
rect 4669 4868 4725 4870
rect 4802 3984 4858 4040
rect 4429 3834 4485 3836
rect 4509 3834 4565 3836
rect 4589 3834 4645 3836
rect 4669 3834 4725 3836
rect 4429 3782 4475 3834
rect 4475 3782 4485 3834
rect 4509 3782 4539 3834
rect 4539 3782 4551 3834
rect 4551 3782 4565 3834
rect 4589 3782 4603 3834
rect 4603 3782 4615 3834
rect 4615 3782 4645 3834
rect 4669 3782 4679 3834
rect 4679 3782 4725 3834
rect 4429 3780 4485 3782
rect 4509 3780 4565 3782
rect 4589 3780 4645 3782
rect 4669 3780 4725 3782
rect 6274 6704 6330 6760
rect 6090 5208 6146 5264
rect 5078 3440 5134 3496
rect 4526 3304 4582 3360
rect 4429 2746 4485 2748
rect 4509 2746 4565 2748
rect 4589 2746 4645 2748
rect 4669 2746 4725 2748
rect 4429 2694 4475 2746
rect 4475 2694 4485 2746
rect 4509 2694 4539 2746
rect 4539 2694 4551 2746
rect 4551 2694 4565 2746
rect 4589 2694 4603 2746
rect 4603 2694 4615 2746
rect 4615 2694 4645 2746
rect 4669 2694 4679 2746
rect 4679 2694 4725 2746
rect 4429 2692 4485 2694
rect 4509 2692 4565 2694
rect 4589 2692 4645 2694
rect 4669 2692 4725 2694
rect 6642 8744 6698 8800
rect 6550 8336 6606 8392
rect 7010 7112 7066 7168
rect 6918 6840 6974 6896
rect 6550 5072 6606 5128
rect 7902 16346 7958 16348
rect 7982 16346 8038 16348
rect 8062 16346 8118 16348
rect 8142 16346 8198 16348
rect 7902 16294 7948 16346
rect 7948 16294 7958 16346
rect 7982 16294 8012 16346
rect 8012 16294 8024 16346
rect 8024 16294 8038 16346
rect 8062 16294 8076 16346
rect 8076 16294 8088 16346
rect 8088 16294 8118 16346
rect 8142 16294 8152 16346
rect 8152 16294 8198 16346
rect 7902 16292 7958 16294
rect 7982 16292 8038 16294
rect 8062 16292 8118 16294
rect 8142 16292 8198 16294
rect 7902 15258 7958 15260
rect 7982 15258 8038 15260
rect 8062 15258 8118 15260
rect 8142 15258 8198 15260
rect 7902 15206 7948 15258
rect 7948 15206 7958 15258
rect 7982 15206 8012 15258
rect 8012 15206 8024 15258
rect 8024 15206 8038 15258
rect 8062 15206 8076 15258
rect 8076 15206 8088 15258
rect 8088 15206 8118 15258
rect 8142 15206 8152 15258
rect 8152 15206 8198 15258
rect 7902 15204 7958 15206
rect 7982 15204 8038 15206
rect 8062 15204 8118 15206
rect 8142 15204 8198 15206
rect 7902 14170 7958 14172
rect 7982 14170 8038 14172
rect 8062 14170 8118 14172
rect 8142 14170 8198 14172
rect 7902 14118 7948 14170
rect 7948 14118 7958 14170
rect 7982 14118 8012 14170
rect 8012 14118 8024 14170
rect 8024 14118 8038 14170
rect 8062 14118 8076 14170
rect 8076 14118 8088 14170
rect 8088 14118 8118 14170
rect 8142 14118 8152 14170
rect 8152 14118 8198 14170
rect 7902 14116 7958 14118
rect 7982 14116 8038 14118
rect 8062 14116 8118 14118
rect 8142 14116 8198 14118
rect 8390 13640 8446 13696
rect 7902 13082 7958 13084
rect 7982 13082 8038 13084
rect 8062 13082 8118 13084
rect 8142 13082 8198 13084
rect 7902 13030 7948 13082
rect 7948 13030 7958 13082
rect 7982 13030 8012 13082
rect 8012 13030 8024 13082
rect 8024 13030 8038 13082
rect 8062 13030 8076 13082
rect 8076 13030 8088 13082
rect 8088 13030 8118 13082
rect 8142 13030 8152 13082
rect 8152 13030 8198 13082
rect 7902 13028 7958 13030
rect 7982 13028 8038 13030
rect 8062 13028 8118 13030
rect 8142 13028 8198 13030
rect 8022 12844 8078 12880
rect 8022 12824 8024 12844
rect 8024 12824 8076 12844
rect 8076 12824 8078 12844
rect 7930 12416 7986 12472
rect 7902 11994 7958 11996
rect 7982 11994 8038 11996
rect 8062 11994 8118 11996
rect 8142 11994 8198 11996
rect 7902 11942 7948 11994
rect 7948 11942 7958 11994
rect 7982 11942 8012 11994
rect 8012 11942 8024 11994
rect 8024 11942 8038 11994
rect 8062 11942 8076 11994
rect 8076 11942 8088 11994
rect 8088 11942 8118 11994
rect 8142 11942 8152 11994
rect 8152 11942 8198 11994
rect 7902 11940 7958 11942
rect 7982 11940 8038 11942
rect 8062 11940 8118 11942
rect 8142 11940 8198 11942
rect 7930 11736 7986 11792
rect 7902 10906 7958 10908
rect 7982 10906 8038 10908
rect 8062 10906 8118 10908
rect 8142 10906 8198 10908
rect 7902 10854 7948 10906
rect 7948 10854 7958 10906
rect 7982 10854 8012 10906
rect 8012 10854 8024 10906
rect 8024 10854 8038 10906
rect 8062 10854 8076 10906
rect 8076 10854 8088 10906
rect 8088 10854 8118 10906
rect 8142 10854 8152 10906
rect 8152 10854 8198 10906
rect 7902 10852 7958 10854
rect 7982 10852 8038 10854
rect 8062 10852 8118 10854
rect 8142 10852 8198 10854
rect 7902 9818 7958 9820
rect 7982 9818 8038 9820
rect 8062 9818 8118 9820
rect 8142 9818 8198 9820
rect 7902 9766 7948 9818
rect 7948 9766 7958 9818
rect 7982 9766 8012 9818
rect 8012 9766 8024 9818
rect 8024 9766 8038 9818
rect 8062 9766 8076 9818
rect 8076 9766 8088 9818
rect 8088 9766 8118 9818
rect 8142 9766 8152 9818
rect 8152 9766 8198 9818
rect 7902 9764 7958 9766
rect 7982 9764 8038 9766
rect 8062 9764 8118 9766
rect 8142 9764 8198 9766
rect 6734 2916 6790 2952
rect 6734 2896 6736 2916
rect 6736 2896 6788 2916
rect 6788 2896 6790 2916
rect 7562 8608 7618 8664
rect 7902 8730 7958 8732
rect 7982 8730 8038 8732
rect 8062 8730 8118 8732
rect 8142 8730 8198 8732
rect 7902 8678 7948 8730
rect 7948 8678 7958 8730
rect 7982 8678 8012 8730
rect 8012 8678 8024 8730
rect 8024 8678 8038 8730
rect 8062 8678 8076 8730
rect 8076 8678 8088 8730
rect 8088 8678 8118 8730
rect 8142 8678 8152 8730
rect 8152 8678 8198 8730
rect 7902 8676 7958 8678
rect 7982 8676 8038 8678
rect 8062 8676 8118 8678
rect 8142 8676 8198 8678
rect 8298 8472 8354 8528
rect 7902 7642 7958 7644
rect 7982 7642 8038 7644
rect 8062 7642 8118 7644
rect 8142 7642 8198 7644
rect 7902 7590 7948 7642
rect 7948 7590 7958 7642
rect 7982 7590 8012 7642
rect 8012 7590 8024 7642
rect 8024 7590 8038 7642
rect 8062 7590 8076 7642
rect 8076 7590 8088 7642
rect 8088 7590 8118 7642
rect 8142 7590 8152 7642
rect 8152 7590 8198 7642
rect 7902 7588 7958 7590
rect 7982 7588 8038 7590
rect 8062 7588 8118 7590
rect 8142 7588 8198 7590
rect 8482 8880 8538 8936
rect 7838 7112 7894 7168
rect 8114 6740 8116 6760
rect 8116 6740 8168 6760
rect 8168 6740 8170 6760
rect 8114 6704 8170 6740
rect 7902 6554 7958 6556
rect 7982 6554 8038 6556
rect 8062 6554 8118 6556
rect 8142 6554 8198 6556
rect 7902 6502 7948 6554
rect 7948 6502 7958 6554
rect 7982 6502 8012 6554
rect 8012 6502 8024 6554
rect 8024 6502 8038 6554
rect 8062 6502 8076 6554
rect 8076 6502 8088 6554
rect 8088 6502 8118 6554
rect 8142 6502 8152 6554
rect 8152 6502 8198 6554
rect 7902 6500 7958 6502
rect 7982 6500 8038 6502
rect 8062 6500 8118 6502
rect 8142 6500 8198 6502
rect 8758 12416 8814 12472
rect 8850 11328 8906 11384
rect 8666 6860 8722 6896
rect 8666 6840 8668 6860
rect 8668 6840 8720 6860
rect 8720 6840 8722 6860
rect 7378 4936 7434 4992
rect 7902 5466 7958 5468
rect 7982 5466 8038 5468
rect 8062 5466 8118 5468
rect 8142 5466 8198 5468
rect 7902 5414 7948 5466
rect 7948 5414 7958 5466
rect 7982 5414 8012 5466
rect 8012 5414 8024 5466
rect 8024 5414 8038 5466
rect 8062 5414 8076 5466
rect 8076 5414 8088 5466
rect 8088 5414 8118 5466
rect 8142 5414 8152 5466
rect 8152 5414 8198 5466
rect 7902 5412 7958 5414
rect 7982 5412 8038 5414
rect 8062 5412 8118 5414
rect 8142 5412 8198 5414
rect 8114 5208 8170 5264
rect 8206 4972 8208 4992
rect 8208 4972 8260 4992
rect 8260 4972 8262 4992
rect 8206 4936 8262 4972
rect 8114 4664 8170 4720
rect 7902 4378 7958 4380
rect 7982 4378 8038 4380
rect 8062 4378 8118 4380
rect 8142 4378 8198 4380
rect 7902 4326 7948 4378
rect 7948 4326 7958 4378
rect 7982 4326 8012 4378
rect 8012 4326 8024 4378
rect 8024 4326 8038 4378
rect 8062 4326 8076 4378
rect 8076 4326 8088 4378
rect 8088 4326 8118 4378
rect 8142 4326 8152 4378
rect 8152 4326 8198 4378
rect 7902 4324 7958 4326
rect 7982 4324 8038 4326
rect 8062 4324 8118 4326
rect 8142 4324 8198 4326
rect 7902 3290 7958 3292
rect 7982 3290 8038 3292
rect 8062 3290 8118 3292
rect 8142 3290 8198 3292
rect 7902 3238 7948 3290
rect 7948 3238 7958 3290
rect 7982 3238 8012 3290
rect 8012 3238 8024 3290
rect 8024 3238 8038 3290
rect 8062 3238 8076 3290
rect 8076 3238 8088 3290
rect 8088 3238 8118 3290
rect 8142 3238 8152 3290
rect 8152 3238 8198 3290
rect 7902 3236 7958 3238
rect 7982 3236 8038 3238
rect 8062 3236 8118 3238
rect 8142 3236 8198 3238
rect 8574 3984 8630 4040
rect 7902 2202 7958 2204
rect 7982 2202 8038 2204
rect 8062 2202 8118 2204
rect 8142 2202 8198 2204
rect 7902 2150 7948 2202
rect 7948 2150 7958 2202
rect 7982 2150 8012 2202
rect 8012 2150 8024 2202
rect 8024 2150 8038 2202
rect 8062 2150 8076 2202
rect 8076 2150 8088 2202
rect 8088 2150 8118 2202
rect 8142 2150 8152 2202
rect 8152 2150 8198 2202
rect 7902 2148 7958 2150
rect 7982 2148 8038 2150
rect 8062 2148 8118 2150
rect 8142 2148 8198 2150
rect 9586 12824 9642 12880
rect 9770 12280 9826 12336
rect 9586 11328 9642 11384
rect 10046 14456 10102 14512
rect 11375 22330 11431 22332
rect 11455 22330 11511 22332
rect 11535 22330 11591 22332
rect 11615 22330 11671 22332
rect 11375 22278 11421 22330
rect 11421 22278 11431 22330
rect 11455 22278 11485 22330
rect 11485 22278 11497 22330
rect 11497 22278 11511 22330
rect 11535 22278 11549 22330
rect 11549 22278 11561 22330
rect 11561 22278 11591 22330
rect 11615 22278 11625 22330
rect 11625 22278 11671 22330
rect 11375 22276 11431 22278
rect 11455 22276 11511 22278
rect 11535 22276 11591 22278
rect 11615 22276 11671 22278
rect 11375 21242 11431 21244
rect 11455 21242 11511 21244
rect 11535 21242 11591 21244
rect 11615 21242 11671 21244
rect 11375 21190 11421 21242
rect 11421 21190 11431 21242
rect 11455 21190 11485 21242
rect 11485 21190 11497 21242
rect 11497 21190 11511 21242
rect 11535 21190 11549 21242
rect 11549 21190 11561 21242
rect 11561 21190 11591 21242
rect 11615 21190 11625 21242
rect 11625 21190 11671 21242
rect 11375 21188 11431 21190
rect 11455 21188 11511 21190
rect 11535 21188 11591 21190
rect 11615 21188 11671 21190
rect 11375 20154 11431 20156
rect 11455 20154 11511 20156
rect 11535 20154 11591 20156
rect 11615 20154 11671 20156
rect 11375 20102 11421 20154
rect 11421 20102 11431 20154
rect 11455 20102 11485 20154
rect 11485 20102 11497 20154
rect 11497 20102 11511 20154
rect 11535 20102 11549 20154
rect 11549 20102 11561 20154
rect 11561 20102 11591 20154
rect 11615 20102 11625 20154
rect 11625 20102 11671 20154
rect 11375 20100 11431 20102
rect 11455 20100 11511 20102
rect 11535 20100 11591 20102
rect 11615 20100 11671 20102
rect 11375 19066 11431 19068
rect 11455 19066 11511 19068
rect 11535 19066 11591 19068
rect 11615 19066 11671 19068
rect 11375 19014 11421 19066
rect 11421 19014 11431 19066
rect 11455 19014 11485 19066
rect 11485 19014 11497 19066
rect 11497 19014 11511 19066
rect 11535 19014 11549 19066
rect 11549 19014 11561 19066
rect 11561 19014 11591 19066
rect 11615 19014 11625 19066
rect 11625 19014 11671 19066
rect 11375 19012 11431 19014
rect 11455 19012 11511 19014
rect 11535 19012 11591 19014
rect 11615 19012 11671 19014
rect 11375 17978 11431 17980
rect 11455 17978 11511 17980
rect 11535 17978 11591 17980
rect 11615 17978 11671 17980
rect 11375 17926 11421 17978
rect 11421 17926 11431 17978
rect 11455 17926 11485 17978
rect 11485 17926 11497 17978
rect 11497 17926 11511 17978
rect 11535 17926 11549 17978
rect 11549 17926 11561 17978
rect 11561 17926 11591 17978
rect 11615 17926 11625 17978
rect 11625 17926 11671 17978
rect 11375 17924 11431 17926
rect 11455 17924 11511 17926
rect 11535 17924 11591 17926
rect 11615 17924 11671 17926
rect 11375 16890 11431 16892
rect 11455 16890 11511 16892
rect 11535 16890 11591 16892
rect 11615 16890 11671 16892
rect 11375 16838 11421 16890
rect 11421 16838 11431 16890
rect 11455 16838 11485 16890
rect 11485 16838 11497 16890
rect 11497 16838 11511 16890
rect 11535 16838 11549 16890
rect 11549 16838 11561 16890
rect 11561 16838 11591 16890
rect 11615 16838 11625 16890
rect 11625 16838 11671 16890
rect 11375 16836 11431 16838
rect 11455 16836 11511 16838
rect 11535 16836 11591 16838
rect 11615 16836 11671 16838
rect 11375 15802 11431 15804
rect 11455 15802 11511 15804
rect 11535 15802 11591 15804
rect 11615 15802 11671 15804
rect 11375 15750 11421 15802
rect 11421 15750 11431 15802
rect 11455 15750 11485 15802
rect 11485 15750 11497 15802
rect 11497 15750 11511 15802
rect 11535 15750 11549 15802
rect 11549 15750 11561 15802
rect 11561 15750 11591 15802
rect 11615 15750 11625 15802
rect 11625 15750 11671 15802
rect 11375 15748 11431 15750
rect 11455 15748 11511 15750
rect 11535 15748 11591 15750
rect 11615 15748 11671 15750
rect 8758 4256 8814 4312
rect 10046 9444 10102 9480
rect 10046 9424 10048 9444
rect 10048 9424 10100 9444
rect 10100 9424 10102 9444
rect 9770 9016 9826 9072
rect 9770 7384 9826 7440
rect 9310 4140 9366 4176
rect 9310 4120 9312 4140
rect 9312 4120 9364 4140
rect 9364 4120 9366 4140
rect 9862 4256 9918 4312
rect 9586 3576 9642 3632
rect 11375 14714 11431 14716
rect 11455 14714 11511 14716
rect 11535 14714 11591 14716
rect 11615 14714 11671 14716
rect 11375 14662 11421 14714
rect 11421 14662 11431 14714
rect 11455 14662 11485 14714
rect 11485 14662 11497 14714
rect 11497 14662 11511 14714
rect 11535 14662 11549 14714
rect 11549 14662 11561 14714
rect 11561 14662 11591 14714
rect 11615 14662 11625 14714
rect 11625 14662 11671 14714
rect 11375 14660 11431 14662
rect 11455 14660 11511 14662
rect 11535 14660 11591 14662
rect 11615 14660 11671 14662
rect 10414 9560 10470 9616
rect 10506 9460 10508 9480
rect 10508 9460 10560 9480
rect 10560 9460 10562 9480
rect 10506 9424 10562 9460
rect 10598 9016 10654 9072
rect 10138 3712 10194 3768
rect 10782 6840 10838 6896
rect 10598 3984 10654 4040
rect 10782 3712 10838 3768
rect 11375 13626 11431 13628
rect 11455 13626 11511 13628
rect 11535 13626 11591 13628
rect 11615 13626 11671 13628
rect 11375 13574 11421 13626
rect 11421 13574 11431 13626
rect 11455 13574 11485 13626
rect 11485 13574 11497 13626
rect 11497 13574 11511 13626
rect 11535 13574 11549 13626
rect 11549 13574 11561 13626
rect 11561 13574 11591 13626
rect 11615 13574 11625 13626
rect 11625 13574 11671 13626
rect 11375 13572 11431 13574
rect 11455 13572 11511 13574
rect 11535 13572 11591 13574
rect 11615 13572 11671 13574
rect 14848 26138 14904 26140
rect 14928 26138 14984 26140
rect 15008 26138 15064 26140
rect 15088 26138 15144 26140
rect 14848 26086 14894 26138
rect 14894 26086 14904 26138
rect 14928 26086 14958 26138
rect 14958 26086 14970 26138
rect 14970 26086 14984 26138
rect 15008 26086 15022 26138
rect 15022 26086 15034 26138
rect 15034 26086 15064 26138
rect 15088 26086 15098 26138
rect 15098 26086 15144 26138
rect 14848 26084 14904 26086
rect 14928 26084 14984 26086
rect 15008 26084 15064 26086
rect 15088 26084 15144 26086
rect 21794 26138 21850 26140
rect 21874 26138 21930 26140
rect 21954 26138 22010 26140
rect 22034 26138 22090 26140
rect 21794 26086 21840 26138
rect 21840 26086 21850 26138
rect 21874 26086 21904 26138
rect 21904 26086 21916 26138
rect 21916 26086 21930 26138
rect 21954 26086 21968 26138
rect 21968 26086 21980 26138
rect 21980 26086 22010 26138
rect 22034 26086 22044 26138
rect 22044 26086 22090 26138
rect 21794 26084 21850 26086
rect 21874 26084 21930 26086
rect 21954 26084 22010 26086
rect 22034 26084 22090 26086
rect 18321 25594 18377 25596
rect 18401 25594 18457 25596
rect 18481 25594 18537 25596
rect 18561 25594 18617 25596
rect 18321 25542 18367 25594
rect 18367 25542 18377 25594
rect 18401 25542 18431 25594
rect 18431 25542 18443 25594
rect 18443 25542 18457 25594
rect 18481 25542 18495 25594
rect 18495 25542 18507 25594
rect 18507 25542 18537 25594
rect 18561 25542 18571 25594
rect 18571 25542 18617 25594
rect 18321 25540 18377 25542
rect 18401 25540 18457 25542
rect 18481 25540 18537 25542
rect 18561 25540 18617 25542
rect 14848 25050 14904 25052
rect 14928 25050 14984 25052
rect 15008 25050 15064 25052
rect 15088 25050 15144 25052
rect 14848 24998 14894 25050
rect 14894 24998 14904 25050
rect 14928 24998 14958 25050
rect 14958 24998 14970 25050
rect 14970 24998 14984 25050
rect 15008 24998 15022 25050
rect 15022 24998 15034 25050
rect 15034 24998 15064 25050
rect 15088 24998 15098 25050
rect 15098 24998 15144 25050
rect 14848 24996 14904 24998
rect 14928 24996 14984 24998
rect 15008 24996 15064 24998
rect 15088 24996 15144 24998
rect 21794 25050 21850 25052
rect 21874 25050 21930 25052
rect 21954 25050 22010 25052
rect 22034 25050 22090 25052
rect 21794 24998 21840 25050
rect 21840 24998 21850 25050
rect 21874 24998 21904 25050
rect 21904 24998 21916 25050
rect 21916 24998 21930 25050
rect 21954 24998 21968 25050
rect 21968 24998 21980 25050
rect 21980 24998 22010 25050
rect 22034 24998 22044 25050
rect 22044 24998 22090 25050
rect 21794 24996 21850 24998
rect 21874 24996 21930 24998
rect 21954 24996 22010 24998
rect 22034 24996 22090 24998
rect 18321 24506 18377 24508
rect 18401 24506 18457 24508
rect 18481 24506 18537 24508
rect 18561 24506 18617 24508
rect 18321 24454 18367 24506
rect 18367 24454 18377 24506
rect 18401 24454 18431 24506
rect 18431 24454 18443 24506
rect 18443 24454 18457 24506
rect 18481 24454 18495 24506
rect 18495 24454 18507 24506
rect 18507 24454 18537 24506
rect 18561 24454 18571 24506
rect 18571 24454 18617 24506
rect 18321 24452 18377 24454
rect 18401 24452 18457 24454
rect 18481 24452 18537 24454
rect 18561 24452 18617 24454
rect 14848 23962 14904 23964
rect 14928 23962 14984 23964
rect 15008 23962 15064 23964
rect 15088 23962 15144 23964
rect 14848 23910 14894 23962
rect 14894 23910 14904 23962
rect 14928 23910 14958 23962
rect 14958 23910 14970 23962
rect 14970 23910 14984 23962
rect 15008 23910 15022 23962
rect 15022 23910 15034 23962
rect 15034 23910 15064 23962
rect 15088 23910 15098 23962
rect 15098 23910 15144 23962
rect 14848 23908 14904 23910
rect 14928 23908 14984 23910
rect 15008 23908 15064 23910
rect 15088 23908 15144 23910
rect 21794 23962 21850 23964
rect 21874 23962 21930 23964
rect 21954 23962 22010 23964
rect 22034 23962 22090 23964
rect 21794 23910 21840 23962
rect 21840 23910 21850 23962
rect 21874 23910 21904 23962
rect 21904 23910 21916 23962
rect 21916 23910 21930 23962
rect 21954 23910 21968 23962
rect 21968 23910 21980 23962
rect 21980 23910 22010 23962
rect 22034 23910 22044 23962
rect 22044 23910 22090 23962
rect 21794 23908 21850 23910
rect 21874 23908 21930 23910
rect 21954 23908 22010 23910
rect 22034 23908 22090 23910
rect 18321 23418 18377 23420
rect 18401 23418 18457 23420
rect 18481 23418 18537 23420
rect 18561 23418 18617 23420
rect 18321 23366 18367 23418
rect 18367 23366 18377 23418
rect 18401 23366 18431 23418
rect 18431 23366 18443 23418
rect 18443 23366 18457 23418
rect 18481 23366 18495 23418
rect 18495 23366 18507 23418
rect 18507 23366 18537 23418
rect 18561 23366 18571 23418
rect 18571 23366 18617 23418
rect 18321 23364 18377 23366
rect 18401 23364 18457 23366
rect 18481 23364 18537 23366
rect 18561 23364 18617 23366
rect 14848 22874 14904 22876
rect 14928 22874 14984 22876
rect 15008 22874 15064 22876
rect 15088 22874 15144 22876
rect 14848 22822 14894 22874
rect 14894 22822 14904 22874
rect 14928 22822 14958 22874
rect 14958 22822 14970 22874
rect 14970 22822 14984 22874
rect 15008 22822 15022 22874
rect 15022 22822 15034 22874
rect 15034 22822 15064 22874
rect 15088 22822 15098 22874
rect 15098 22822 15144 22874
rect 14848 22820 14904 22822
rect 14928 22820 14984 22822
rect 15008 22820 15064 22822
rect 15088 22820 15144 22822
rect 14848 21786 14904 21788
rect 14928 21786 14984 21788
rect 15008 21786 15064 21788
rect 15088 21786 15144 21788
rect 14848 21734 14894 21786
rect 14894 21734 14904 21786
rect 14928 21734 14958 21786
rect 14958 21734 14970 21786
rect 14970 21734 14984 21786
rect 15008 21734 15022 21786
rect 15022 21734 15034 21786
rect 15034 21734 15064 21786
rect 15088 21734 15098 21786
rect 15098 21734 15144 21786
rect 14848 21732 14904 21734
rect 14928 21732 14984 21734
rect 15008 21732 15064 21734
rect 15088 21732 15144 21734
rect 14848 20698 14904 20700
rect 14928 20698 14984 20700
rect 15008 20698 15064 20700
rect 15088 20698 15144 20700
rect 14848 20646 14894 20698
rect 14894 20646 14904 20698
rect 14928 20646 14958 20698
rect 14958 20646 14970 20698
rect 14970 20646 14984 20698
rect 15008 20646 15022 20698
rect 15022 20646 15034 20698
rect 15034 20646 15064 20698
rect 15088 20646 15098 20698
rect 15098 20646 15144 20698
rect 14848 20644 14904 20646
rect 14928 20644 14984 20646
rect 15008 20644 15064 20646
rect 15088 20644 15144 20646
rect 14848 19610 14904 19612
rect 14928 19610 14984 19612
rect 15008 19610 15064 19612
rect 15088 19610 15144 19612
rect 14848 19558 14894 19610
rect 14894 19558 14904 19610
rect 14928 19558 14958 19610
rect 14958 19558 14970 19610
rect 14970 19558 14984 19610
rect 15008 19558 15022 19610
rect 15022 19558 15034 19610
rect 15034 19558 15064 19610
rect 15088 19558 15098 19610
rect 15098 19558 15144 19610
rect 14848 19556 14904 19558
rect 14928 19556 14984 19558
rect 15008 19556 15064 19558
rect 15088 19556 15144 19558
rect 14848 18522 14904 18524
rect 14928 18522 14984 18524
rect 15008 18522 15064 18524
rect 15088 18522 15144 18524
rect 14848 18470 14894 18522
rect 14894 18470 14904 18522
rect 14928 18470 14958 18522
rect 14958 18470 14970 18522
rect 14970 18470 14984 18522
rect 15008 18470 15022 18522
rect 15022 18470 15034 18522
rect 15034 18470 15064 18522
rect 15088 18470 15098 18522
rect 15098 18470 15144 18522
rect 14848 18468 14904 18470
rect 14928 18468 14984 18470
rect 15008 18468 15064 18470
rect 15088 18468 15144 18470
rect 14848 17434 14904 17436
rect 14928 17434 14984 17436
rect 15008 17434 15064 17436
rect 15088 17434 15144 17436
rect 14848 17382 14894 17434
rect 14894 17382 14904 17434
rect 14928 17382 14958 17434
rect 14958 17382 14970 17434
rect 14970 17382 14984 17434
rect 15008 17382 15022 17434
rect 15022 17382 15034 17434
rect 15034 17382 15064 17434
rect 15088 17382 15098 17434
rect 15098 17382 15144 17434
rect 14848 17380 14904 17382
rect 14928 17380 14984 17382
rect 15008 17380 15064 17382
rect 15088 17380 15144 17382
rect 13726 14320 13782 14376
rect 11375 12538 11431 12540
rect 11455 12538 11511 12540
rect 11535 12538 11591 12540
rect 11615 12538 11671 12540
rect 11375 12486 11421 12538
rect 11421 12486 11431 12538
rect 11455 12486 11485 12538
rect 11485 12486 11497 12538
rect 11497 12486 11511 12538
rect 11535 12486 11549 12538
rect 11549 12486 11561 12538
rect 11561 12486 11591 12538
rect 11615 12486 11625 12538
rect 11625 12486 11671 12538
rect 11375 12484 11431 12486
rect 11455 12484 11511 12486
rect 11535 12484 11591 12486
rect 11615 12484 11671 12486
rect 14848 16346 14904 16348
rect 14928 16346 14984 16348
rect 15008 16346 15064 16348
rect 15088 16346 15144 16348
rect 14848 16294 14894 16346
rect 14894 16294 14904 16346
rect 14928 16294 14958 16346
rect 14958 16294 14970 16346
rect 14970 16294 14984 16346
rect 15008 16294 15022 16346
rect 15022 16294 15034 16346
rect 15034 16294 15064 16346
rect 15088 16294 15098 16346
rect 15098 16294 15144 16346
rect 14848 16292 14904 16294
rect 14928 16292 14984 16294
rect 15008 16292 15064 16294
rect 15088 16292 15144 16294
rect 21794 22874 21850 22876
rect 21874 22874 21930 22876
rect 21954 22874 22010 22876
rect 22034 22874 22090 22876
rect 21794 22822 21840 22874
rect 21840 22822 21850 22874
rect 21874 22822 21904 22874
rect 21904 22822 21916 22874
rect 21916 22822 21930 22874
rect 21954 22822 21968 22874
rect 21968 22822 21980 22874
rect 21980 22822 22010 22874
rect 22034 22822 22044 22874
rect 22044 22822 22090 22874
rect 21794 22820 21850 22822
rect 21874 22820 21930 22822
rect 21954 22820 22010 22822
rect 22034 22820 22090 22822
rect 18321 22330 18377 22332
rect 18401 22330 18457 22332
rect 18481 22330 18537 22332
rect 18561 22330 18617 22332
rect 18321 22278 18367 22330
rect 18367 22278 18377 22330
rect 18401 22278 18431 22330
rect 18431 22278 18443 22330
rect 18443 22278 18457 22330
rect 18481 22278 18495 22330
rect 18495 22278 18507 22330
rect 18507 22278 18537 22330
rect 18561 22278 18571 22330
rect 18571 22278 18617 22330
rect 18321 22276 18377 22278
rect 18401 22276 18457 22278
rect 18481 22276 18537 22278
rect 18561 22276 18617 22278
rect 21794 21786 21850 21788
rect 21874 21786 21930 21788
rect 21954 21786 22010 21788
rect 22034 21786 22090 21788
rect 21794 21734 21840 21786
rect 21840 21734 21850 21786
rect 21874 21734 21904 21786
rect 21904 21734 21916 21786
rect 21916 21734 21930 21786
rect 21954 21734 21968 21786
rect 21968 21734 21980 21786
rect 21980 21734 22010 21786
rect 22034 21734 22044 21786
rect 22044 21734 22090 21786
rect 21794 21732 21850 21734
rect 21874 21732 21930 21734
rect 21954 21732 22010 21734
rect 22034 21732 22090 21734
rect 18321 21242 18377 21244
rect 18401 21242 18457 21244
rect 18481 21242 18537 21244
rect 18561 21242 18617 21244
rect 18321 21190 18367 21242
rect 18367 21190 18377 21242
rect 18401 21190 18431 21242
rect 18431 21190 18443 21242
rect 18443 21190 18457 21242
rect 18481 21190 18495 21242
rect 18495 21190 18507 21242
rect 18507 21190 18537 21242
rect 18561 21190 18571 21242
rect 18571 21190 18617 21242
rect 18321 21188 18377 21190
rect 18401 21188 18457 21190
rect 18481 21188 18537 21190
rect 18561 21188 18617 21190
rect 21794 20698 21850 20700
rect 21874 20698 21930 20700
rect 21954 20698 22010 20700
rect 22034 20698 22090 20700
rect 21794 20646 21840 20698
rect 21840 20646 21850 20698
rect 21874 20646 21904 20698
rect 21904 20646 21916 20698
rect 21916 20646 21930 20698
rect 21954 20646 21968 20698
rect 21968 20646 21980 20698
rect 21980 20646 22010 20698
rect 22034 20646 22044 20698
rect 22044 20646 22090 20698
rect 21794 20644 21850 20646
rect 21874 20644 21930 20646
rect 21954 20644 22010 20646
rect 22034 20644 22090 20646
rect 14848 15258 14904 15260
rect 14928 15258 14984 15260
rect 15008 15258 15064 15260
rect 15088 15258 15144 15260
rect 14848 15206 14894 15258
rect 14894 15206 14904 15258
rect 14928 15206 14958 15258
rect 14958 15206 14970 15258
rect 14970 15206 14984 15258
rect 15008 15206 15022 15258
rect 15022 15206 15034 15258
rect 15034 15206 15064 15258
rect 15088 15206 15098 15258
rect 15098 15206 15144 15258
rect 14848 15204 14904 15206
rect 14928 15204 14984 15206
rect 15008 15204 15064 15206
rect 15088 15204 15144 15206
rect 14848 14170 14904 14172
rect 14928 14170 14984 14172
rect 15008 14170 15064 14172
rect 15088 14170 15144 14172
rect 14848 14118 14894 14170
rect 14894 14118 14904 14170
rect 14928 14118 14958 14170
rect 14958 14118 14970 14170
rect 14970 14118 14984 14170
rect 15008 14118 15022 14170
rect 15022 14118 15034 14170
rect 15034 14118 15064 14170
rect 15088 14118 15098 14170
rect 15098 14118 15144 14170
rect 14848 14116 14904 14118
rect 14928 14116 14984 14118
rect 15008 14116 15064 14118
rect 15088 14116 15144 14118
rect 14848 13082 14904 13084
rect 14928 13082 14984 13084
rect 15008 13082 15064 13084
rect 15088 13082 15144 13084
rect 14848 13030 14894 13082
rect 14894 13030 14904 13082
rect 14928 13030 14958 13082
rect 14958 13030 14970 13082
rect 14970 13030 14984 13082
rect 15008 13030 15022 13082
rect 15022 13030 15034 13082
rect 15034 13030 15064 13082
rect 15088 13030 15098 13082
rect 15098 13030 15144 13082
rect 14848 13028 14904 13030
rect 14928 13028 14984 13030
rect 15008 13028 15064 13030
rect 15088 13028 15144 13030
rect 13726 12688 13782 12744
rect 11375 11450 11431 11452
rect 11455 11450 11511 11452
rect 11535 11450 11591 11452
rect 11615 11450 11671 11452
rect 11375 11398 11421 11450
rect 11421 11398 11431 11450
rect 11455 11398 11485 11450
rect 11485 11398 11497 11450
rect 11497 11398 11511 11450
rect 11535 11398 11549 11450
rect 11549 11398 11561 11450
rect 11561 11398 11591 11450
rect 11615 11398 11625 11450
rect 11625 11398 11671 11450
rect 11375 11396 11431 11398
rect 11455 11396 11511 11398
rect 11535 11396 11591 11398
rect 11615 11396 11671 11398
rect 11518 11192 11574 11248
rect 11375 10362 11431 10364
rect 11455 10362 11511 10364
rect 11535 10362 11591 10364
rect 11615 10362 11671 10364
rect 11375 10310 11421 10362
rect 11421 10310 11431 10362
rect 11455 10310 11485 10362
rect 11485 10310 11497 10362
rect 11497 10310 11511 10362
rect 11535 10310 11549 10362
rect 11549 10310 11561 10362
rect 11561 10310 11591 10362
rect 11615 10310 11625 10362
rect 11625 10310 11671 10362
rect 11375 10308 11431 10310
rect 11455 10308 11511 10310
rect 11535 10308 11591 10310
rect 11615 10308 11671 10310
rect 11978 11192 12034 11248
rect 11375 9274 11431 9276
rect 11455 9274 11511 9276
rect 11535 9274 11591 9276
rect 11615 9274 11671 9276
rect 11375 9222 11421 9274
rect 11421 9222 11431 9274
rect 11455 9222 11485 9274
rect 11485 9222 11497 9274
rect 11497 9222 11511 9274
rect 11535 9222 11549 9274
rect 11549 9222 11561 9274
rect 11561 9222 11591 9274
rect 11615 9222 11625 9274
rect 11625 9222 11671 9274
rect 11375 9220 11431 9222
rect 11455 9220 11511 9222
rect 11535 9220 11591 9222
rect 11615 9220 11671 9222
rect 11375 8186 11431 8188
rect 11455 8186 11511 8188
rect 11535 8186 11591 8188
rect 11615 8186 11671 8188
rect 11375 8134 11421 8186
rect 11421 8134 11431 8186
rect 11455 8134 11485 8186
rect 11485 8134 11497 8186
rect 11497 8134 11511 8186
rect 11535 8134 11549 8186
rect 11549 8134 11561 8186
rect 11561 8134 11591 8186
rect 11615 8134 11625 8186
rect 11625 8134 11671 8186
rect 11375 8132 11431 8134
rect 11455 8132 11511 8134
rect 11535 8132 11591 8134
rect 11615 8132 11671 8134
rect 15290 13368 15346 13424
rect 15750 13268 15752 13288
rect 15752 13268 15804 13288
rect 15804 13268 15806 13288
rect 15750 13232 15806 13268
rect 14848 11994 14904 11996
rect 14928 11994 14984 11996
rect 15008 11994 15064 11996
rect 15088 11994 15144 11996
rect 14848 11942 14894 11994
rect 14894 11942 14904 11994
rect 14928 11942 14958 11994
rect 14958 11942 14970 11994
rect 14970 11942 14984 11994
rect 15008 11942 15022 11994
rect 15022 11942 15034 11994
rect 15034 11942 15064 11994
rect 15088 11942 15098 11994
rect 15098 11942 15144 11994
rect 14848 11940 14904 11942
rect 14928 11940 14984 11942
rect 15008 11940 15064 11942
rect 15088 11940 15144 11942
rect 11375 7098 11431 7100
rect 11455 7098 11511 7100
rect 11535 7098 11591 7100
rect 11615 7098 11671 7100
rect 11375 7046 11421 7098
rect 11421 7046 11431 7098
rect 11455 7046 11485 7098
rect 11485 7046 11497 7098
rect 11497 7046 11511 7098
rect 11535 7046 11549 7098
rect 11549 7046 11561 7098
rect 11561 7046 11591 7098
rect 11615 7046 11625 7098
rect 11625 7046 11671 7098
rect 11375 7044 11431 7046
rect 11455 7044 11511 7046
rect 11535 7044 11591 7046
rect 11615 7044 11671 7046
rect 11375 6010 11431 6012
rect 11455 6010 11511 6012
rect 11535 6010 11591 6012
rect 11615 6010 11671 6012
rect 11375 5958 11421 6010
rect 11421 5958 11431 6010
rect 11455 5958 11485 6010
rect 11485 5958 11497 6010
rect 11497 5958 11511 6010
rect 11535 5958 11549 6010
rect 11549 5958 11561 6010
rect 11561 5958 11591 6010
rect 11615 5958 11625 6010
rect 11625 5958 11671 6010
rect 11375 5956 11431 5958
rect 11455 5956 11511 5958
rect 11535 5956 11591 5958
rect 11615 5956 11671 5958
rect 11375 4922 11431 4924
rect 11455 4922 11511 4924
rect 11535 4922 11591 4924
rect 11615 4922 11671 4924
rect 11375 4870 11421 4922
rect 11421 4870 11431 4922
rect 11455 4870 11485 4922
rect 11485 4870 11497 4922
rect 11497 4870 11511 4922
rect 11535 4870 11549 4922
rect 11549 4870 11561 4922
rect 11561 4870 11591 4922
rect 11615 4870 11625 4922
rect 11625 4870 11671 4922
rect 11375 4868 11431 4870
rect 11455 4868 11511 4870
rect 11535 4868 11591 4870
rect 11615 4868 11671 4870
rect 11334 4140 11390 4176
rect 11334 4120 11336 4140
rect 11336 4120 11388 4140
rect 11388 4120 11390 4140
rect 11375 3834 11431 3836
rect 11455 3834 11511 3836
rect 11535 3834 11591 3836
rect 11615 3834 11671 3836
rect 11375 3782 11421 3834
rect 11421 3782 11431 3834
rect 11455 3782 11485 3834
rect 11485 3782 11497 3834
rect 11497 3782 11511 3834
rect 11535 3782 11549 3834
rect 11549 3782 11561 3834
rect 11561 3782 11591 3834
rect 11615 3782 11625 3834
rect 11625 3782 11671 3834
rect 11375 3780 11431 3782
rect 11455 3780 11511 3782
rect 11535 3780 11591 3782
rect 11615 3780 11671 3782
rect 11375 2746 11431 2748
rect 11455 2746 11511 2748
rect 11535 2746 11591 2748
rect 11615 2746 11671 2748
rect 11375 2694 11421 2746
rect 11421 2694 11431 2746
rect 11455 2694 11485 2746
rect 11485 2694 11497 2746
rect 11497 2694 11511 2746
rect 11535 2694 11549 2746
rect 11549 2694 11561 2746
rect 11561 2694 11591 2746
rect 11615 2694 11625 2746
rect 11625 2694 11671 2746
rect 11375 2692 11431 2694
rect 11455 2692 11511 2694
rect 11535 2692 11591 2694
rect 11615 2692 11671 2694
rect 12254 3576 12310 3632
rect 13174 7384 13230 7440
rect 13266 7248 13322 7304
rect 14186 9580 14242 9616
rect 14186 9560 14188 9580
rect 14188 9560 14240 9580
rect 14240 9560 14242 9580
rect 14848 10906 14904 10908
rect 14928 10906 14984 10908
rect 15008 10906 15064 10908
rect 15088 10906 15144 10908
rect 14848 10854 14894 10906
rect 14894 10854 14904 10906
rect 14928 10854 14958 10906
rect 14958 10854 14970 10906
rect 14970 10854 14984 10906
rect 15008 10854 15022 10906
rect 15022 10854 15034 10906
rect 15034 10854 15064 10906
rect 15088 10854 15098 10906
rect 15098 10854 15144 10906
rect 14848 10852 14904 10854
rect 14928 10852 14984 10854
rect 15008 10852 15064 10854
rect 15088 10852 15144 10854
rect 14848 9818 14904 9820
rect 14928 9818 14984 9820
rect 15008 9818 15064 9820
rect 15088 9818 15144 9820
rect 14848 9766 14894 9818
rect 14894 9766 14904 9818
rect 14928 9766 14958 9818
rect 14958 9766 14970 9818
rect 14970 9766 14984 9818
rect 15008 9766 15022 9818
rect 15022 9766 15034 9818
rect 15034 9766 15064 9818
rect 15088 9766 15098 9818
rect 15098 9766 15144 9818
rect 14848 9764 14904 9766
rect 14928 9764 14984 9766
rect 15008 9764 15064 9766
rect 15088 9764 15144 9766
rect 14848 8730 14904 8732
rect 14928 8730 14984 8732
rect 15008 8730 15064 8732
rect 15088 8730 15144 8732
rect 14848 8678 14894 8730
rect 14894 8678 14904 8730
rect 14928 8678 14958 8730
rect 14958 8678 14970 8730
rect 14970 8678 14984 8730
rect 15008 8678 15022 8730
rect 15022 8678 15034 8730
rect 15034 8678 15064 8730
rect 15088 8678 15098 8730
rect 15098 8678 15144 8730
rect 14848 8676 14904 8678
rect 14928 8676 14984 8678
rect 15008 8676 15064 8678
rect 15088 8676 15144 8678
rect 15566 12280 15622 12336
rect 14848 7642 14904 7644
rect 14928 7642 14984 7644
rect 15008 7642 15064 7644
rect 15088 7642 15144 7644
rect 14848 7590 14894 7642
rect 14894 7590 14904 7642
rect 14928 7590 14958 7642
rect 14958 7590 14970 7642
rect 14970 7590 14984 7642
rect 15008 7590 15022 7642
rect 15022 7590 15034 7642
rect 15034 7590 15064 7642
rect 15088 7590 15098 7642
rect 15098 7590 15144 7642
rect 14848 7588 14904 7590
rect 14928 7588 14984 7590
rect 15008 7588 15064 7590
rect 15088 7588 15144 7590
rect 14848 6554 14904 6556
rect 14928 6554 14984 6556
rect 15008 6554 15064 6556
rect 15088 6554 15144 6556
rect 14848 6502 14894 6554
rect 14894 6502 14904 6554
rect 14928 6502 14958 6554
rect 14958 6502 14970 6554
rect 14970 6502 14984 6554
rect 15008 6502 15022 6554
rect 15022 6502 15034 6554
rect 15034 6502 15064 6554
rect 15088 6502 15098 6554
rect 15098 6502 15144 6554
rect 14848 6500 14904 6502
rect 14928 6500 14984 6502
rect 15008 6500 15064 6502
rect 15088 6500 15144 6502
rect 14848 5466 14904 5468
rect 14928 5466 14984 5468
rect 15008 5466 15064 5468
rect 15088 5466 15144 5468
rect 14848 5414 14894 5466
rect 14894 5414 14904 5466
rect 14928 5414 14958 5466
rect 14958 5414 14970 5466
rect 14970 5414 14984 5466
rect 15008 5414 15022 5466
rect 15022 5414 15034 5466
rect 15034 5414 15064 5466
rect 15088 5414 15098 5466
rect 15098 5414 15144 5466
rect 14848 5412 14904 5414
rect 14928 5412 14984 5414
rect 15008 5412 15064 5414
rect 15088 5412 15144 5414
rect 14848 4378 14904 4380
rect 14928 4378 14984 4380
rect 15008 4378 15064 4380
rect 15088 4378 15144 4380
rect 14848 4326 14894 4378
rect 14894 4326 14904 4378
rect 14928 4326 14958 4378
rect 14958 4326 14970 4378
rect 14970 4326 14984 4378
rect 15008 4326 15022 4378
rect 15022 4326 15034 4378
rect 15034 4326 15064 4378
rect 15088 4326 15098 4378
rect 15098 4326 15144 4378
rect 14848 4324 14904 4326
rect 14928 4324 14984 4326
rect 15008 4324 15064 4326
rect 15088 4324 15144 4326
rect 15198 3440 15254 3496
rect 14848 3290 14904 3292
rect 14928 3290 14984 3292
rect 15008 3290 15064 3292
rect 15088 3290 15144 3292
rect 14848 3238 14894 3290
rect 14894 3238 14904 3290
rect 14928 3238 14958 3290
rect 14958 3238 14970 3290
rect 14970 3238 14984 3290
rect 15008 3238 15022 3290
rect 15022 3238 15034 3290
rect 15034 3238 15064 3290
rect 15088 3238 15098 3290
rect 15098 3238 15144 3290
rect 14848 3236 14904 3238
rect 14928 3236 14984 3238
rect 15008 3236 15064 3238
rect 15088 3236 15144 3238
rect 18321 20154 18377 20156
rect 18401 20154 18457 20156
rect 18481 20154 18537 20156
rect 18561 20154 18617 20156
rect 18321 20102 18367 20154
rect 18367 20102 18377 20154
rect 18401 20102 18431 20154
rect 18431 20102 18443 20154
rect 18443 20102 18457 20154
rect 18481 20102 18495 20154
rect 18495 20102 18507 20154
rect 18507 20102 18537 20154
rect 18561 20102 18571 20154
rect 18571 20102 18617 20154
rect 18321 20100 18377 20102
rect 18401 20100 18457 20102
rect 18481 20100 18537 20102
rect 18561 20100 18617 20102
rect 21794 19610 21850 19612
rect 21874 19610 21930 19612
rect 21954 19610 22010 19612
rect 22034 19610 22090 19612
rect 21794 19558 21840 19610
rect 21840 19558 21850 19610
rect 21874 19558 21904 19610
rect 21904 19558 21916 19610
rect 21916 19558 21930 19610
rect 21954 19558 21968 19610
rect 21968 19558 21980 19610
rect 21980 19558 22010 19610
rect 22034 19558 22044 19610
rect 22044 19558 22090 19610
rect 21794 19556 21850 19558
rect 21874 19556 21930 19558
rect 21954 19556 22010 19558
rect 22034 19556 22090 19558
rect 18321 19066 18377 19068
rect 18401 19066 18457 19068
rect 18481 19066 18537 19068
rect 18561 19066 18617 19068
rect 18321 19014 18367 19066
rect 18367 19014 18377 19066
rect 18401 19014 18431 19066
rect 18431 19014 18443 19066
rect 18443 19014 18457 19066
rect 18481 19014 18495 19066
rect 18495 19014 18507 19066
rect 18507 19014 18537 19066
rect 18561 19014 18571 19066
rect 18571 19014 18617 19066
rect 18321 19012 18377 19014
rect 18401 19012 18457 19014
rect 18481 19012 18537 19014
rect 18561 19012 18617 19014
rect 16118 13776 16174 13832
rect 15934 11736 15990 11792
rect 15934 10512 15990 10568
rect 17130 12144 17186 12200
rect 21794 18522 21850 18524
rect 21874 18522 21930 18524
rect 21954 18522 22010 18524
rect 22034 18522 22090 18524
rect 21794 18470 21840 18522
rect 21840 18470 21850 18522
rect 21874 18470 21904 18522
rect 21904 18470 21916 18522
rect 21916 18470 21930 18522
rect 21954 18470 21968 18522
rect 21968 18470 21980 18522
rect 21980 18470 22010 18522
rect 22034 18470 22044 18522
rect 22044 18470 22090 18522
rect 21794 18468 21850 18470
rect 21874 18468 21930 18470
rect 21954 18468 22010 18470
rect 22034 18468 22090 18470
rect 18321 17978 18377 17980
rect 18401 17978 18457 17980
rect 18481 17978 18537 17980
rect 18561 17978 18617 17980
rect 18321 17926 18367 17978
rect 18367 17926 18377 17978
rect 18401 17926 18431 17978
rect 18431 17926 18443 17978
rect 18443 17926 18457 17978
rect 18481 17926 18495 17978
rect 18495 17926 18507 17978
rect 18507 17926 18537 17978
rect 18561 17926 18571 17978
rect 18571 17926 18617 17978
rect 18321 17924 18377 17926
rect 18401 17924 18457 17926
rect 18481 17924 18537 17926
rect 18561 17924 18617 17926
rect 21794 17434 21850 17436
rect 21874 17434 21930 17436
rect 21954 17434 22010 17436
rect 22034 17434 22090 17436
rect 21794 17382 21840 17434
rect 21840 17382 21850 17434
rect 21874 17382 21904 17434
rect 21904 17382 21916 17434
rect 21916 17382 21930 17434
rect 21954 17382 21968 17434
rect 21968 17382 21980 17434
rect 21980 17382 22010 17434
rect 22034 17382 22044 17434
rect 22044 17382 22090 17434
rect 21794 17380 21850 17382
rect 21874 17380 21930 17382
rect 21954 17380 22010 17382
rect 22034 17380 22090 17382
rect 18321 16890 18377 16892
rect 18401 16890 18457 16892
rect 18481 16890 18537 16892
rect 18561 16890 18617 16892
rect 18321 16838 18367 16890
rect 18367 16838 18377 16890
rect 18401 16838 18431 16890
rect 18431 16838 18443 16890
rect 18443 16838 18457 16890
rect 18481 16838 18495 16890
rect 18495 16838 18507 16890
rect 18507 16838 18537 16890
rect 18561 16838 18571 16890
rect 18571 16838 18617 16890
rect 18321 16836 18377 16838
rect 18401 16836 18457 16838
rect 18481 16836 18537 16838
rect 18561 16836 18617 16838
rect 21794 16346 21850 16348
rect 21874 16346 21930 16348
rect 21954 16346 22010 16348
rect 22034 16346 22090 16348
rect 21794 16294 21840 16346
rect 21840 16294 21850 16346
rect 21874 16294 21904 16346
rect 21904 16294 21916 16346
rect 21916 16294 21930 16346
rect 21954 16294 21968 16346
rect 21968 16294 21980 16346
rect 21980 16294 22010 16346
rect 22034 16294 22044 16346
rect 22044 16294 22090 16346
rect 21794 16292 21850 16294
rect 21874 16292 21930 16294
rect 21954 16292 22010 16294
rect 22034 16292 22090 16294
rect 18321 15802 18377 15804
rect 18401 15802 18457 15804
rect 18481 15802 18537 15804
rect 18561 15802 18617 15804
rect 18321 15750 18367 15802
rect 18367 15750 18377 15802
rect 18401 15750 18431 15802
rect 18431 15750 18443 15802
rect 18443 15750 18457 15802
rect 18481 15750 18495 15802
rect 18495 15750 18507 15802
rect 18507 15750 18537 15802
rect 18561 15750 18571 15802
rect 18571 15750 18617 15802
rect 18321 15748 18377 15750
rect 18401 15748 18457 15750
rect 18481 15748 18537 15750
rect 18561 15748 18617 15750
rect 21794 15258 21850 15260
rect 21874 15258 21930 15260
rect 21954 15258 22010 15260
rect 22034 15258 22090 15260
rect 21794 15206 21840 15258
rect 21840 15206 21850 15258
rect 21874 15206 21904 15258
rect 21904 15206 21916 15258
rect 21916 15206 21930 15258
rect 21954 15206 21968 15258
rect 21968 15206 21980 15258
rect 21980 15206 22010 15258
rect 22034 15206 22044 15258
rect 22044 15206 22090 15258
rect 21794 15204 21850 15206
rect 21874 15204 21930 15206
rect 21954 15204 22010 15206
rect 22034 15204 22090 15206
rect 18321 14714 18377 14716
rect 18401 14714 18457 14716
rect 18481 14714 18537 14716
rect 18561 14714 18617 14716
rect 18321 14662 18367 14714
rect 18367 14662 18377 14714
rect 18401 14662 18431 14714
rect 18431 14662 18443 14714
rect 18443 14662 18457 14714
rect 18481 14662 18495 14714
rect 18495 14662 18507 14714
rect 18507 14662 18537 14714
rect 18561 14662 18571 14714
rect 18571 14662 18617 14714
rect 18321 14660 18377 14662
rect 18401 14660 18457 14662
rect 18481 14660 18537 14662
rect 18561 14660 18617 14662
rect 28354 26696 28410 26752
rect 25267 26682 25323 26684
rect 25347 26682 25403 26684
rect 25427 26682 25483 26684
rect 25507 26682 25563 26684
rect 25267 26630 25313 26682
rect 25313 26630 25323 26682
rect 25347 26630 25377 26682
rect 25377 26630 25389 26682
rect 25389 26630 25403 26682
rect 25427 26630 25441 26682
rect 25441 26630 25453 26682
rect 25453 26630 25483 26682
rect 25507 26630 25517 26682
rect 25517 26630 25563 26682
rect 25267 26628 25323 26630
rect 25347 26628 25403 26630
rect 25427 26628 25483 26630
rect 25507 26628 25563 26630
rect 28740 26138 28796 26140
rect 28820 26138 28876 26140
rect 28900 26138 28956 26140
rect 28980 26138 29036 26140
rect 28740 26086 28786 26138
rect 28786 26086 28796 26138
rect 28820 26086 28850 26138
rect 28850 26086 28862 26138
rect 28862 26086 28876 26138
rect 28900 26086 28914 26138
rect 28914 26086 28926 26138
rect 28926 26086 28956 26138
rect 28980 26086 28990 26138
rect 28990 26086 29036 26138
rect 28740 26084 28796 26086
rect 28820 26084 28876 26086
rect 28900 26084 28956 26086
rect 28980 26084 29036 26086
rect 28354 25880 28410 25936
rect 25267 25594 25323 25596
rect 25347 25594 25403 25596
rect 25427 25594 25483 25596
rect 25507 25594 25563 25596
rect 25267 25542 25313 25594
rect 25313 25542 25323 25594
rect 25347 25542 25377 25594
rect 25377 25542 25389 25594
rect 25389 25542 25403 25594
rect 25427 25542 25441 25594
rect 25441 25542 25453 25594
rect 25453 25542 25483 25594
rect 25507 25542 25517 25594
rect 25517 25542 25563 25594
rect 25267 25540 25323 25542
rect 25347 25540 25403 25542
rect 25427 25540 25483 25542
rect 25507 25540 25563 25542
rect 25267 24506 25323 24508
rect 25347 24506 25403 24508
rect 25427 24506 25483 24508
rect 25507 24506 25563 24508
rect 25267 24454 25313 24506
rect 25313 24454 25323 24506
rect 25347 24454 25377 24506
rect 25377 24454 25389 24506
rect 25389 24454 25403 24506
rect 25427 24454 25441 24506
rect 25441 24454 25453 24506
rect 25453 24454 25483 24506
rect 25507 24454 25517 24506
rect 25517 24454 25563 24506
rect 25267 24452 25323 24454
rect 25347 24452 25403 24454
rect 25427 24452 25483 24454
rect 25507 24452 25563 24454
rect 25267 23418 25323 23420
rect 25347 23418 25403 23420
rect 25427 23418 25483 23420
rect 25507 23418 25563 23420
rect 25267 23366 25313 23418
rect 25313 23366 25323 23418
rect 25347 23366 25377 23418
rect 25377 23366 25389 23418
rect 25389 23366 25403 23418
rect 25427 23366 25441 23418
rect 25441 23366 25453 23418
rect 25453 23366 25483 23418
rect 25507 23366 25517 23418
rect 25517 23366 25563 23418
rect 25267 23364 25323 23366
rect 25347 23364 25403 23366
rect 25427 23364 25483 23366
rect 25507 23364 25563 23366
rect 25267 22330 25323 22332
rect 25347 22330 25403 22332
rect 25427 22330 25483 22332
rect 25507 22330 25563 22332
rect 25267 22278 25313 22330
rect 25313 22278 25323 22330
rect 25347 22278 25377 22330
rect 25377 22278 25389 22330
rect 25389 22278 25403 22330
rect 25427 22278 25441 22330
rect 25441 22278 25453 22330
rect 25453 22278 25483 22330
rect 25507 22278 25517 22330
rect 25517 22278 25563 22330
rect 25267 22276 25323 22278
rect 25347 22276 25403 22278
rect 25427 22276 25483 22278
rect 25507 22276 25563 22278
rect 25267 21242 25323 21244
rect 25347 21242 25403 21244
rect 25427 21242 25483 21244
rect 25507 21242 25563 21244
rect 25267 21190 25313 21242
rect 25313 21190 25323 21242
rect 25347 21190 25377 21242
rect 25377 21190 25389 21242
rect 25389 21190 25403 21242
rect 25427 21190 25441 21242
rect 25441 21190 25453 21242
rect 25453 21190 25483 21242
rect 25507 21190 25517 21242
rect 25517 21190 25563 21242
rect 25267 21188 25323 21190
rect 25347 21188 25403 21190
rect 25427 21188 25483 21190
rect 25507 21188 25563 21190
rect 25267 20154 25323 20156
rect 25347 20154 25403 20156
rect 25427 20154 25483 20156
rect 25507 20154 25563 20156
rect 25267 20102 25313 20154
rect 25313 20102 25323 20154
rect 25347 20102 25377 20154
rect 25377 20102 25389 20154
rect 25389 20102 25403 20154
rect 25427 20102 25441 20154
rect 25441 20102 25453 20154
rect 25453 20102 25483 20154
rect 25507 20102 25517 20154
rect 25517 20102 25563 20154
rect 25267 20100 25323 20102
rect 25347 20100 25403 20102
rect 25427 20100 25483 20102
rect 25507 20100 25563 20102
rect 25267 19066 25323 19068
rect 25347 19066 25403 19068
rect 25427 19066 25483 19068
rect 25507 19066 25563 19068
rect 25267 19014 25313 19066
rect 25313 19014 25323 19066
rect 25347 19014 25377 19066
rect 25377 19014 25389 19066
rect 25389 19014 25403 19066
rect 25427 19014 25441 19066
rect 25441 19014 25453 19066
rect 25453 19014 25483 19066
rect 25507 19014 25517 19066
rect 25517 19014 25563 19066
rect 25267 19012 25323 19014
rect 25347 19012 25403 19014
rect 25427 19012 25483 19014
rect 25507 19012 25563 19014
rect 25267 17978 25323 17980
rect 25347 17978 25403 17980
rect 25427 17978 25483 17980
rect 25507 17978 25563 17980
rect 25267 17926 25313 17978
rect 25313 17926 25323 17978
rect 25347 17926 25377 17978
rect 25377 17926 25389 17978
rect 25389 17926 25403 17978
rect 25427 17926 25441 17978
rect 25441 17926 25453 17978
rect 25453 17926 25483 17978
rect 25507 17926 25517 17978
rect 25517 17926 25563 17978
rect 25267 17924 25323 17926
rect 25347 17924 25403 17926
rect 25427 17924 25483 17926
rect 25507 17924 25563 17926
rect 25267 16890 25323 16892
rect 25347 16890 25403 16892
rect 25427 16890 25483 16892
rect 25507 16890 25563 16892
rect 25267 16838 25313 16890
rect 25313 16838 25323 16890
rect 25347 16838 25377 16890
rect 25377 16838 25389 16890
rect 25389 16838 25403 16890
rect 25427 16838 25441 16890
rect 25441 16838 25453 16890
rect 25453 16838 25483 16890
rect 25507 16838 25517 16890
rect 25517 16838 25563 16890
rect 25267 16836 25323 16838
rect 25347 16836 25403 16838
rect 25427 16836 25483 16838
rect 25507 16836 25563 16838
rect 21794 14170 21850 14172
rect 21874 14170 21930 14172
rect 21954 14170 22010 14172
rect 22034 14170 22090 14172
rect 21794 14118 21840 14170
rect 21840 14118 21850 14170
rect 21874 14118 21904 14170
rect 21904 14118 21916 14170
rect 21916 14118 21930 14170
rect 21954 14118 21968 14170
rect 21968 14118 21980 14170
rect 21980 14118 22010 14170
rect 22034 14118 22044 14170
rect 22044 14118 22090 14170
rect 21794 14116 21850 14118
rect 21874 14116 21930 14118
rect 21954 14116 22010 14118
rect 22034 14116 22090 14118
rect 18321 13626 18377 13628
rect 18401 13626 18457 13628
rect 18481 13626 18537 13628
rect 18561 13626 18617 13628
rect 18321 13574 18367 13626
rect 18367 13574 18377 13626
rect 18401 13574 18431 13626
rect 18431 13574 18443 13626
rect 18443 13574 18457 13626
rect 18481 13574 18495 13626
rect 18495 13574 18507 13626
rect 18507 13574 18537 13626
rect 18561 13574 18571 13626
rect 18571 13574 18617 13626
rect 18321 13572 18377 13574
rect 18401 13572 18457 13574
rect 18481 13572 18537 13574
rect 18561 13572 18617 13574
rect 21794 13082 21850 13084
rect 21874 13082 21930 13084
rect 21954 13082 22010 13084
rect 22034 13082 22090 13084
rect 21794 13030 21840 13082
rect 21840 13030 21850 13082
rect 21874 13030 21904 13082
rect 21904 13030 21916 13082
rect 21916 13030 21930 13082
rect 21954 13030 21968 13082
rect 21968 13030 21980 13082
rect 21980 13030 22010 13082
rect 22034 13030 22044 13082
rect 22044 13030 22090 13082
rect 21794 13028 21850 13030
rect 21874 13028 21930 13030
rect 21954 13028 22010 13030
rect 22034 13028 22090 13030
rect 18321 12538 18377 12540
rect 18401 12538 18457 12540
rect 18481 12538 18537 12540
rect 18561 12538 18617 12540
rect 18321 12486 18367 12538
rect 18367 12486 18377 12538
rect 18401 12486 18431 12538
rect 18431 12486 18443 12538
rect 18443 12486 18457 12538
rect 18481 12486 18495 12538
rect 18495 12486 18507 12538
rect 18507 12486 18537 12538
rect 18561 12486 18571 12538
rect 18571 12486 18617 12538
rect 18321 12484 18377 12486
rect 18401 12484 18457 12486
rect 18481 12484 18537 12486
rect 18561 12484 18617 12486
rect 18321 11450 18377 11452
rect 18401 11450 18457 11452
rect 18481 11450 18537 11452
rect 18561 11450 18617 11452
rect 18321 11398 18367 11450
rect 18367 11398 18377 11450
rect 18401 11398 18431 11450
rect 18431 11398 18443 11450
rect 18443 11398 18457 11450
rect 18481 11398 18495 11450
rect 18495 11398 18507 11450
rect 18507 11398 18537 11450
rect 18561 11398 18571 11450
rect 18571 11398 18617 11450
rect 18321 11396 18377 11398
rect 18401 11396 18457 11398
rect 18481 11396 18537 11398
rect 18561 11396 18617 11398
rect 18321 10362 18377 10364
rect 18401 10362 18457 10364
rect 18481 10362 18537 10364
rect 18561 10362 18617 10364
rect 18321 10310 18367 10362
rect 18367 10310 18377 10362
rect 18401 10310 18431 10362
rect 18431 10310 18443 10362
rect 18443 10310 18457 10362
rect 18481 10310 18495 10362
rect 18495 10310 18507 10362
rect 18507 10310 18537 10362
rect 18561 10310 18571 10362
rect 18571 10310 18617 10362
rect 18321 10308 18377 10310
rect 18401 10308 18457 10310
rect 18481 10308 18537 10310
rect 18561 10308 18617 10310
rect 18321 9274 18377 9276
rect 18401 9274 18457 9276
rect 18481 9274 18537 9276
rect 18561 9274 18617 9276
rect 18321 9222 18367 9274
rect 18367 9222 18377 9274
rect 18401 9222 18431 9274
rect 18431 9222 18443 9274
rect 18443 9222 18457 9274
rect 18481 9222 18495 9274
rect 18495 9222 18507 9274
rect 18507 9222 18537 9274
rect 18561 9222 18571 9274
rect 18571 9222 18617 9274
rect 18321 9220 18377 9222
rect 18401 9220 18457 9222
rect 18481 9220 18537 9222
rect 18561 9220 18617 9222
rect 18321 8186 18377 8188
rect 18401 8186 18457 8188
rect 18481 8186 18537 8188
rect 18561 8186 18617 8188
rect 18321 8134 18367 8186
rect 18367 8134 18377 8186
rect 18401 8134 18431 8186
rect 18431 8134 18443 8186
rect 18443 8134 18457 8186
rect 18481 8134 18495 8186
rect 18495 8134 18507 8186
rect 18507 8134 18537 8186
rect 18561 8134 18571 8186
rect 18571 8134 18617 8186
rect 18321 8132 18377 8134
rect 18401 8132 18457 8134
rect 18481 8132 18537 8134
rect 18561 8132 18617 8134
rect 18321 7098 18377 7100
rect 18401 7098 18457 7100
rect 18481 7098 18537 7100
rect 18561 7098 18617 7100
rect 18321 7046 18367 7098
rect 18367 7046 18377 7098
rect 18401 7046 18431 7098
rect 18431 7046 18443 7098
rect 18443 7046 18457 7098
rect 18481 7046 18495 7098
rect 18495 7046 18507 7098
rect 18507 7046 18537 7098
rect 18561 7046 18571 7098
rect 18571 7046 18617 7098
rect 18321 7044 18377 7046
rect 18401 7044 18457 7046
rect 18481 7044 18537 7046
rect 18561 7044 18617 7046
rect 18321 6010 18377 6012
rect 18401 6010 18457 6012
rect 18481 6010 18537 6012
rect 18561 6010 18617 6012
rect 18321 5958 18367 6010
rect 18367 5958 18377 6010
rect 18401 5958 18431 6010
rect 18431 5958 18443 6010
rect 18443 5958 18457 6010
rect 18481 5958 18495 6010
rect 18495 5958 18507 6010
rect 18507 5958 18537 6010
rect 18561 5958 18571 6010
rect 18571 5958 18617 6010
rect 18321 5956 18377 5958
rect 18401 5956 18457 5958
rect 18481 5956 18537 5958
rect 18561 5956 18617 5958
rect 18321 4922 18377 4924
rect 18401 4922 18457 4924
rect 18481 4922 18537 4924
rect 18561 4922 18617 4924
rect 18321 4870 18367 4922
rect 18367 4870 18377 4922
rect 18401 4870 18431 4922
rect 18431 4870 18443 4922
rect 18443 4870 18457 4922
rect 18481 4870 18495 4922
rect 18495 4870 18507 4922
rect 18507 4870 18537 4922
rect 18561 4870 18571 4922
rect 18571 4870 18617 4922
rect 18321 4868 18377 4870
rect 18401 4868 18457 4870
rect 18481 4868 18537 4870
rect 18561 4868 18617 4870
rect 18321 3834 18377 3836
rect 18401 3834 18457 3836
rect 18481 3834 18537 3836
rect 18561 3834 18617 3836
rect 18321 3782 18367 3834
rect 18367 3782 18377 3834
rect 18401 3782 18431 3834
rect 18431 3782 18443 3834
rect 18443 3782 18457 3834
rect 18481 3782 18495 3834
rect 18495 3782 18507 3834
rect 18507 3782 18537 3834
rect 18561 3782 18571 3834
rect 18571 3782 18617 3834
rect 18321 3780 18377 3782
rect 18401 3780 18457 3782
rect 18481 3780 18537 3782
rect 18561 3780 18617 3782
rect 21794 11994 21850 11996
rect 21874 11994 21930 11996
rect 21954 11994 22010 11996
rect 22034 11994 22090 11996
rect 21794 11942 21840 11994
rect 21840 11942 21850 11994
rect 21874 11942 21904 11994
rect 21904 11942 21916 11994
rect 21916 11942 21930 11994
rect 21954 11942 21968 11994
rect 21968 11942 21980 11994
rect 21980 11942 22010 11994
rect 22034 11942 22044 11994
rect 22044 11942 22090 11994
rect 21794 11940 21850 11942
rect 21874 11940 21930 11942
rect 21954 11940 22010 11942
rect 22034 11940 22090 11942
rect 21794 10906 21850 10908
rect 21874 10906 21930 10908
rect 21954 10906 22010 10908
rect 22034 10906 22090 10908
rect 21794 10854 21840 10906
rect 21840 10854 21850 10906
rect 21874 10854 21904 10906
rect 21904 10854 21916 10906
rect 21916 10854 21930 10906
rect 21954 10854 21968 10906
rect 21968 10854 21980 10906
rect 21980 10854 22010 10906
rect 22034 10854 22044 10906
rect 22044 10854 22090 10906
rect 21794 10852 21850 10854
rect 21874 10852 21930 10854
rect 21954 10852 22010 10854
rect 22034 10852 22090 10854
rect 21794 9818 21850 9820
rect 21874 9818 21930 9820
rect 21954 9818 22010 9820
rect 22034 9818 22090 9820
rect 21794 9766 21840 9818
rect 21840 9766 21850 9818
rect 21874 9766 21904 9818
rect 21904 9766 21916 9818
rect 21916 9766 21930 9818
rect 21954 9766 21968 9818
rect 21968 9766 21980 9818
rect 21980 9766 22010 9818
rect 22034 9766 22044 9818
rect 22044 9766 22090 9818
rect 21794 9764 21850 9766
rect 21874 9764 21930 9766
rect 21954 9764 22010 9766
rect 22034 9764 22090 9766
rect 21794 8730 21850 8732
rect 21874 8730 21930 8732
rect 21954 8730 22010 8732
rect 22034 8730 22090 8732
rect 21794 8678 21840 8730
rect 21840 8678 21850 8730
rect 21874 8678 21904 8730
rect 21904 8678 21916 8730
rect 21916 8678 21930 8730
rect 21954 8678 21968 8730
rect 21968 8678 21980 8730
rect 21980 8678 22010 8730
rect 22034 8678 22044 8730
rect 22044 8678 22090 8730
rect 21794 8676 21850 8678
rect 21874 8676 21930 8678
rect 21954 8676 22010 8678
rect 22034 8676 22090 8678
rect 21794 7642 21850 7644
rect 21874 7642 21930 7644
rect 21954 7642 22010 7644
rect 22034 7642 22090 7644
rect 21794 7590 21840 7642
rect 21840 7590 21850 7642
rect 21874 7590 21904 7642
rect 21904 7590 21916 7642
rect 21916 7590 21930 7642
rect 21954 7590 21968 7642
rect 21968 7590 21980 7642
rect 21980 7590 22010 7642
rect 22034 7590 22044 7642
rect 22044 7590 22090 7642
rect 21794 7588 21850 7590
rect 21874 7588 21930 7590
rect 21954 7588 22010 7590
rect 22034 7588 22090 7590
rect 21794 6554 21850 6556
rect 21874 6554 21930 6556
rect 21954 6554 22010 6556
rect 22034 6554 22090 6556
rect 21794 6502 21840 6554
rect 21840 6502 21850 6554
rect 21874 6502 21904 6554
rect 21904 6502 21916 6554
rect 21916 6502 21930 6554
rect 21954 6502 21968 6554
rect 21968 6502 21980 6554
rect 21980 6502 22010 6554
rect 22034 6502 22044 6554
rect 22044 6502 22090 6554
rect 21794 6500 21850 6502
rect 21874 6500 21930 6502
rect 21954 6500 22010 6502
rect 22034 6500 22090 6502
rect 21794 5466 21850 5468
rect 21874 5466 21930 5468
rect 21954 5466 22010 5468
rect 22034 5466 22090 5468
rect 21794 5414 21840 5466
rect 21840 5414 21850 5466
rect 21874 5414 21904 5466
rect 21904 5414 21916 5466
rect 21916 5414 21930 5466
rect 21954 5414 21968 5466
rect 21968 5414 21980 5466
rect 21980 5414 22010 5466
rect 22034 5414 22044 5466
rect 22044 5414 22090 5466
rect 21794 5412 21850 5414
rect 21874 5412 21930 5414
rect 21954 5412 22010 5414
rect 22034 5412 22090 5414
rect 20902 4684 20958 4720
rect 20902 4664 20904 4684
rect 20904 4664 20956 4684
rect 20956 4664 20958 4684
rect 21794 4378 21850 4380
rect 21874 4378 21930 4380
rect 21954 4378 22010 4380
rect 22034 4378 22090 4380
rect 21794 4326 21840 4378
rect 21840 4326 21850 4378
rect 21874 4326 21904 4378
rect 21904 4326 21916 4378
rect 21916 4326 21930 4378
rect 21954 4326 21968 4378
rect 21968 4326 21980 4378
rect 21980 4326 22010 4378
rect 22034 4326 22044 4378
rect 22044 4326 22090 4378
rect 21794 4324 21850 4326
rect 21874 4324 21930 4326
rect 21954 4324 22010 4326
rect 22034 4324 22090 4326
rect 25267 15802 25323 15804
rect 25347 15802 25403 15804
rect 25427 15802 25483 15804
rect 25507 15802 25563 15804
rect 25267 15750 25313 15802
rect 25313 15750 25323 15802
rect 25347 15750 25377 15802
rect 25377 15750 25389 15802
rect 25389 15750 25403 15802
rect 25427 15750 25441 15802
rect 25441 15750 25453 15802
rect 25453 15750 25483 15802
rect 25507 15750 25517 15802
rect 25517 15750 25563 15802
rect 25267 15748 25323 15750
rect 25347 15748 25403 15750
rect 25427 15748 25483 15750
rect 25507 15748 25563 15750
rect 25267 14714 25323 14716
rect 25347 14714 25403 14716
rect 25427 14714 25483 14716
rect 25507 14714 25563 14716
rect 25267 14662 25313 14714
rect 25313 14662 25323 14714
rect 25347 14662 25377 14714
rect 25377 14662 25389 14714
rect 25389 14662 25403 14714
rect 25427 14662 25441 14714
rect 25441 14662 25453 14714
rect 25453 14662 25483 14714
rect 25507 14662 25517 14714
rect 25517 14662 25563 14714
rect 25267 14660 25323 14662
rect 25347 14660 25403 14662
rect 25427 14660 25483 14662
rect 25507 14660 25563 14662
rect 25267 13626 25323 13628
rect 25347 13626 25403 13628
rect 25427 13626 25483 13628
rect 25507 13626 25563 13628
rect 25267 13574 25313 13626
rect 25313 13574 25323 13626
rect 25347 13574 25377 13626
rect 25377 13574 25389 13626
rect 25389 13574 25403 13626
rect 25427 13574 25441 13626
rect 25441 13574 25453 13626
rect 25453 13574 25483 13626
rect 25507 13574 25517 13626
rect 25517 13574 25563 13626
rect 25267 13572 25323 13574
rect 25347 13572 25403 13574
rect 25427 13572 25483 13574
rect 25507 13572 25563 13574
rect 28354 25064 28410 25120
rect 28740 25050 28796 25052
rect 28820 25050 28876 25052
rect 28900 25050 28956 25052
rect 28980 25050 29036 25052
rect 28740 24998 28786 25050
rect 28786 24998 28796 25050
rect 28820 24998 28850 25050
rect 28850 24998 28862 25050
rect 28862 24998 28876 25050
rect 28900 24998 28914 25050
rect 28914 24998 28926 25050
rect 28926 24998 28956 25050
rect 28980 24998 28990 25050
rect 28990 24998 29036 25050
rect 28740 24996 28796 24998
rect 28820 24996 28876 24998
rect 28900 24996 28956 24998
rect 28980 24996 29036 24998
rect 28354 24248 28410 24304
rect 28740 23962 28796 23964
rect 28820 23962 28876 23964
rect 28900 23962 28956 23964
rect 28980 23962 29036 23964
rect 28740 23910 28786 23962
rect 28786 23910 28796 23962
rect 28820 23910 28850 23962
rect 28850 23910 28862 23962
rect 28862 23910 28876 23962
rect 28900 23910 28914 23962
rect 28914 23910 28926 23962
rect 28926 23910 28956 23962
rect 28980 23910 28990 23962
rect 28990 23910 29036 23962
rect 28740 23908 28796 23910
rect 28820 23908 28876 23910
rect 28900 23908 28956 23910
rect 28980 23908 29036 23910
rect 28722 23432 28778 23488
rect 28740 22874 28796 22876
rect 28820 22874 28876 22876
rect 28900 22874 28956 22876
rect 28980 22874 29036 22876
rect 28740 22822 28786 22874
rect 28786 22822 28796 22874
rect 28820 22822 28850 22874
rect 28850 22822 28862 22874
rect 28862 22822 28876 22874
rect 28900 22822 28914 22874
rect 28914 22822 28926 22874
rect 28926 22822 28956 22874
rect 28980 22822 28990 22874
rect 28990 22822 29036 22874
rect 28740 22820 28796 22822
rect 28820 22820 28876 22822
rect 28900 22820 28956 22822
rect 28980 22820 29036 22822
rect 28354 22616 28410 22672
rect 28814 22092 28870 22128
rect 28814 22072 28816 22092
rect 28816 22072 28868 22092
rect 28868 22072 28870 22092
rect 28740 21786 28796 21788
rect 28820 21786 28876 21788
rect 28900 21786 28956 21788
rect 28980 21786 29036 21788
rect 28740 21734 28786 21786
rect 28786 21734 28796 21786
rect 28820 21734 28850 21786
rect 28850 21734 28862 21786
rect 28862 21734 28876 21786
rect 28900 21734 28914 21786
rect 28914 21734 28926 21786
rect 28926 21734 28956 21786
rect 28980 21734 28990 21786
rect 28990 21734 29036 21786
rect 28740 21732 28796 21734
rect 28820 21732 28876 21734
rect 28900 21732 28956 21734
rect 28980 21732 29036 21734
rect 28354 20984 28410 21040
rect 28740 20698 28796 20700
rect 28820 20698 28876 20700
rect 28900 20698 28956 20700
rect 28980 20698 29036 20700
rect 28740 20646 28786 20698
rect 28786 20646 28796 20698
rect 28820 20646 28850 20698
rect 28850 20646 28862 20698
rect 28862 20646 28876 20698
rect 28900 20646 28914 20698
rect 28914 20646 28926 20698
rect 28926 20646 28956 20698
rect 28980 20646 28990 20698
rect 28990 20646 29036 20698
rect 28740 20644 28796 20646
rect 28820 20644 28876 20646
rect 28900 20644 28956 20646
rect 28980 20644 29036 20646
rect 28354 20168 28410 20224
rect 28740 19610 28796 19612
rect 28820 19610 28876 19612
rect 28900 19610 28956 19612
rect 28980 19610 29036 19612
rect 28740 19558 28786 19610
rect 28786 19558 28796 19610
rect 28820 19558 28850 19610
rect 28850 19558 28862 19610
rect 28862 19558 28876 19610
rect 28900 19558 28914 19610
rect 28914 19558 28926 19610
rect 28926 19558 28956 19610
rect 28980 19558 28990 19610
rect 28990 19558 29036 19610
rect 28740 19556 28796 19558
rect 28820 19556 28876 19558
rect 28900 19556 28956 19558
rect 28980 19556 29036 19558
rect 28354 19352 28410 19408
rect 28814 18828 28870 18864
rect 28814 18808 28816 18828
rect 28816 18808 28868 18828
rect 28868 18808 28870 18828
rect 28740 18522 28796 18524
rect 28820 18522 28876 18524
rect 28900 18522 28956 18524
rect 28980 18522 29036 18524
rect 28740 18470 28786 18522
rect 28786 18470 28796 18522
rect 28820 18470 28850 18522
rect 28850 18470 28862 18522
rect 28862 18470 28876 18522
rect 28900 18470 28914 18522
rect 28914 18470 28926 18522
rect 28926 18470 28956 18522
rect 28980 18470 28990 18522
rect 28990 18470 29036 18522
rect 28740 18468 28796 18470
rect 28820 18468 28876 18470
rect 28900 18468 28956 18470
rect 28980 18468 29036 18470
rect 28354 17720 28410 17776
rect 28740 17434 28796 17436
rect 28820 17434 28876 17436
rect 28900 17434 28956 17436
rect 28980 17434 29036 17436
rect 28740 17382 28786 17434
rect 28786 17382 28796 17434
rect 28820 17382 28850 17434
rect 28850 17382 28862 17434
rect 28862 17382 28876 17434
rect 28900 17382 28914 17434
rect 28914 17382 28926 17434
rect 28926 17382 28956 17434
rect 28980 17382 28990 17434
rect 28990 17382 29036 17434
rect 28740 17380 28796 17382
rect 28820 17380 28876 17382
rect 28900 17380 28956 17382
rect 28980 17380 29036 17382
rect 28354 16904 28410 16960
rect 28740 16346 28796 16348
rect 28820 16346 28876 16348
rect 28900 16346 28956 16348
rect 28980 16346 29036 16348
rect 28740 16294 28786 16346
rect 28786 16294 28796 16346
rect 28820 16294 28850 16346
rect 28850 16294 28862 16346
rect 28862 16294 28876 16346
rect 28900 16294 28914 16346
rect 28914 16294 28926 16346
rect 28926 16294 28956 16346
rect 28980 16294 28990 16346
rect 28990 16294 29036 16346
rect 28740 16292 28796 16294
rect 28820 16292 28876 16294
rect 28900 16292 28956 16294
rect 28980 16292 29036 16294
rect 28354 16088 28410 16144
rect 28354 15272 28410 15328
rect 28740 15258 28796 15260
rect 28820 15258 28876 15260
rect 28900 15258 28956 15260
rect 28980 15258 29036 15260
rect 28740 15206 28786 15258
rect 28786 15206 28796 15258
rect 28820 15206 28850 15258
rect 28850 15206 28862 15258
rect 28862 15206 28876 15258
rect 28900 15206 28914 15258
rect 28914 15206 28926 15258
rect 28926 15206 28956 15258
rect 28980 15206 28990 15258
rect 28990 15206 29036 15258
rect 28740 15204 28796 15206
rect 28820 15204 28876 15206
rect 28900 15204 28956 15206
rect 28980 15204 29036 15206
rect 26974 14456 27030 14512
rect 28354 14456 28410 14512
rect 28740 14170 28796 14172
rect 28820 14170 28876 14172
rect 28900 14170 28956 14172
rect 28980 14170 29036 14172
rect 28740 14118 28786 14170
rect 28786 14118 28796 14170
rect 28820 14118 28850 14170
rect 28850 14118 28862 14170
rect 28862 14118 28876 14170
rect 28900 14118 28914 14170
rect 28914 14118 28926 14170
rect 28926 14118 28956 14170
rect 28980 14118 28990 14170
rect 28990 14118 29036 14170
rect 28740 14116 28796 14118
rect 28820 14116 28876 14118
rect 28900 14116 28956 14118
rect 28980 14116 29036 14118
rect 28354 13640 28410 13696
rect 28740 13082 28796 13084
rect 28820 13082 28876 13084
rect 28900 13082 28956 13084
rect 28980 13082 29036 13084
rect 28740 13030 28786 13082
rect 28786 13030 28796 13082
rect 28820 13030 28850 13082
rect 28850 13030 28862 13082
rect 28862 13030 28876 13082
rect 28900 13030 28914 13082
rect 28914 13030 28926 13082
rect 28926 13030 28956 13082
rect 28980 13030 28990 13082
rect 28990 13030 29036 13082
rect 28740 13028 28796 13030
rect 28820 13028 28876 13030
rect 28900 13028 28956 13030
rect 28980 13028 29036 13030
rect 28354 12824 28410 12880
rect 25267 12538 25323 12540
rect 25347 12538 25403 12540
rect 25427 12538 25483 12540
rect 25507 12538 25563 12540
rect 25267 12486 25313 12538
rect 25313 12486 25323 12538
rect 25347 12486 25377 12538
rect 25377 12486 25389 12538
rect 25389 12486 25403 12538
rect 25427 12486 25441 12538
rect 25441 12486 25453 12538
rect 25453 12486 25483 12538
rect 25507 12486 25517 12538
rect 25517 12486 25563 12538
rect 25267 12484 25323 12486
rect 25347 12484 25403 12486
rect 25427 12484 25483 12486
rect 25507 12484 25563 12486
rect 28354 12008 28410 12064
rect 28740 11994 28796 11996
rect 28820 11994 28876 11996
rect 28900 11994 28956 11996
rect 28980 11994 29036 11996
rect 28740 11942 28786 11994
rect 28786 11942 28796 11994
rect 28820 11942 28850 11994
rect 28850 11942 28862 11994
rect 28862 11942 28876 11994
rect 28900 11942 28914 11994
rect 28914 11942 28926 11994
rect 28926 11942 28956 11994
rect 28980 11942 28990 11994
rect 28990 11942 29036 11994
rect 28740 11940 28796 11942
rect 28820 11940 28876 11942
rect 28900 11940 28956 11942
rect 28980 11940 29036 11942
rect 25267 11450 25323 11452
rect 25347 11450 25403 11452
rect 25427 11450 25483 11452
rect 25507 11450 25563 11452
rect 25267 11398 25313 11450
rect 25313 11398 25323 11450
rect 25347 11398 25377 11450
rect 25377 11398 25389 11450
rect 25389 11398 25403 11450
rect 25427 11398 25441 11450
rect 25441 11398 25453 11450
rect 25453 11398 25483 11450
rect 25507 11398 25517 11450
rect 25517 11398 25563 11450
rect 25267 11396 25323 11398
rect 25347 11396 25403 11398
rect 25427 11396 25483 11398
rect 25507 11396 25563 11398
rect 28354 11192 28410 11248
rect 28740 10906 28796 10908
rect 28820 10906 28876 10908
rect 28900 10906 28956 10908
rect 28980 10906 29036 10908
rect 28740 10854 28786 10906
rect 28786 10854 28796 10906
rect 28820 10854 28850 10906
rect 28850 10854 28862 10906
rect 28862 10854 28876 10906
rect 28900 10854 28914 10906
rect 28914 10854 28926 10906
rect 28926 10854 28956 10906
rect 28980 10854 28990 10906
rect 28990 10854 29036 10906
rect 28740 10852 28796 10854
rect 28820 10852 28876 10854
rect 28900 10852 28956 10854
rect 28980 10852 29036 10854
rect 28354 10376 28410 10432
rect 25267 10362 25323 10364
rect 25347 10362 25403 10364
rect 25427 10362 25483 10364
rect 25507 10362 25563 10364
rect 25267 10310 25313 10362
rect 25313 10310 25323 10362
rect 25347 10310 25377 10362
rect 25377 10310 25389 10362
rect 25389 10310 25403 10362
rect 25427 10310 25441 10362
rect 25441 10310 25453 10362
rect 25453 10310 25483 10362
rect 25507 10310 25517 10362
rect 25517 10310 25563 10362
rect 25267 10308 25323 10310
rect 25347 10308 25403 10310
rect 25427 10308 25483 10310
rect 25507 10308 25563 10310
rect 28740 9818 28796 9820
rect 28820 9818 28876 9820
rect 28900 9818 28956 9820
rect 28980 9818 29036 9820
rect 28740 9766 28786 9818
rect 28786 9766 28796 9818
rect 28820 9766 28850 9818
rect 28850 9766 28862 9818
rect 28862 9766 28876 9818
rect 28900 9766 28914 9818
rect 28914 9766 28926 9818
rect 28926 9766 28956 9818
rect 28980 9766 28990 9818
rect 28990 9766 29036 9818
rect 28740 9764 28796 9766
rect 28820 9764 28876 9766
rect 28900 9764 28956 9766
rect 28980 9764 29036 9766
rect 28354 9560 28410 9616
rect 18321 2746 18377 2748
rect 18401 2746 18457 2748
rect 18481 2746 18537 2748
rect 18561 2746 18617 2748
rect 18321 2694 18367 2746
rect 18367 2694 18377 2746
rect 18401 2694 18431 2746
rect 18431 2694 18443 2746
rect 18443 2694 18457 2746
rect 18481 2694 18495 2746
rect 18495 2694 18507 2746
rect 18507 2694 18537 2746
rect 18561 2694 18571 2746
rect 18571 2694 18617 2746
rect 18321 2692 18377 2694
rect 18401 2692 18457 2694
rect 18481 2692 18537 2694
rect 18561 2692 18617 2694
rect 14848 2202 14904 2204
rect 14928 2202 14984 2204
rect 15008 2202 15064 2204
rect 15088 2202 15144 2204
rect 14848 2150 14894 2202
rect 14894 2150 14904 2202
rect 14928 2150 14958 2202
rect 14958 2150 14970 2202
rect 14970 2150 14984 2202
rect 15008 2150 15022 2202
rect 15022 2150 15034 2202
rect 15034 2150 15064 2202
rect 15088 2150 15098 2202
rect 15098 2150 15144 2202
rect 14848 2148 14904 2150
rect 14928 2148 14984 2150
rect 15008 2148 15064 2150
rect 15088 2148 15144 2150
rect 21794 3290 21850 3292
rect 21874 3290 21930 3292
rect 21954 3290 22010 3292
rect 22034 3290 22090 3292
rect 21794 3238 21840 3290
rect 21840 3238 21850 3290
rect 21874 3238 21904 3290
rect 21904 3238 21916 3290
rect 21916 3238 21930 3290
rect 21954 3238 21968 3290
rect 21968 3238 21980 3290
rect 21980 3238 22010 3290
rect 22034 3238 22044 3290
rect 22044 3238 22090 3290
rect 21794 3236 21850 3238
rect 21874 3236 21930 3238
rect 21954 3236 22010 3238
rect 22034 3236 22090 3238
rect 21822 2896 21878 2952
rect 21794 2202 21850 2204
rect 21874 2202 21930 2204
rect 21954 2202 22010 2204
rect 22034 2202 22090 2204
rect 21794 2150 21840 2202
rect 21840 2150 21850 2202
rect 21874 2150 21904 2202
rect 21904 2150 21916 2202
rect 21916 2150 21930 2202
rect 21954 2150 21968 2202
rect 21968 2150 21980 2202
rect 21980 2150 22010 2202
rect 22034 2150 22044 2202
rect 22044 2150 22090 2202
rect 21794 2148 21850 2150
rect 21874 2148 21930 2150
rect 21954 2148 22010 2150
rect 22034 2148 22090 2150
rect 23386 2896 23442 2952
rect 25267 9274 25323 9276
rect 25347 9274 25403 9276
rect 25427 9274 25483 9276
rect 25507 9274 25563 9276
rect 25267 9222 25313 9274
rect 25313 9222 25323 9274
rect 25347 9222 25377 9274
rect 25377 9222 25389 9274
rect 25389 9222 25403 9274
rect 25427 9222 25441 9274
rect 25441 9222 25453 9274
rect 25453 9222 25483 9274
rect 25507 9222 25517 9274
rect 25517 9222 25563 9274
rect 25267 9220 25323 9222
rect 25347 9220 25403 9222
rect 25427 9220 25483 9222
rect 25507 9220 25563 9222
rect 25267 8186 25323 8188
rect 25347 8186 25403 8188
rect 25427 8186 25483 8188
rect 25507 8186 25563 8188
rect 25267 8134 25313 8186
rect 25313 8134 25323 8186
rect 25347 8134 25377 8186
rect 25377 8134 25389 8186
rect 25389 8134 25403 8186
rect 25427 8134 25441 8186
rect 25441 8134 25453 8186
rect 25453 8134 25483 8186
rect 25507 8134 25517 8186
rect 25517 8134 25563 8186
rect 25267 8132 25323 8134
rect 25347 8132 25403 8134
rect 25427 8132 25483 8134
rect 25507 8132 25563 8134
rect 24122 6160 24178 6216
rect 25267 7098 25323 7100
rect 25347 7098 25403 7100
rect 25427 7098 25483 7100
rect 25507 7098 25563 7100
rect 25267 7046 25313 7098
rect 25313 7046 25323 7098
rect 25347 7046 25377 7098
rect 25377 7046 25389 7098
rect 25389 7046 25403 7098
rect 25427 7046 25441 7098
rect 25441 7046 25453 7098
rect 25453 7046 25483 7098
rect 25507 7046 25517 7098
rect 25517 7046 25563 7098
rect 25267 7044 25323 7046
rect 25347 7044 25403 7046
rect 25427 7044 25483 7046
rect 25507 7044 25563 7046
rect 24674 3032 24730 3088
rect 25267 6010 25323 6012
rect 25347 6010 25403 6012
rect 25427 6010 25483 6012
rect 25507 6010 25563 6012
rect 25267 5958 25313 6010
rect 25313 5958 25323 6010
rect 25347 5958 25377 6010
rect 25377 5958 25389 6010
rect 25389 5958 25403 6010
rect 25427 5958 25441 6010
rect 25441 5958 25453 6010
rect 25453 5958 25483 6010
rect 25507 5958 25517 6010
rect 25517 5958 25563 6010
rect 25267 5956 25323 5958
rect 25347 5956 25403 5958
rect 25427 5956 25483 5958
rect 25507 5956 25563 5958
rect 25267 4922 25323 4924
rect 25347 4922 25403 4924
rect 25427 4922 25483 4924
rect 25507 4922 25563 4924
rect 25267 4870 25313 4922
rect 25313 4870 25323 4922
rect 25347 4870 25377 4922
rect 25377 4870 25389 4922
rect 25389 4870 25403 4922
rect 25427 4870 25441 4922
rect 25441 4870 25453 4922
rect 25453 4870 25483 4922
rect 25507 4870 25517 4922
rect 25517 4870 25563 4922
rect 25267 4868 25323 4870
rect 25347 4868 25403 4870
rect 25427 4868 25483 4870
rect 25507 4868 25563 4870
rect 28814 9036 28870 9072
rect 28814 9016 28816 9036
rect 28816 9016 28868 9036
rect 28868 9016 28870 9036
rect 25870 4664 25926 4720
rect 25267 3834 25323 3836
rect 25347 3834 25403 3836
rect 25427 3834 25483 3836
rect 25507 3834 25563 3836
rect 25267 3782 25313 3834
rect 25313 3782 25323 3834
rect 25347 3782 25377 3834
rect 25377 3782 25389 3834
rect 25389 3782 25403 3834
rect 25427 3782 25441 3834
rect 25441 3782 25453 3834
rect 25453 3782 25483 3834
rect 25507 3782 25517 3834
rect 25517 3782 25563 3834
rect 25267 3780 25323 3782
rect 25347 3780 25403 3782
rect 25427 3780 25483 3782
rect 25507 3780 25563 3782
rect 25267 2746 25323 2748
rect 25347 2746 25403 2748
rect 25427 2746 25483 2748
rect 25507 2746 25563 2748
rect 25267 2694 25313 2746
rect 25313 2694 25323 2746
rect 25347 2694 25377 2746
rect 25377 2694 25389 2746
rect 25389 2694 25403 2746
rect 25427 2694 25441 2746
rect 25441 2694 25453 2746
rect 25453 2694 25483 2746
rect 25507 2694 25517 2746
rect 25517 2694 25563 2746
rect 25267 2692 25323 2694
rect 25347 2692 25403 2694
rect 25427 2692 25483 2694
rect 25507 2692 25563 2694
rect 25594 2352 25650 2408
rect 28740 8730 28796 8732
rect 28820 8730 28876 8732
rect 28900 8730 28956 8732
rect 28980 8730 29036 8732
rect 28740 8678 28786 8730
rect 28786 8678 28796 8730
rect 28820 8678 28850 8730
rect 28850 8678 28862 8730
rect 28862 8678 28876 8730
rect 28900 8678 28914 8730
rect 28914 8678 28926 8730
rect 28926 8678 28956 8730
rect 28980 8678 28990 8730
rect 28990 8678 29036 8730
rect 28740 8676 28796 8678
rect 28820 8676 28876 8678
rect 28900 8676 28956 8678
rect 28980 8676 29036 8678
rect 26882 3848 26938 3904
rect 28354 7928 28410 7984
rect 28740 7642 28796 7644
rect 28820 7642 28876 7644
rect 28900 7642 28956 7644
rect 28980 7642 29036 7644
rect 28740 7590 28786 7642
rect 28786 7590 28796 7642
rect 28820 7590 28850 7642
rect 28850 7590 28862 7642
rect 28862 7590 28876 7642
rect 28900 7590 28914 7642
rect 28914 7590 28926 7642
rect 28926 7590 28956 7642
rect 28980 7590 28990 7642
rect 28990 7590 29036 7642
rect 28740 7588 28796 7590
rect 28820 7588 28876 7590
rect 28900 7588 28956 7590
rect 28980 7588 29036 7590
rect 28354 7112 28410 7168
rect 28740 6554 28796 6556
rect 28820 6554 28876 6556
rect 28900 6554 28956 6556
rect 28980 6554 29036 6556
rect 28740 6502 28786 6554
rect 28786 6502 28796 6554
rect 28820 6502 28850 6554
rect 28850 6502 28862 6554
rect 28862 6502 28876 6554
rect 28900 6502 28914 6554
rect 28914 6502 28926 6554
rect 28926 6502 28956 6554
rect 28980 6502 28990 6554
rect 28990 6502 29036 6554
rect 28740 6500 28796 6502
rect 28820 6500 28876 6502
rect 28900 6500 28956 6502
rect 28980 6500 29036 6502
rect 28354 6296 28410 6352
rect 28814 5772 28870 5808
rect 28814 5752 28816 5772
rect 28816 5752 28868 5772
rect 28868 5752 28870 5772
rect 28740 5466 28796 5468
rect 28820 5466 28876 5468
rect 28900 5466 28956 5468
rect 28980 5466 29036 5468
rect 28740 5414 28786 5466
rect 28786 5414 28796 5466
rect 28820 5414 28850 5466
rect 28850 5414 28862 5466
rect 28862 5414 28876 5466
rect 28900 5414 28914 5466
rect 28914 5414 28926 5466
rect 28926 5414 28956 5466
rect 28980 5414 28990 5466
rect 28990 5414 29036 5466
rect 28740 5412 28796 5414
rect 28820 5412 28876 5414
rect 28900 5412 28956 5414
rect 28980 5412 29036 5414
rect 28722 4664 28778 4720
rect 28740 4378 28796 4380
rect 28820 4378 28876 4380
rect 28900 4378 28956 4380
rect 28980 4378 29036 4380
rect 28740 4326 28786 4378
rect 28786 4326 28796 4378
rect 28820 4326 28850 4378
rect 28850 4326 28862 4378
rect 28862 4326 28876 4378
rect 28900 4326 28914 4378
rect 28914 4326 28926 4378
rect 28926 4326 28956 4378
rect 28980 4326 28990 4378
rect 28990 4326 29036 4378
rect 28740 4324 28796 4326
rect 28820 4324 28876 4326
rect 28900 4324 28956 4326
rect 28980 4324 29036 4326
rect 28740 3290 28796 3292
rect 28820 3290 28876 3292
rect 28900 3290 28956 3292
rect 28980 3290 29036 3292
rect 28740 3238 28786 3290
rect 28786 3238 28796 3290
rect 28820 3238 28850 3290
rect 28850 3238 28862 3290
rect 28862 3238 28876 3290
rect 28900 3238 28914 3290
rect 28914 3238 28926 3290
rect 28926 3238 28956 3290
rect 28980 3238 28990 3290
rect 28990 3238 29036 3290
rect 28740 3236 28796 3238
rect 28820 3236 28876 3238
rect 28900 3236 28956 3238
rect 28980 3236 29036 3238
rect 28630 2896 28686 2952
rect 28740 2202 28796 2204
rect 28820 2202 28876 2204
rect 28900 2202 28956 2204
rect 28980 2202 29036 2204
rect 28740 2150 28786 2202
rect 28786 2150 28796 2202
rect 28820 2150 28850 2202
rect 28850 2150 28862 2202
rect 28862 2150 28876 2202
rect 28900 2150 28914 2202
rect 28914 2150 28926 2202
rect 28926 2150 28956 2202
rect 28980 2150 28990 2202
rect 28990 2150 29036 2202
rect 28740 2148 28796 2150
rect 28820 2148 28876 2150
rect 28900 2148 28956 2150
rect 28980 2148 29036 2150
<< metal3 >>
rect 4419 27776 4735 27777
rect 4419 27712 4425 27776
rect 4489 27712 4505 27776
rect 4569 27712 4585 27776
rect 4649 27712 4665 27776
rect 4729 27712 4735 27776
rect 4419 27711 4735 27712
rect 11365 27776 11681 27777
rect 11365 27712 11371 27776
rect 11435 27712 11451 27776
rect 11515 27712 11531 27776
rect 11595 27712 11611 27776
rect 11675 27712 11681 27776
rect 11365 27711 11681 27712
rect 18311 27776 18627 27777
rect 18311 27712 18317 27776
rect 18381 27712 18397 27776
rect 18461 27712 18477 27776
rect 18541 27712 18557 27776
rect 18621 27712 18627 27776
rect 18311 27711 18627 27712
rect 25257 27776 25573 27777
rect 25257 27712 25263 27776
rect 25327 27712 25343 27776
rect 25407 27712 25423 27776
rect 25487 27712 25503 27776
rect 25567 27712 25573 27776
rect 25257 27711 25573 27712
rect 28533 27570 28599 27573
rect 29200 27570 30000 27600
rect 28533 27568 30000 27570
rect 28533 27512 28538 27568
rect 28594 27512 30000 27568
rect 28533 27510 30000 27512
rect 28533 27507 28599 27510
rect 29200 27480 30000 27510
rect 7892 27232 8208 27233
rect 7892 27168 7898 27232
rect 7962 27168 7978 27232
rect 8042 27168 8058 27232
rect 8122 27168 8138 27232
rect 8202 27168 8208 27232
rect 7892 27167 8208 27168
rect 14838 27232 15154 27233
rect 14838 27168 14844 27232
rect 14908 27168 14924 27232
rect 14988 27168 15004 27232
rect 15068 27168 15084 27232
rect 15148 27168 15154 27232
rect 14838 27167 15154 27168
rect 21784 27232 22100 27233
rect 21784 27168 21790 27232
rect 21854 27168 21870 27232
rect 21934 27168 21950 27232
rect 22014 27168 22030 27232
rect 22094 27168 22100 27232
rect 21784 27167 22100 27168
rect 28730 27232 29046 27233
rect 28730 27168 28736 27232
rect 28800 27168 28816 27232
rect 28880 27168 28896 27232
rect 28960 27168 28976 27232
rect 29040 27168 29046 27232
rect 28730 27167 29046 27168
rect 28349 26754 28415 26757
rect 29200 26754 30000 26784
rect 28349 26752 30000 26754
rect 28349 26696 28354 26752
rect 28410 26696 30000 26752
rect 28349 26694 30000 26696
rect 28349 26691 28415 26694
rect 4419 26688 4735 26689
rect 4419 26624 4425 26688
rect 4489 26624 4505 26688
rect 4569 26624 4585 26688
rect 4649 26624 4665 26688
rect 4729 26624 4735 26688
rect 4419 26623 4735 26624
rect 11365 26688 11681 26689
rect 11365 26624 11371 26688
rect 11435 26624 11451 26688
rect 11515 26624 11531 26688
rect 11595 26624 11611 26688
rect 11675 26624 11681 26688
rect 11365 26623 11681 26624
rect 18311 26688 18627 26689
rect 18311 26624 18317 26688
rect 18381 26624 18397 26688
rect 18461 26624 18477 26688
rect 18541 26624 18557 26688
rect 18621 26624 18627 26688
rect 18311 26623 18627 26624
rect 25257 26688 25573 26689
rect 25257 26624 25263 26688
rect 25327 26624 25343 26688
rect 25407 26624 25423 26688
rect 25487 26624 25503 26688
rect 25567 26624 25573 26688
rect 29200 26664 30000 26694
rect 25257 26623 25573 26624
rect 7892 26144 8208 26145
rect 7892 26080 7898 26144
rect 7962 26080 7978 26144
rect 8042 26080 8058 26144
rect 8122 26080 8138 26144
rect 8202 26080 8208 26144
rect 7892 26079 8208 26080
rect 14838 26144 15154 26145
rect 14838 26080 14844 26144
rect 14908 26080 14924 26144
rect 14988 26080 15004 26144
rect 15068 26080 15084 26144
rect 15148 26080 15154 26144
rect 14838 26079 15154 26080
rect 21784 26144 22100 26145
rect 21784 26080 21790 26144
rect 21854 26080 21870 26144
rect 21934 26080 21950 26144
rect 22014 26080 22030 26144
rect 22094 26080 22100 26144
rect 21784 26079 22100 26080
rect 28730 26144 29046 26145
rect 28730 26080 28736 26144
rect 28800 26080 28816 26144
rect 28880 26080 28896 26144
rect 28960 26080 28976 26144
rect 29040 26080 29046 26144
rect 28730 26079 29046 26080
rect 28349 25938 28415 25941
rect 29200 25938 30000 25968
rect 28349 25936 30000 25938
rect 28349 25880 28354 25936
rect 28410 25880 30000 25936
rect 28349 25878 30000 25880
rect 28349 25875 28415 25878
rect 29200 25848 30000 25878
rect 4419 25600 4735 25601
rect 4419 25536 4425 25600
rect 4489 25536 4505 25600
rect 4569 25536 4585 25600
rect 4649 25536 4665 25600
rect 4729 25536 4735 25600
rect 4419 25535 4735 25536
rect 11365 25600 11681 25601
rect 11365 25536 11371 25600
rect 11435 25536 11451 25600
rect 11515 25536 11531 25600
rect 11595 25536 11611 25600
rect 11675 25536 11681 25600
rect 11365 25535 11681 25536
rect 18311 25600 18627 25601
rect 18311 25536 18317 25600
rect 18381 25536 18397 25600
rect 18461 25536 18477 25600
rect 18541 25536 18557 25600
rect 18621 25536 18627 25600
rect 18311 25535 18627 25536
rect 25257 25600 25573 25601
rect 25257 25536 25263 25600
rect 25327 25536 25343 25600
rect 25407 25536 25423 25600
rect 25487 25536 25503 25600
rect 25567 25536 25573 25600
rect 25257 25535 25573 25536
rect 28352 25198 29194 25258
rect 28352 25125 28412 25198
rect 29134 25156 29194 25198
rect 29134 25152 29378 25156
rect 28349 25120 28415 25125
rect 28349 25064 28354 25120
rect 28410 25064 28415 25120
rect 29134 25096 30000 25152
rect 28349 25059 28415 25064
rect 7892 25056 8208 25057
rect 7892 24992 7898 25056
rect 7962 24992 7978 25056
rect 8042 24992 8058 25056
rect 8122 24992 8138 25056
rect 8202 24992 8208 25056
rect 7892 24991 8208 24992
rect 14838 25056 15154 25057
rect 14838 24992 14844 25056
rect 14908 24992 14924 25056
rect 14988 24992 15004 25056
rect 15068 24992 15084 25056
rect 15148 24992 15154 25056
rect 14838 24991 15154 24992
rect 21784 25056 22100 25057
rect 21784 24992 21790 25056
rect 21854 24992 21870 25056
rect 21934 24992 21950 25056
rect 22014 24992 22030 25056
rect 22094 24992 22100 25056
rect 21784 24991 22100 24992
rect 28730 25056 29046 25057
rect 28730 24992 28736 25056
rect 28800 24992 28816 25056
rect 28880 24992 28896 25056
rect 28960 24992 28976 25056
rect 29040 24992 29046 25056
rect 29200 25032 30000 25096
rect 28730 24991 29046 24992
rect 4419 24512 4735 24513
rect 4419 24448 4425 24512
rect 4489 24448 4505 24512
rect 4569 24448 4585 24512
rect 4649 24448 4665 24512
rect 4729 24448 4735 24512
rect 4419 24447 4735 24448
rect 11365 24512 11681 24513
rect 11365 24448 11371 24512
rect 11435 24448 11451 24512
rect 11515 24448 11531 24512
rect 11595 24448 11611 24512
rect 11675 24448 11681 24512
rect 11365 24447 11681 24448
rect 18311 24512 18627 24513
rect 18311 24448 18317 24512
rect 18381 24448 18397 24512
rect 18461 24448 18477 24512
rect 18541 24448 18557 24512
rect 18621 24448 18627 24512
rect 18311 24447 18627 24448
rect 25257 24512 25573 24513
rect 25257 24448 25263 24512
rect 25327 24448 25343 24512
rect 25407 24448 25423 24512
rect 25487 24448 25503 24512
rect 25567 24448 25573 24512
rect 25257 24447 25573 24448
rect 28349 24306 28415 24309
rect 29200 24306 30000 24336
rect 28349 24304 30000 24306
rect 28349 24248 28354 24304
rect 28410 24248 30000 24304
rect 28349 24246 30000 24248
rect 28349 24243 28415 24246
rect 29200 24216 30000 24246
rect 7892 23968 8208 23969
rect 7892 23904 7898 23968
rect 7962 23904 7978 23968
rect 8042 23904 8058 23968
rect 8122 23904 8138 23968
rect 8202 23904 8208 23968
rect 7892 23903 8208 23904
rect 14838 23968 15154 23969
rect 14838 23904 14844 23968
rect 14908 23904 14924 23968
rect 14988 23904 15004 23968
rect 15068 23904 15084 23968
rect 15148 23904 15154 23968
rect 14838 23903 15154 23904
rect 21784 23968 22100 23969
rect 21784 23904 21790 23968
rect 21854 23904 21870 23968
rect 21934 23904 21950 23968
rect 22014 23904 22030 23968
rect 22094 23904 22100 23968
rect 21784 23903 22100 23904
rect 28730 23968 29046 23969
rect 28730 23904 28736 23968
rect 28800 23904 28816 23968
rect 28880 23904 28896 23968
rect 28960 23904 28976 23968
rect 29040 23904 29046 23968
rect 28730 23903 29046 23904
rect 0 23400 800 23520
rect 1393 23490 1459 23493
rect 936 23488 1459 23490
rect 936 23432 1398 23488
rect 1454 23432 1459 23488
rect 936 23430 1459 23432
rect 0 23218 800 23248
rect 936 23218 996 23430
rect 1393 23427 1459 23430
rect 28717 23490 28783 23493
rect 29200 23490 30000 23520
rect 28717 23488 30000 23490
rect 28717 23432 28722 23488
rect 28778 23432 30000 23488
rect 28717 23430 30000 23432
rect 28717 23427 28783 23430
rect 4419 23424 4735 23425
rect 4419 23360 4425 23424
rect 4489 23360 4505 23424
rect 4569 23360 4585 23424
rect 4649 23360 4665 23424
rect 4729 23360 4735 23424
rect 4419 23359 4735 23360
rect 11365 23424 11681 23425
rect 11365 23360 11371 23424
rect 11435 23360 11451 23424
rect 11515 23360 11531 23424
rect 11595 23360 11611 23424
rect 11675 23360 11681 23424
rect 11365 23359 11681 23360
rect 18311 23424 18627 23425
rect 18311 23360 18317 23424
rect 18381 23360 18397 23424
rect 18461 23360 18477 23424
rect 18541 23360 18557 23424
rect 18621 23360 18627 23424
rect 18311 23359 18627 23360
rect 25257 23424 25573 23425
rect 25257 23360 25263 23424
rect 25327 23360 25343 23424
rect 25407 23360 25423 23424
rect 25487 23360 25503 23424
rect 25567 23360 25573 23424
rect 29200 23400 30000 23430
rect 25257 23359 25573 23360
rect 0 23158 996 23218
rect 0 23128 800 23158
rect 0 22946 800 22976
rect 1025 22946 1091 22949
rect 0 22944 1091 22946
rect 0 22888 1030 22944
rect 1086 22888 1091 22944
rect 0 22886 1091 22888
rect 0 22856 800 22886
rect 1025 22883 1091 22886
rect 7892 22880 8208 22881
rect 7892 22816 7898 22880
rect 7962 22816 7978 22880
rect 8042 22816 8058 22880
rect 8122 22816 8138 22880
rect 8202 22816 8208 22880
rect 7892 22815 8208 22816
rect 14838 22880 15154 22881
rect 14838 22816 14844 22880
rect 14908 22816 14924 22880
rect 14988 22816 15004 22880
rect 15068 22816 15084 22880
rect 15148 22816 15154 22880
rect 14838 22815 15154 22816
rect 21784 22880 22100 22881
rect 21784 22816 21790 22880
rect 21854 22816 21870 22880
rect 21934 22816 21950 22880
rect 22014 22816 22030 22880
rect 22094 22816 22100 22880
rect 21784 22815 22100 22816
rect 28730 22880 29046 22881
rect 28730 22816 28736 22880
rect 28800 22816 28816 22880
rect 28880 22816 28896 22880
rect 28960 22816 28976 22880
rect 29040 22816 29046 22880
rect 28730 22815 29046 22816
rect 0 22674 800 22704
rect 933 22674 999 22677
rect 0 22672 999 22674
rect 0 22616 938 22672
rect 994 22616 999 22672
rect 0 22614 999 22616
rect 0 22584 800 22614
rect 933 22611 999 22614
rect 28349 22674 28415 22677
rect 29200 22674 30000 22704
rect 28349 22672 30000 22674
rect 28349 22616 28354 22672
rect 28410 22616 30000 22672
rect 28349 22614 30000 22616
rect 28349 22611 28415 22614
rect 29200 22584 30000 22614
rect 0 22402 800 22432
rect 933 22402 999 22405
rect 0 22400 999 22402
rect 0 22344 938 22400
rect 994 22344 999 22400
rect 0 22342 999 22344
rect 0 22312 800 22342
rect 933 22339 999 22342
rect 4419 22336 4735 22337
rect 4419 22272 4425 22336
rect 4489 22272 4505 22336
rect 4569 22272 4585 22336
rect 4649 22272 4665 22336
rect 4729 22272 4735 22336
rect 4419 22271 4735 22272
rect 11365 22336 11681 22337
rect 11365 22272 11371 22336
rect 11435 22272 11451 22336
rect 11515 22272 11531 22336
rect 11595 22272 11611 22336
rect 11675 22272 11681 22336
rect 11365 22271 11681 22272
rect 18311 22336 18627 22337
rect 18311 22272 18317 22336
rect 18381 22272 18397 22336
rect 18461 22272 18477 22336
rect 18541 22272 18557 22336
rect 18621 22272 18627 22336
rect 18311 22271 18627 22272
rect 25257 22336 25573 22337
rect 25257 22272 25263 22336
rect 25327 22272 25343 22336
rect 25407 22272 25423 22336
rect 25487 22272 25503 22336
rect 25567 22272 25573 22336
rect 25257 22271 25573 22272
rect 0 22130 800 22160
rect 1025 22130 1091 22133
rect 0 22128 1091 22130
rect 0 22072 1030 22128
rect 1086 22072 1091 22128
rect 0 22070 1091 22072
rect 0 22040 800 22070
rect 1025 22067 1091 22070
rect 28809 22130 28875 22133
rect 28809 22128 29378 22130
rect 28809 22072 28814 22128
rect 28870 22072 29378 22128
rect 28809 22070 29378 22072
rect 28809 22067 28875 22070
rect 29318 21888 29378 22070
rect 0 21858 800 21888
rect 1025 21858 1091 21861
rect 0 21856 1091 21858
rect 0 21800 1030 21856
rect 1086 21800 1091 21856
rect 0 21798 1091 21800
rect 0 21768 800 21798
rect 1025 21795 1091 21798
rect 7892 21792 8208 21793
rect 7892 21728 7898 21792
rect 7962 21728 7978 21792
rect 8042 21728 8058 21792
rect 8122 21728 8138 21792
rect 8202 21728 8208 21792
rect 7892 21727 8208 21728
rect 14838 21792 15154 21793
rect 14838 21728 14844 21792
rect 14908 21728 14924 21792
rect 14988 21728 15004 21792
rect 15068 21728 15084 21792
rect 15148 21728 15154 21792
rect 14838 21727 15154 21728
rect 21784 21792 22100 21793
rect 21784 21728 21790 21792
rect 21854 21728 21870 21792
rect 21934 21728 21950 21792
rect 22014 21728 22030 21792
rect 22094 21728 22100 21792
rect 21784 21727 22100 21728
rect 28730 21792 29046 21793
rect 28730 21728 28736 21792
rect 28800 21728 28816 21792
rect 28880 21728 28896 21792
rect 28960 21728 28976 21792
rect 29040 21728 29046 21792
rect 29200 21768 30000 21888
rect 28730 21727 29046 21728
rect 0 21586 800 21616
rect 933 21586 999 21589
rect 0 21584 999 21586
rect 0 21528 938 21584
rect 994 21528 999 21584
rect 0 21526 999 21528
rect 0 21496 800 21526
rect 933 21523 999 21526
rect 0 21314 800 21344
rect 933 21314 999 21317
rect 0 21312 999 21314
rect 0 21256 938 21312
rect 994 21256 999 21312
rect 0 21254 999 21256
rect 0 21224 800 21254
rect 933 21251 999 21254
rect 4419 21248 4735 21249
rect 4419 21184 4425 21248
rect 4489 21184 4505 21248
rect 4569 21184 4585 21248
rect 4649 21184 4665 21248
rect 4729 21184 4735 21248
rect 4419 21183 4735 21184
rect 11365 21248 11681 21249
rect 11365 21184 11371 21248
rect 11435 21184 11451 21248
rect 11515 21184 11531 21248
rect 11595 21184 11611 21248
rect 11675 21184 11681 21248
rect 11365 21183 11681 21184
rect 18311 21248 18627 21249
rect 18311 21184 18317 21248
rect 18381 21184 18397 21248
rect 18461 21184 18477 21248
rect 18541 21184 18557 21248
rect 18621 21184 18627 21248
rect 18311 21183 18627 21184
rect 25257 21248 25573 21249
rect 25257 21184 25263 21248
rect 25327 21184 25343 21248
rect 25407 21184 25423 21248
rect 25487 21184 25503 21248
rect 25567 21184 25573 21248
rect 25257 21183 25573 21184
rect 0 21042 800 21072
rect 1025 21042 1091 21045
rect 0 21040 1091 21042
rect 0 20984 1030 21040
rect 1086 20984 1091 21040
rect 0 20982 1091 20984
rect 0 20952 800 20982
rect 1025 20979 1091 20982
rect 28349 21042 28415 21045
rect 29200 21042 30000 21072
rect 28349 21040 30000 21042
rect 28349 20984 28354 21040
rect 28410 20984 30000 21040
rect 28349 20982 30000 20984
rect 28349 20979 28415 20982
rect 29200 20952 30000 20982
rect 0 20770 800 20800
rect 933 20770 999 20773
rect 0 20768 999 20770
rect 0 20712 938 20768
rect 994 20712 999 20768
rect 0 20710 999 20712
rect 0 20680 800 20710
rect 933 20707 999 20710
rect 7892 20704 8208 20705
rect 7892 20640 7898 20704
rect 7962 20640 7978 20704
rect 8042 20640 8058 20704
rect 8122 20640 8138 20704
rect 8202 20640 8208 20704
rect 7892 20639 8208 20640
rect 14838 20704 15154 20705
rect 14838 20640 14844 20704
rect 14908 20640 14924 20704
rect 14988 20640 15004 20704
rect 15068 20640 15084 20704
rect 15148 20640 15154 20704
rect 14838 20639 15154 20640
rect 21784 20704 22100 20705
rect 21784 20640 21790 20704
rect 21854 20640 21870 20704
rect 21934 20640 21950 20704
rect 22014 20640 22030 20704
rect 22094 20640 22100 20704
rect 21784 20639 22100 20640
rect 28730 20704 29046 20705
rect 28730 20640 28736 20704
rect 28800 20640 28816 20704
rect 28880 20640 28896 20704
rect 28960 20640 28976 20704
rect 29040 20640 29046 20704
rect 28730 20639 29046 20640
rect 1393 20634 1459 20637
rect 936 20632 1459 20634
rect 936 20576 1398 20632
rect 1454 20576 1459 20632
rect 936 20574 1459 20576
rect 0 20498 800 20528
rect 936 20498 996 20574
rect 1393 20571 1459 20574
rect 0 20438 996 20498
rect 0 20408 800 20438
rect 0 20226 800 20256
rect 1025 20226 1091 20229
rect 0 20224 1091 20226
rect 0 20168 1030 20224
rect 1086 20168 1091 20224
rect 0 20166 1091 20168
rect 0 20136 800 20166
rect 1025 20163 1091 20166
rect 28349 20226 28415 20229
rect 29200 20226 30000 20256
rect 28349 20224 30000 20226
rect 28349 20168 28354 20224
rect 28410 20168 30000 20224
rect 28349 20166 30000 20168
rect 28349 20163 28415 20166
rect 4419 20160 4735 20161
rect 4419 20096 4425 20160
rect 4489 20096 4505 20160
rect 4569 20096 4585 20160
rect 4649 20096 4665 20160
rect 4729 20096 4735 20160
rect 4419 20095 4735 20096
rect 11365 20160 11681 20161
rect 11365 20096 11371 20160
rect 11435 20096 11451 20160
rect 11515 20096 11531 20160
rect 11595 20096 11611 20160
rect 11675 20096 11681 20160
rect 11365 20095 11681 20096
rect 18311 20160 18627 20161
rect 18311 20096 18317 20160
rect 18381 20096 18397 20160
rect 18461 20096 18477 20160
rect 18541 20096 18557 20160
rect 18621 20096 18627 20160
rect 18311 20095 18627 20096
rect 25257 20160 25573 20161
rect 25257 20096 25263 20160
rect 25327 20096 25343 20160
rect 25407 20096 25423 20160
rect 25487 20096 25503 20160
rect 25567 20096 25573 20160
rect 29200 20136 30000 20166
rect 25257 20095 25573 20096
rect 0 19954 800 19984
rect 933 19954 999 19957
rect 0 19952 999 19954
rect 0 19896 938 19952
rect 994 19896 999 19952
rect 0 19894 999 19896
rect 0 19864 800 19894
rect 933 19891 999 19894
rect 0 19682 800 19712
rect 1025 19682 1091 19685
rect 0 19680 1091 19682
rect 0 19624 1030 19680
rect 1086 19624 1091 19680
rect 0 19622 1091 19624
rect 0 19592 800 19622
rect 1025 19619 1091 19622
rect 7892 19616 8208 19617
rect 7892 19552 7898 19616
rect 7962 19552 7978 19616
rect 8042 19552 8058 19616
rect 8122 19552 8138 19616
rect 8202 19552 8208 19616
rect 7892 19551 8208 19552
rect 14838 19616 15154 19617
rect 14838 19552 14844 19616
rect 14908 19552 14924 19616
rect 14988 19552 15004 19616
rect 15068 19552 15084 19616
rect 15148 19552 15154 19616
rect 14838 19551 15154 19552
rect 21784 19616 22100 19617
rect 21784 19552 21790 19616
rect 21854 19552 21870 19616
rect 21934 19552 21950 19616
rect 22014 19552 22030 19616
rect 22094 19552 22100 19616
rect 21784 19551 22100 19552
rect 28730 19616 29046 19617
rect 28730 19552 28736 19616
rect 28800 19552 28816 19616
rect 28880 19552 28896 19616
rect 28960 19552 28976 19616
rect 29040 19552 29046 19616
rect 28730 19551 29046 19552
rect 0 19410 800 19440
rect 933 19410 999 19413
rect 0 19408 999 19410
rect 0 19352 938 19408
rect 994 19352 999 19408
rect 0 19350 999 19352
rect 0 19320 800 19350
rect 933 19347 999 19350
rect 28349 19410 28415 19413
rect 29200 19410 30000 19440
rect 28349 19408 30000 19410
rect 28349 19352 28354 19408
rect 28410 19352 30000 19408
rect 28349 19350 30000 19352
rect 28349 19347 28415 19350
rect 29200 19320 30000 19350
rect 1669 19274 1735 19277
rect 1534 19272 1735 19274
rect 1534 19216 1674 19272
rect 1730 19216 1735 19272
rect 1534 19214 1735 19216
rect 0 19138 800 19168
rect 1534 19138 1594 19214
rect 1669 19211 1735 19214
rect 0 19078 1594 19138
rect 0 19048 800 19078
rect 4419 19072 4735 19073
rect 4419 19008 4425 19072
rect 4489 19008 4505 19072
rect 4569 19008 4585 19072
rect 4649 19008 4665 19072
rect 4729 19008 4735 19072
rect 4419 19007 4735 19008
rect 11365 19072 11681 19073
rect 11365 19008 11371 19072
rect 11435 19008 11451 19072
rect 11515 19008 11531 19072
rect 11595 19008 11611 19072
rect 11675 19008 11681 19072
rect 11365 19007 11681 19008
rect 18311 19072 18627 19073
rect 18311 19008 18317 19072
rect 18381 19008 18397 19072
rect 18461 19008 18477 19072
rect 18541 19008 18557 19072
rect 18621 19008 18627 19072
rect 18311 19007 18627 19008
rect 25257 19072 25573 19073
rect 25257 19008 25263 19072
rect 25327 19008 25343 19072
rect 25407 19008 25423 19072
rect 25487 19008 25503 19072
rect 25567 19008 25573 19072
rect 25257 19007 25573 19008
rect 1393 19002 1459 19005
rect 936 19000 1459 19002
rect 936 18944 1398 19000
rect 1454 18944 1459 19000
rect 936 18942 1459 18944
rect 0 18866 800 18896
rect 936 18866 996 18942
rect 1393 18939 1459 18942
rect 0 18806 996 18866
rect 4061 18866 4127 18869
rect 8334 18866 8340 18868
rect 4061 18864 8340 18866
rect 4061 18808 4066 18864
rect 4122 18808 8340 18864
rect 4061 18806 8340 18808
rect 0 18776 800 18806
rect 4061 18803 4127 18806
rect 8334 18804 8340 18806
rect 8404 18804 8410 18868
rect 28809 18866 28875 18869
rect 28809 18864 29378 18866
rect 28809 18808 28814 18864
rect 28870 18808 29378 18864
rect 28809 18806 29378 18808
rect 28809 18803 28875 18806
rect 29318 18624 29378 18806
rect 0 18594 800 18624
rect 1025 18594 1091 18597
rect 0 18592 1091 18594
rect 0 18536 1030 18592
rect 1086 18536 1091 18592
rect 0 18534 1091 18536
rect 0 18504 800 18534
rect 1025 18531 1091 18534
rect 7892 18528 8208 18529
rect 7892 18464 7898 18528
rect 7962 18464 7978 18528
rect 8042 18464 8058 18528
rect 8122 18464 8138 18528
rect 8202 18464 8208 18528
rect 7892 18463 8208 18464
rect 14838 18528 15154 18529
rect 14838 18464 14844 18528
rect 14908 18464 14924 18528
rect 14988 18464 15004 18528
rect 15068 18464 15084 18528
rect 15148 18464 15154 18528
rect 14838 18463 15154 18464
rect 21784 18528 22100 18529
rect 21784 18464 21790 18528
rect 21854 18464 21870 18528
rect 21934 18464 21950 18528
rect 22014 18464 22030 18528
rect 22094 18464 22100 18528
rect 21784 18463 22100 18464
rect 28730 18528 29046 18529
rect 28730 18464 28736 18528
rect 28800 18464 28816 18528
rect 28880 18464 28896 18528
rect 28960 18464 28976 18528
rect 29040 18464 29046 18528
rect 29200 18504 30000 18624
rect 28730 18463 29046 18464
rect 0 18322 800 18352
rect 933 18322 999 18325
rect 0 18320 999 18322
rect 0 18264 938 18320
rect 994 18264 999 18320
rect 0 18262 999 18264
rect 0 18232 800 18262
rect 933 18259 999 18262
rect 0 18050 800 18080
rect 933 18050 999 18053
rect 0 18048 999 18050
rect 0 17992 938 18048
rect 994 17992 999 18048
rect 0 17990 999 17992
rect 0 17960 800 17990
rect 933 17987 999 17990
rect 4419 17984 4735 17985
rect 4419 17920 4425 17984
rect 4489 17920 4505 17984
rect 4569 17920 4585 17984
rect 4649 17920 4665 17984
rect 4729 17920 4735 17984
rect 4419 17919 4735 17920
rect 11365 17984 11681 17985
rect 11365 17920 11371 17984
rect 11435 17920 11451 17984
rect 11515 17920 11531 17984
rect 11595 17920 11611 17984
rect 11675 17920 11681 17984
rect 11365 17919 11681 17920
rect 18311 17984 18627 17985
rect 18311 17920 18317 17984
rect 18381 17920 18397 17984
rect 18461 17920 18477 17984
rect 18541 17920 18557 17984
rect 18621 17920 18627 17984
rect 18311 17919 18627 17920
rect 25257 17984 25573 17985
rect 25257 17920 25263 17984
rect 25327 17920 25343 17984
rect 25407 17920 25423 17984
rect 25487 17920 25503 17984
rect 25567 17920 25573 17984
rect 25257 17919 25573 17920
rect 1393 17914 1459 17917
rect 936 17912 1459 17914
rect 936 17856 1398 17912
rect 1454 17856 1459 17912
rect 936 17854 1459 17856
rect 0 17778 800 17808
rect 936 17778 996 17854
rect 1393 17851 1459 17854
rect 0 17718 996 17778
rect 28349 17778 28415 17781
rect 29200 17778 30000 17808
rect 28349 17776 30000 17778
rect 28349 17720 28354 17776
rect 28410 17720 30000 17776
rect 28349 17718 30000 17720
rect 0 17688 800 17718
rect 28349 17715 28415 17718
rect 29200 17688 30000 17718
rect 0 17506 800 17536
rect 933 17506 999 17509
rect 0 17504 999 17506
rect 0 17448 938 17504
rect 994 17448 999 17504
rect 0 17446 999 17448
rect 0 17416 800 17446
rect 933 17443 999 17446
rect 7892 17440 8208 17441
rect 7892 17376 7898 17440
rect 7962 17376 7978 17440
rect 8042 17376 8058 17440
rect 8122 17376 8138 17440
rect 8202 17376 8208 17440
rect 7892 17375 8208 17376
rect 14838 17440 15154 17441
rect 14838 17376 14844 17440
rect 14908 17376 14924 17440
rect 14988 17376 15004 17440
rect 15068 17376 15084 17440
rect 15148 17376 15154 17440
rect 14838 17375 15154 17376
rect 21784 17440 22100 17441
rect 21784 17376 21790 17440
rect 21854 17376 21870 17440
rect 21934 17376 21950 17440
rect 22014 17376 22030 17440
rect 22094 17376 22100 17440
rect 21784 17375 22100 17376
rect 28730 17440 29046 17441
rect 28730 17376 28736 17440
rect 28800 17376 28816 17440
rect 28880 17376 28896 17440
rect 28960 17376 28976 17440
rect 29040 17376 29046 17440
rect 28730 17375 29046 17376
rect 0 17234 800 17264
rect 1025 17234 1091 17237
rect 0 17232 1091 17234
rect 0 17176 1030 17232
rect 1086 17176 1091 17232
rect 0 17174 1091 17176
rect 0 17144 800 17174
rect 1025 17171 1091 17174
rect 0 16962 800 16992
rect 933 16962 999 16965
rect 0 16960 999 16962
rect 0 16904 938 16960
rect 994 16904 999 16960
rect 0 16902 999 16904
rect 0 16872 800 16902
rect 933 16899 999 16902
rect 28349 16962 28415 16965
rect 29200 16962 30000 16992
rect 28349 16960 30000 16962
rect 28349 16904 28354 16960
rect 28410 16904 30000 16960
rect 28349 16902 30000 16904
rect 28349 16899 28415 16902
rect 4419 16896 4735 16897
rect 4419 16832 4425 16896
rect 4489 16832 4505 16896
rect 4569 16832 4585 16896
rect 4649 16832 4665 16896
rect 4729 16832 4735 16896
rect 4419 16831 4735 16832
rect 11365 16896 11681 16897
rect 11365 16832 11371 16896
rect 11435 16832 11451 16896
rect 11515 16832 11531 16896
rect 11595 16832 11611 16896
rect 11675 16832 11681 16896
rect 11365 16831 11681 16832
rect 18311 16896 18627 16897
rect 18311 16832 18317 16896
rect 18381 16832 18397 16896
rect 18461 16832 18477 16896
rect 18541 16832 18557 16896
rect 18621 16832 18627 16896
rect 18311 16831 18627 16832
rect 25257 16896 25573 16897
rect 25257 16832 25263 16896
rect 25327 16832 25343 16896
rect 25407 16832 25423 16896
rect 25487 16832 25503 16896
rect 25567 16832 25573 16896
rect 29200 16872 30000 16902
rect 25257 16831 25573 16832
rect 0 16690 800 16720
rect 1025 16690 1091 16693
rect 0 16688 1091 16690
rect 0 16632 1030 16688
rect 1086 16632 1091 16688
rect 0 16630 1091 16632
rect 0 16600 800 16630
rect 1025 16627 1091 16630
rect 0 16418 800 16448
rect 933 16418 999 16421
rect 0 16416 999 16418
rect 0 16360 938 16416
rect 994 16360 999 16416
rect 0 16358 999 16360
rect 0 16328 800 16358
rect 933 16355 999 16358
rect 7892 16352 8208 16353
rect 7892 16288 7898 16352
rect 7962 16288 7978 16352
rect 8042 16288 8058 16352
rect 8122 16288 8138 16352
rect 8202 16288 8208 16352
rect 7892 16287 8208 16288
rect 14838 16352 15154 16353
rect 14838 16288 14844 16352
rect 14908 16288 14924 16352
rect 14988 16288 15004 16352
rect 15068 16288 15084 16352
rect 15148 16288 15154 16352
rect 14838 16287 15154 16288
rect 21784 16352 22100 16353
rect 21784 16288 21790 16352
rect 21854 16288 21870 16352
rect 21934 16288 21950 16352
rect 22014 16288 22030 16352
rect 22094 16288 22100 16352
rect 21784 16287 22100 16288
rect 28730 16352 29046 16353
rect 28730 16288 28736 16352
rect 28800 16288 28816 16352
rect 28880 16288 28896 16352
rect 28960 16288 28976 16352
rect 29040 16288 29046 16352
rect 28730 16287 29046 16288
rect 0 16146 800 16176
rect 1025 16146 1091 16149
rect 0 16144 1091 16146
rect 0 16088 1030 16144
rect 1086 16088 1091 16144
rect 0 16086 1091 16088
rect 0 16056 800 16086
rect 1025 16083 1091 16086
rect 28349 16146 28415 16149
rect 29200 16146 30000 16176
rect 28349 16144 30000 16146
rect 28349 16088 28354 16144
rect 28410 16088 30000 16144
rect 28349 16086 30000 16088
rect 28349 16083 28415 16086
rect 29200 16056 30000 16086
rect 0 15874 800 15904
rect 933 15874 999 15877
rect 0 15872 999 15874
rect 0 15816 938 15872
rect 994 15816 999 15872
rect 0 15814 999 15816
rect 0 15784 800 15814
rect 933 15811 999 15814
rect 4419 15808 4735 15809
rect 4419 15744 4425 15808
rect 4489 15744 4505 15808
rect 4569 15744 4585 15808
rect 4649 15744 4665 15808
rect 4729 15744 4735 15808
rect 4419 15743 4735 15744
rect 11365 15808 11681 15809
rect 11365 15744 11371 15808
rect 11435 15744 11451 15808
rect 11515 15744 11531 15808
rect 11595 15744 11611 15808
rect 11675 15744 11681 15808
rect 11365 15743 11681 15744
rect 18311 15808 18627 15809
rect 18311 15744 18317 15808
rect 18381 15744 18397 15808
rect 18461 15744 18477 15808
rect 18541 15744 18557 15808
rect 18621 15744 18627 15808
rect 18311 15743 18627 15744
rect 25257 15808 25573 15809
rect 25257 15744 25263 15808
rect 25327 15744 25343 15808
rect 25407 15744 25423 15808
rect 25487 15744 25503 15808
rect 25567 15744 25573 15808
rect 25257 15743 25573 15744
rect 0 15602 800 15632
rect 1025 15602 1091 15605
rect 0 15600 1091 15602
rect 0 15544 1030 15600
rect 1086 15544 1091 15600
rect 0 15542 1091 15544
rect 0 15512 800 15542
rect 1025 15539 1091 15542
rect 28352 15406 29194 15466
rect 0 15330 800 15360
rect 28352 15333 28412 15406
rect 29134 15364 29194 15406
rect 29134 15360 29378 15364
rect 933 15330 999 15333
rect 0 15328 999 15330
rect 0 15272 938 15328
rect 994 15272 999 15328
rect 0 15270 999 15272
rect 0 15240 800 15270
rect 933 15267 999 15270
rect 1669 15330 1735 15333
rect 4102 15330 4108 15332
rect 1669 15328 4108 15330
rect 1669 15272 1674 15328
rect 1730 15272 4108 15328
rect 1669 15270 4108 15272
rect 1669 15267 1735 15270
rect 4102 15268 4108 15270
rect 4172 15268 4178 15332
rect 28349 15328 28415 15333
rect 28349 15272 28354 15328
rect 28410 15272 28415 15328
rect 29134 15304 30000 15360
rect 28349 15267 28415 15272
rect 7892 15264 8208 15265
rect 7892 15200 7898 15264
rect 7962 15200 7978 15264
rect 8042 15200 8058 15264
rect 8122 15200 8138 15264
rect 8202 15200 8208 15264
rect 7892 15199 8208 15200
rect 14838 15264 15154 15265
rect 14838 15200 14844 15264
rect 14908 15200 14924 15264
rect 14988 15200 15004 15264
rect 15068 15200 15084 15264
rect 15148 15200 15154 15264
rect 14838 15199 15154 15200
rect 21784 15264 22100 15265
rect 21784 15200 21790 15264
rect 21854 15200 21870 15264
rect 21934 15200 21950 15264
rect 22014 15200 22030 15264
rect 22094 15200 22100 15264
rect 21784 15199 22100 15200
rect 28730 15264 29046 15265
rect 28730 15200 28736 15264
rect 28800 15200 28816 15264
rect 28880 15200 28896 15264
rect 28960 15200 28976 15264
rect 29040 15200 29046 15264
rect 29200 15240 30000 15304
rect 28730 15199 29046 15200
rect 1853 15194 1919 15197
rect 936 15192 1919 15194
rect 936 15136 1858 15192
rect 1914 15136 1919 15192
rect 936 15134 1919 15136
rect 0 15058 800 15088
rect 936 15058 996 15134
rect 1853 15131 1919 15134
rect 0 14998 996 15058
rect 0 14968 800 14998
rect 0 14696 800 14816
rect 4419 14720 4735 14721
rect 4419 14656 4425 14720
rect 4489 14656 4505 14720
rect 4569 14656 4585 14720
rect 4649 14656 4665 14720
rect 4729 14656 4735 14720
rect 4419 14655 4735 14656
rect 11365 14720 11681 14721
rect 11365 14656 11371 14720
rect 11435 14656 11451 14720
rect 11515 14656 11531 14720
rect 11595 14656 11611 14720
rect 11675 14656 11681 14720
rect 11365 14655 11681 14656
rect 18311 14720 18627 14721
rect 18311 14656 18317 14720
rect 18381 14656 18397 14720
rect 18461 14656 18477 14720
rect 18541 14656 18557 14720
rect 18621 14656 18627 14720
rect 18311 14655 18627 14656
rect 25257 14720 25573 14721
rect 25257 14656 25263 14720
rect 25327 14656 25343 14720
rect 25407 14656 25423 14720
rect 25487 14656 25503 14720
rect 25567 14656 25573 14720
rect 25257 14655 25573 14656
rect 0 14514 800 14544
rect 933 14514 999 14517
rect 0 14512 999 14514
rect 0 14456 938 14512
rect 994 14456 999 14512
rect 0 14454 999 14456
rect 0 14424 800 14454
rect 933 14451 999 14454
rect 10041 14514 10107 14517
rect 26969 14514 27035 14517
rect 10041 14512 27035 14514
rect 10041 14456 10046 14512
rect 10102 14456 26974 14512
rect 27030 14456 27035 14512
rect 10041 14454 27035 14456
rect 10041 14451 10107 14454
rect 26969 14451 27035 14454
rect 28349 14514 28415 14517
rect 29200 14514 30000 14544
rect 28349 14512 30000 14514
rect 28349 14456 28354 14512
rect 28410 14456 30000 14512
rect 28349 14454 30000 14456
rect 28349 14451 28415 14454
rect 29200 14424 30000 14454
rect 1853 14378 1919 14381
rect 13721 14378 13787 14381
rect 1853 14376 13787 14378
rect 1853 14320 1858 14376
rect 1914 14320 13726 14376
rect 13782 14320 13787 14376
rect 1853 14318 13787 14320
rect 1853 14315 1919 14318
rect 13721 14315 13787 14318
rect 0 14242 800 14272
rect 933 14242 999 14245
rect 0 14240 999 14242
rect 0 14184 938 14240
rect 994 14184 999 14240
rect 0 14182 999 14184
rect 0 14152 800 14182
rect 933 14179 999 14182
rect 7892 14176 8208 14177
rect 7892 14112 7898 14176
rect 7962 14112 7978 14176
rect 8042 14112 8058 14176
rect 8122 14112 8138 14176
rect 8202 14112 8208 14176
rect 7892 14111 8208 14112
rect 14838 14176 15154 14177
rect 14838 14112 14844 14176
rect 14908 14112 14924 14176
rect 14988 14112 15004 14176
rect 15068 14112 15084 14176
rect 15148 14112 15154 14176
rect 14838 14111 15154 14112
rect 21784 14176 22100 14177
rect 21784 14112 21790 14176
rect 21854 14112 21870 14176
rect 21934 14112 21950 14176
rect 22014 14112 22030 14176
rect 22094 14112 22100 14176
rect 21784 14111 22100 14112
rect 28730 14176 29046 14177
rect 28730 14112 28736 14176
rect 28800 14112 28816 14176
rect 28880 14112 28896 14176
rect 28960 14112 28976 14176
rect 29040 14112 29046 14176
rect 28730 14111 29046 14112
rect 0 13970 800 14000
rect 1025 13970 1091 13973
rect 0 13968 1091 13970
rect 0 13912 1030 13968
rect 1086 13912 1091 13968
rect 0 13910 1091 13912
rect 0 13880 800 13910
rect 1025 13907 1091 13910
rect 1853 13834 1919 13837
rect 16113 13834 16179 13837
rect 1853 13832 16179 13834
rect 1853 13776 1858 13832
rect 1914 13776 16118 13832
rect 16174 13776 16179 13832
rect 1853 13774 16179 13776
rect 1853 13771 1919 13774
rect 16113 13771 16179 13774
rect 0 13698 800 13728
rect 1393 13698 1459 13701
rect 1669 13698 1735 13701
rect 8385 13700 8451 13701
rect 8334 13698 8340 13700
rect 0 13696 1459 13698
rect 0 13640 1398 13696
rect 1454 13640 1459 13696
rect 0 13638 1459 13640
rect 0 13608 800 13638
rect 1393 13635 1459 13638
rect 1534 13696 1735 13698
rect 1534 13640 1674 13696
rect 1730 13640 1735 13696
rect 1534 13638 1735 13640
rect 8294 13638 8340 13698
rect 8404 13696 8451 13700
rect 8446 13640 8451 13696
rect 0 13426 800 13456
rect 1534 13426 1594 13638
rect 1669 13635 1735 13638
rect 8334 13636 8340 13638
rect 8404 13636 8451 13640
rect 8385 13635 8451 13636
rect 28349 13698 28415 13701
rect 29200 13698 30000 13728
rect 28349 13696 30000 13698
rect 28349 13640 28354 13696
rect 28410 13640 30000 13696
rect 28349 13638 30000 13640
rect 28349 13635 28415 13638
rect 4419 13632 4735 13633
rect 4419 13568 4425 13632
rect 4489 13568 4505 13632
rect 4569 13568 4585 13632
rect 4649 13568 4665 13632
rect 4729 13568 4735 13632
rect 4419 13567 4735 13568
rect 11365 13632 11681 13633
rect 11365 13568 11371 13632
rect 11435 13568 11451 13632
rect 11515 13568 11531 13632
rect 11595 13568 11611 13632
rect 11675 13568 11681 13632
rect 11365 13567 11681 13568
rect 18311 13632 18627 13633
rect 18311 13568 18317 13632
rect 18381 13568 18397 13632
rect 18461 13568 18477 13632
rect 18541 13568 18557 13632
rect 18621 13568 18627 13632
rect 18311 13567 18627 13568
rect 25257 13632 25573 13633
rect 25257 13568 25263 13632
rect 25327 13568 25343 13632
rect 25407 13568 25423 13632
rect 25487 13568 25503 13632
rect 25567 13568 25573 13632
rect 29200 13608 30000 13638
rect 25257 13567 25573 13568
rect 0 13366 1594 13426
rect 1853 13426 1919 13429
rect 15285 13426 15351 13429
rect 1853 13424 15351 13426
rect 1853 13368 1858 13424
rect 1914 13368 15290 13424
rect 15346 13368 15351 13424
rect 1853 13366 15351 13368
rect 0 13336 800 13366
rect 1853 13363 1919 13366
rect 15285 13363 15351 13366
rect 1577 13290 1643 13293
rect 15745 13290 15811 13293
rect 1577 13288 15811 13290
rect 1577 13232 1582 13288
rect 1638 13232 15750 13288
rect 15806 13232 15811 13288
rect 1577 13230 15811 13232
rect 1577 13227 1643 13230
rect 15745 13227 15811 13230
rect 0 13154 800 13184
rect 933 13154 999 13157
rect 0 13152 999 13154
rect 0 13096 938 13152
rect 994 13096 999 13152
rect 0 13094 999 13096
rect 0 13064 800 13094
rect 933 13091 999 13094
rect 7892 13088 8208 13089
rect 7892 13024 7898 13088
rect 7962 13024 7978 13088
rect 8042 13024 8058 13088
rect 8122 13024 8138 13088
rect 8202 13024 8208 13088
rect 7892 13023 8208 13024
rect 14838 13088 15154 13089
rect 14838 13024 14844 13088
rect 14908 13024 14924 13088
rect 14988 13024 15004 13088
rect 15068 13024 15084 13088
rect 15148 13024 15154 13088
rect 14838 13023 15154 13024
rect 21784 13088 22100 13089
rect 21784 13024 21790 13088
rect 21854 13024 21870 13088
rect 21934 13024 21950 13088
rect 22014 13024 22030 13088
rect 22094 13024 22100 13088
rect 21784 13023 22100 13024
rect 28730 13088 29046 13089
rect 28730 13024 28736 13088
rect 28800 13024 28816 13088
rect 28880 13024 28896 13088
rect 28960 13024 28976 13088
rect 29040 13024 29046 13088
rect 28730 13023 29046 13024
rect 0 12882 800 12912
rect 1025 12882 1091 12885
rect 0 12880 1091 12882
rect 0 12824 1030 12880
rect 1086 12824 1091 12880
rect 0 12822 1091 12824
rect 0 12792 800 12822
rect 1025 12819 1091 12822
rect 8017 12882 8083 12885
rect 9581 12882 9647 12885
rect 8017 12880 9647 12882
rect 8017 12824 8022 12880
rect 8078 12824 9586 12880
rect 9642 12824 9647 12880
rect 8017 12822 9647 12824
rect 8017 12819 8083 12822
rect 9581 12819 9647 12822
rect 28349 12882 28415 12885
rect 29200 12882 30000 12912
rect 28349 12880 30000 12882
rect 28349 12824 28354 12880
rect 28410 12824 30000 12880
rect 28349 12822 30000 12824
rect 28349 12819 28415 12822
rect 29200 12792 30000 12822
rect 1853 12746 1919 12749
rect 13721 12746 13787 12749
rect 1853 12744 13787 12746
rect 1853 12688 1858 12744
rect 1914 12688 13726 12744
rect 13782 12688 13787 12744
rect 1853 12686 13787 12688
rect 1853 12683 1919 12686
rect 13721 12683 13787 12686
rect 0 12610 800 12640
rect 933 12610 999 12613
rect 0 12608 999 12610
rect 0 12552 938 12608
rect 994 12552 999 12608
rect 0 12550 999 12552
rect 0 12520 800 12550
rect 933 12547 999 12550
rect 4419 12544 4735 12545
rect 4419 12480 4425 12544
rect 4489 12480 4505 12544
rect 4569 12480 4585 12544
rect 4649 12480 4665 12544
rect 4729 12480 4735 12544
rect 4419 12479 4735 12480
rect 11365 12544 11681 12545
rect 11365 12480 11371 12544
rect 11435 12480 11451 12544
rect 11515 12480 11531 12544
rect 11595 12480 11611 12544
rect 11675 12480 11681 12544
rect 11365 12479 11681 12480
rect 18311 12544 18627 12545
rect 18311 12480 18317 12544
rect 18381 12480 18397 12544
rect 18461 12480 18477 12544
rect 18541 12480 18557 12544
rect 18621 12480 18627 12544
rect 18311 12479 18627 12480
rect 25257 12544 25573 12545
rect 25257 12480 25263 12544
rect 25327 12480 25343 12544
rect 25407 12480 25423 12544
rect 25487 12480 25503 12544
rect 25567 12480 25573 12544
rect 25257 12479 25573 12480
rect 7925 12474 7991 12477
rect 8753 12474 8819 12477
rect 7925 12472 8819 12474
rect 7925 12416 7930 12472
rect 7986 12416 8758 12472
rect 8814 12416 8819 12472
rect 7925 12414 8819 12416
rect 7925 12411 7991 12414
rect 8753 12411 8819 12414
rect 0 12338 800 12368
rect 1669 12338 1735 12341
rect 0 12336 1735 12338
rect 0 12280 1674 12336
rect 1730 12280 1735 12336
rect 0 12278 1735 12280
rect 0 12248 800 12278
rect 1669 12275 1735 12278
rect 9765 12338 9831 12341
rect 15561 12338 15627 12341
rect 9765 12336 15627 12338
rect 9765 12280 9770 12336
rect 9826 12280 15566 12336
rect 15622 12280 15627 12336
rect 9765 12278 15627 12280
rect 9765 12275 9831 12278
rect 15561 12275 15627 12278
rect 1853 12202 1919 12205
rect 17125 12202 17191 12205
rect 1853 12200 17191 12202
rect 1853 12144 1858 12200
rect 1914 12144 17130 12200
rect 17186 12144 17191 12200
rect 1853 12142 17191 12144
rect 1853 12139 1919 12142
rect 17125 12139 17191 12142
rect 28352 12142 29194 12202
rect 0 12066 800 12096
rect 28352 12069 28412 12142
rect 29134 12100 29194 12142
rect 29134 12096 29378 12100
rect 933 12066 999 12069
rect 0 12064 999 12066
rect 0 12008 938 12064
rect 994 12008 999 12064
rect 0 12006 999 12008
rect 0 11976 800 12006
rect 933 12003 999 12006
rect 28349 12064 28415 12069
rect 28349 12008 28354 12064
rect 28410 12008 28415 12064
rect 29134 12040 30000 12096
rect 28349 12003 28415 12008
rect 7892 12000 8208 12001
rect 7892 11936 7898 12000
rect 7962 11936 7978 12000
rect 8042 11936 8058 12000
rect 8122 11936 8138 12000
rect 8202 11936 8208 12000
rect 7892 11935 8208 11936
rect 14838 12000 15154 12001
rect 14838 11936 14844 12000
rect 14908 11936 14924 12000
rect 14988 11936 15004 12000
rect 15068 11936 15084 12000
rect 15148 11936 15154 12000
rect 14838 11935 15154 11936
rect 21784 12000 22100 12001
rect 21784 11936 21790 12000
rect 21854 11936 21870 12000
rect 21934 11936 21950 12000
rect 22014 11936 22030 12000
rect 22094 11936 22100 12000
rect 21784 11935 22100 11936
rect 28730 12000 29046 12001
rect 28730 11936 28736 12000
rect 28800 11936 28816 12000
rect 28880 11936 28896 12000
rect 28960 11936 28976 12000
rect 29040 11936 29046 12000
rect 29200 11976 30000 12040
rect 28730 11935 29046 11936
rect 0 11794 800 11824
rect 1025 11794 1091 11797
rect 0 11792 1091 11794
rect 0 11736 1030 11792
rect 1086 11736 1091 11792
rect 0 11734 1091 11736
rect 0 11704 800 11734
rect 1025 11731 1091 11734
rect 5165 11794 5231 11797
rect 7925 11794 7991 11797
rect 15929 11794 15995 11797
rect 5165 11792 15995 11794
rect 5165 11736 5170 11792
rect 5226 11736 7930 11792
rect 7986 11736 15934 11792
rect 15990 11736 15995 11792
rect 5165 11734 15995 11736
rect 5165 11731 5231 11734
rect 7925 11731 7991 11734
rect 15929 11731 15995 11734
rect 0 11522 800 11552
rect 933 11522 999 11525
rect 0 11520 999 11522
rect 0 11464 938 11520
rect 994 11464 999 11520
rect 0 11462 999 11464
rect 0 11432 800 11462
rect 933 11459 999 11462
rect 4419 11456 4735 11457
rect 4419 11392 4425 11456
rect 4489 11392 4505 11456
rect 4569 11392 4585 11456
rect 4649 11392 4665 11456
rect 4729 11392 4735 11456
rect 4419 11391 4735 11392
rect 11365 11456 11681 11457
rect 11365 11392 11371 11456
rect 11435 11392 11451 11456
rect 11515 11392 11531 11456
rect 11595 11392 11611 11456
rect 11675 11392 11681 11456
rect 11365 11391 11681 11392
rect 18311 11456 18627 11457
rect 18311 11392 18317 11456
rect 18381 11392 18397 11456
rect 18461 11392 18477 11456
rect 18541 11392 18557 11456
rect 18621 11392 18627 11456
rect 18311 11391 18627 11392
rect 25257 11456 25573 11457
rect 25257 11392 25263 11456
rect 25327 11392 25343 11456
rect 25407 11392 25423 11456
rect 25487 11392 25503 11456
rect 25567 11392 25573 11456
rect 25257 11391 25573 11392
rect 8845 11386 8911 11389
rect 9581 11386 9647 11389
rect 8845 11384 9647 11386
rect 8845 11328 8850 11384
rect 8906 11328 9586 11384
rect 9642 11328 9647 11384
rect 8845 11326 9647 11328
rect 8845 11323 8911 11326
rect 9581 11323 9647 11326
rect 0 11250 800 11280
rect 1025 11250 1091 11253
rect 0 11248 1091 11250
rect 0 11192 1030 11248
rect 1086 11192 1091 11248
rect 0 11190 1091 11192
rect 0 11160 800 11190
rect 1025 11187 1091 11190
rect 11513 11250 11579 11253
rect 11973 11250 12039 11253
rect 11513 11248 12039 11250
rect 11513 11192 11518 11248
rect 11574 11192 11978 11248
rect 12034 11192 12039 11248
rect 11513 11190 12039 11192
rect 11513 11187 11579 11190
rect 11973 11187 12039 11190
rect 28349 11250 28415 11253
rect 29200 11250 30000 11280
rect 28349 11248 30000 11250
rect 28349 11192 28354 11248
rect 28410 11192 30000 11248
rect 28349 11190 30000 11192
rect 28349 11187 28415 11190
rect 29200 11160 30000 11190
rect 0 10978 800 11008
rect 1393 10978 1459 10981
rect 1669 10978 1735 10981
rect 0 10976 1459 10978
rect 0 10920 1398 10976
rect 1454 10920 1459 10976
rect 0 10918 1459 10920
rect 0 10888 800 10918
rect 1393 10915 1459 10918
rect 1534 10976 1735 10978
rect 1534 10920 1674 10976
rect 1730 10920 1735 10976
rect 1534 10918 1735 10920
rect 0 10706 800 10736
rect 1534 10706 1594 10918
rect 1669 10915 1735 10918
rect 7892 10912 8208 10913
rect 7892 10848 7898 10912
rect 7962 10848 7978 10912
rect 8042 10848 8058 10912
rect 8122 10848 8138 10912
rect 8202 10848 8208 10912
rect 7892 10847 8208 10848
rect 14838 10912 15154 10913
rect 14838 10848 14844 10912
rect 14908 10848 14924 10912
rect 14988 10848 15004 10912
rect 15068 10848 15084 10912
rect 15148 10848 15154 10912
rect 14838 10847 15154 10848
rect 21784 10912 22100 10913
rect 21784 10848 21790 10912
rect 21854 10848 21870 10912
rect 21934 10848 21950 10912
rect 22014 10848 22030 10912
rect 22094 10848 22100 10912
rect 21784 10847 22100 10848
rect 28730 10912 29046 10913
rect 28730 10848 28736 10912
rect 28800 10848 28816 10912
rect 28880 10848 28896 10912
rect 28960 10848 28976 10912
rect 29040 10848 29046 10912
rect 28730 10847 29046 10848
rect 0 10646 1594 10706
rect 0 10616 800 10646
rect 1577 10570 1643 10573
rect 15929 10570 15995 10573
rect 1577 10568 15995 10570
rect 1577 10512 1582 10568
rect 1638 10512 15934 10568
rect 15990 10512 15995 10568
rect 1577 10510 15995 10512
rect 1577 10507 1643 10510
rect 15929 10507 15995 10510
rect 0 10434 800 10464
rect 933 10434 999 10437
rect 0 10432 999 10434
rect 0 10376 938 10432
rect 994 10376 999 10432
rect 0 10374 999 10376
rect 0 10344 800 10374
rect 933 10371 999 10374
rect 28349 10434 28415 10437
rect 29200 10434 30000 10464
rect 28349 10432 30000 10434
rect 28349 10376 28354 10432
rect 28410 10376 30000 10432
rect 28349 10374 30000 10376
rect 28349 10371 28415 10374
rect 4419 10368 4735 10369
rect 4419 10304 4425 10368
rect 4489 10304 4505 10368
rect 4569 10304 4585 10368
rect 4649 10304 4665 10368
rect 4729 10304 4735 10368
rect 4419 10303 4735 10304
rect 11365 10368 11681 10369
rect 11365 10304 11371 10368
rect 11435 10304 11451 10368
rect 11515 10304 11531 10368
rect 11595 10304 11611 10368
rect 11675 10304 11681 10368
rect 11365 10303 11681 10304
rect 18311 10368 18627 10369
rect 18311 10304 18317 10368
rect 18381 10304 18397 10368
rect 18461 10304 18477 10368
rect 18541 10304 18557 10368
rect 18621 10304 18627 10368
rect 18311 10303 18627 10304
rect 25257 10368 25573 10369
rect 25257 10304 25263 10368
rect 25327 10304 25343 10368
rect 25407 10304 25423 10368
rect 25487 10304 25503 10368
rect 25567 10304 25573 10368
rect 29200 10344 30000 10374
rect 25257 10303 25573 10304
rect 0 10162 800 10192
rect 1025 10162 1091 10165
rect 0 10160 1091 10162
rect 0 10104 1030 10160
rect 1086 10104 1091 10160
rect 0 10102 1091 10104
rect 0 10072 800 10102
rect 1025 10099 1091 10102
rect 4797 10026 4863 10029
rect 5717 10026 5783 10029
rect 4797 10024 5783 10026
rect 4797 9968 4802 10024
rect 4858 9968 5722 10024
rect 5778 9968 5783 10024
rect 4797 9966 5783 9968
rect 4797 9963 4863 9966
rect 5717 9963 5783 9966
rect 0 9890 800 9920
rect 933 9890 999 9893
rect 0 9888 999 9890
rect 0 9832 938 9888
rect 994 9832 999 9888
rect 0 9830 999 9832
rect 0 9800 800 9830
rect 933 9827 999 9830
rect 7892 9824 8208 9825
rect 7892 9760 7898 9824
rect 7962 9760 7978 9824
rect 8042 9760 8058 9824
rect 8122 9760 8138 9824
rect 8202 9760 8208 9824
rect 7892 9759 8208 9760
rect 14838 9824 15154 9825
rect 14838 9760 14844 9824
rect 14908 9760 14924 9824
rect 14988 9760 15004 9824
rect 15068 9760 15084 9824
rect 15148 9760 15154 9824
rect 14838 9759 15154 9760
rect 21784 9824 22100 9825
rect 21784 9760 21790 9824
rect 21854 9760 21870 9824
rect 21934 9760 21950 9824
rect 22014 9760 22030 9824
rect 22094 9760 22100 9824
rect 21784 9759 22100 9760
rect 28730 9824 29046 9825
rect 28730 9760 28736 9824
rect 28800 9760 28816 9824
rect 28880 9760 28896 9824
rect 28960 9760 28976 9824
rect 29040 9760 29046 9824
rect 28730 9759 29046 9760
rect 0 9618 800 9648
rect 1669 9618 1735 9621
rect 0 9616 1735 9618
rect 0 9560 1674 9616
rect 1730 9560 1735 9616
rect 0 9558 1735 9560
rect 0 9528 800 9558
rect 1669 9555 1735 9558
rect 4613 9618 4679 9621
rect 5073 9618 5139 9621
rect 4613 9616 5139 9618
rect 4613 9560 4618 9616
rect 4674 9560 5078 9616
rect 5134 9560 5139 9616
rect 4613 9558 5139 9560
rect 4613 9555 4679 9558
rect 5073 9555 5139 9558
rect 10409 9618 10475 9621
rect 14181 9618 14247 9621
rect 10409 9616 14247 9618
rect 10409 9560 10414 9616
rect 10470 9560 14186 9616
rect 14242 9560 14247 9616
rect 10409 9558 14247 9560
rect 10409 9555 10475 9558
rect 14181 9555 14247 9558
rect 28349 9618 28415 9621
rect 29200 9618 30000 9648
rect 28349 9616 30000 9618
rect 28349 9560 28354 9616
rect 28410 9560 30000 9616
rect 28349 9558 30000 9560
rect 28349 9555 28415 9558
rect 29200 9528 30000 9558
rect 10041 9482 10107 9485
rect 10501 9482 10567 9485
rect 10041 9480 10567 9482
rect 10041 9424 10046 9480
rect 10102 9424 10506 9480
rect 10562 9424 10567 9480
rect 10041 9422 10567 9424
rect 10041 9419 10107 9422
rect 10501 9419 10567 9422
rect 0 9346 800 9376
rect 933 9346 999 9349
rect 0 9344 999 9346
rect 0 9288 938 9344
rect 994 9288 999 9344
rect 0 9286 999 9288
rect 0 9256 800 9286
rect 933 9283 999 9286
rect 4419 9280 4735 9281
rect 4419 9216 4425 9280
rect 4489 9216 4505 9280
rect 4569 9216 4585 9280
rect 4649 9216 4665 9280
rect 4729 9216 4735 9280
rect 4419 9215 4735 9216
rect 11365 9280 11681 9281
rect 11365 9216 11371 9280
rect 11435 9216 11451 9280
rect 11515 9216 11531 9280
rect 11595 9216 11611 9280
rect 11675 9216 11681 9280
rect 11365 9215 11681 9216
rect 18311 9280 18627 9281
rect 18311 9216 18317 9280
rect 18381 9216 18397 9280
rect 18461 9216 18477 9280
rect 18541 9216 18557 9280
rect 18621 9216 18627 9280
rect 18311 9215 18627 9216
rect 25257 9280 25573 9281
rect 25257 9216 25263 9280
rect 25327 9216 25343 9280
rect 25407 9216 25423 9280
rect 25487 9216 25503 9280
rect 25567 9216 25573 9280
rect 25257 9215 25573 9216
rect 5349 9212 5415 9213
rect 5349 9208 5396 9212
rect 5460 9210 5466 9212
rect 5349 9152 5354 9208
rect 5349 9148 5396 9152
rect 5460 9150 5506 9210
rect 5460 9148 5466 9150
rect 5349 9147 5415 9148
rect 0 9074 800 9104
rect 1025 9074 1091 9077
rect 0 9072 1091 9074
rect 0 9016 1030 9072
rect 1086 9016 1091 9072
rect 0 9014 1091 9016
rect 0 8984 800 9014
rect 1025 9011 1091 9014
rect 9765 9074 9831 9077
rect 10593 9074 10659 9077
rect 9765 9072 10659 9074
rect 9765 9016 9770 9072
rect 9826 9016 10598 9072
rect 10654 9016 10659 9072
rect 9765 9014 10659 9016
rect 9765 9011 9831 9014
rect 10593 9011 10659 9014
rect 28809 9074 28875 9077
rect 28809 9072 29378 9074
rect 28809 9016 28814 9072
rect 28870 9016 29378 9072
rect 28809 9014 29378 9016
rect 28809 9011 28875 9014
rect 2129 8938 2195 8941
rect 8477 8938 8543 8941
rect 2129 8936 8543 8938
rect 2129 8880 2134 8936
rect 2190 8880 8482 8936
rect 8538 8880 8543 8936
rect 2129 8878 8543 8880
rect 2129 8875 2195 8878
rect 8477 8875 8543 8878
rect 29318 8832 29378 9014
rect 0 8802 800 8832
rect 933 8802 999 8805
rect 0 8800 999 8802
rect 0 8744 938 8800
rect 994 8744 999 8800
rect 0 8742 999 8744
rect 0 8712 800 8742
rect 933 8739 999 8742
rect 1577 8802 1643 8805
rect 6637 8802 6703 8805
rect 1577 8800 6703 8802
rect 1577 8744 1582 8800
rect 1638 8744 6642 8800
rect 6698 8744 6703 8800
rect 1577 8742 6703 8744
rect 1577 8739 1643 8742
rect 6637 8739 6703 8742
rect 7892 8736 8208 8737
rect 7892 8672 7898 8736
rect 7962 8672 7978 8736
rect 8042 8672 8058 8736
rect 8122 8672 8138 8736
rect 8202 8672 8208 8736
rect 7892 8671 8208 8672
rect 14838 8736 15154 8737
rect 14838 8672 14844 8736
rect 14908 8672 14924 8736
rect 14988 8672 15004 8736
rect 15068 8672 15084 8736
rect 15148 8672 15154 8736
rect 14838 8671 15154 8672
rect 21784 8736 22100 8737
rect 21784 8672 21790 8736
rect 21854 8672 21870 8736
rect 21934 8672 21950 8736
rect 22014 8672 22030 8736
rect 22094 8672 22100 8736
rect 21784 8671 22100 8672
rect 28730 8736 29046 8737
rect 28730 8672 28736 8736
rect 28800 8672 28816 8736
rect 28880 8672 28896 8736
rect 28960 8672 28976 8736
rect 29040 8672 29046 8736
rect 29200 8712 30000 8832
rect 28730 8671 29046 8672
rect 2405 8666 2471 8669
rect 7557 8666 7623 8669
rect 2405 8664 7623 8666
rect 2405 8608 2410 8664
rect 2466 8608 7562 8664
rect 7618 8608 7623 8664
rect 2405 8606 7623 8608
rect 2405 8603 2471 8606
rect 7557 8603 7623 8606
rect 0 8530 800 8560
rect 1025 8530 1091 8533
rect 0 8528 1091 8530
rect 0 8472 1030 8528
rect 1086 8472 1091 8528
rect 0 8470 1091 8472
rect 0 8440 800 8470
rect 1025 8467 1091 8470
rect 1577 8530 1643 8533
rect 8293 8530 8359 8533
rect 1577 8528 8359 8530
rect 1577 8472 1582 8528
rect 1638 8472 8298 8528
rect 8354 8472 8359 8528
rect 1577 8470 8359 8472
rect 1577 8467 1643 8470
rect 8293 8467 8359 8470
rect 1025 8394 1091 8397
rect 6545 8394 6611 8397
rect 1025 8392 6611 8394
rect 1025 8336 1030 8392
rect 1086 8336 6550 8392
rect 6606 8336 6611 8392
rect 1025 8334 6611 8336
rect 1025 8331 1091 8334
rect 6545 8331 6611 8334
rect 0 8258 800 8288
rect 1393 8258 1459 8261
rect 1669 8258 1735 8261
rect 0 8256 1459 8258
rect 0 8200 1398 8256
rect 1454 8200 1459 8256
rect 0 8198 1459 8200
rect 0 8168 800 8198
rect 1393 8195 1459 8198
rect 1534 8256 1735 8258
rect 1534 8200 1674 8256
rect 1730 8200 1735 8256
rect 1534 8198 1735 8200
rect 0 7986 800 8016
rect 1534 7986 1594 8198
rect 1669 8195 1735 8198
rect 4419 8192 4735 8193
rect 4419 8128 4425 8192
rect 4489 8128 4505 8192
rect 4569 8128 4585 8192
rect 4649 8128 4665 8192
rect 4729 8128 4735 8192
rect 4419 8127 4735 8128
rect 11365 8192 11681 8193
rect 11365 8128 11371 8192
rect 11435 8128 11451 8192
rect 11515 8128 11531 8192
rect 11595 8128 11611 8192
rect 11675 8128 11681 8192
rect 11365 8127 11681 8128
rect 18311 8192 18627 8193
rect 18311 8128 18317 8192
rect 18381 8128 18397 8192
rect 18461 8128 18477 8192
rect 18541 8128 18557 8192
rect 18621 8128 18627 8192
rect 18311 8127 18627 8128
rect 25257 8192 25573 8193
rect 25257 8128 25263 8192
rect 25327 8128 25343 8192
rect 25407 8128 25423 8192
rect 25487 8128 25503 8192
rect 25567 8128 25573 8192
rect 25257 8127 25573 8128
rect 0 7926 1594 7986
rect 28349 7986 28415 7989
rect 29200 7986 30000 8016
rect 28349 7984 30000 7986
rect 28349 7928 28354 7984
rect 28410 7928 30000 7984
rect 28349 7926 30000 7928
rect 0 7896 800 7926
rect 28349 7923 28415 7926
rect 29200 7896 30000 7926
rect 0 7714 800 7744
rect 1761 7714 1827 7717
rect 0 7712 1827 7714
rect 0 7656 1766 7712
rect 1822 7656 1827 7712
rect 0 7654 1827 7656
rect 0 7624 800 7654
rect 1761 7651 1827 7654
rect 2773 7714 2839 7717
rect 3325 7714 3391 7717
rect 2773 7712 3391 7714
rect 2773 7656 2778 7712
rect 2834 7656 3330 7712
rect 3386 7656 3391 7712
rect 2773 7654 3391 7656
rect 2773 7651 2839 7654
rect 3325 7651 3391 7654
rect 7892 7648 8208 7649
rect 7892 7584 7898 7648
rect 7962 7584 7978 7648
rect 8042 7584 8058 7648
rect 8122 7584 8138 7648
rect 8202 7584 8208 7648
rect 7892 7583 8208 7584
rect 14838 7648 15154 7649
rect 14838 7584 14844 7648
rect 14908 7584 14924 7648
rect 14988 7584 15004 7648
rect 15068 7584 15084 7648
rect 15148 7584 15154 7648
rect 14838 7583 15154 7584
rect 21784 7648 22100 7649
rect 21784 7584 21790 7648
rect 21854 7584 21870 7648
rect 21934 7584 21950 7648
rect 22014 7584 22030 7648
rect 22094 7584 22100 7648
rect 21784 7583 22100 7584
rect 28730 7648 29046 7649
rect 28730 7584 28736 7648
rect 28800 7584 28816 7648
rect 28880 7584 28896 7648
rect 28960 7584 28976 7648
rect 29040 7584 29046 7648
rect 28730 7583 29046 7584
rect 0 7442 800 7472
rect 2773 7442 2839 7445
rect 0 7440 2839 7442
rect 0 7384 2778 7440
rect 2834 7384 2839 7440
rect 0 7382 2839 7384
rect 0 7352 800 7382
rect 2773 7379 2839 7382
rect 9765 7442 9831 7445
rect 13169 7442 13235 7445
rect 9765 7440 13235 7442
rect 9765 7384 9770 7440
rect 9826 7384 13174 7440
rect 13230 7384 13235 7440
rect 9765 7382 13235 7384
rect 9765 7379 9831 7382
rect 13169 7379 13235 7382
rect 2497 7306 2563 7309
rect 13261 7306 13327 7309
rect 2497 7304 13327 7306
rect 2497 7248 2502 7304
rect 2558 7248 13266 7304
rect 13322 7248 13327 7304
rect 2497 7246 13327 7248
rect 2497 7243 2563 7246
rect 13261 7243 13327 7246
rect 0 7170 800 7200
rect 933 7170 999 7173
rect 0 7168 999 7170
rect 0 7112 938 7168
rect 994 7112 999 7168
rect 0 7110 999 7112
rect 0 7080 800 7110
rect 933 7107 999 7110
rect 1301 7170 1367 7173
rect 3049 7170 3115 7173
rect 1301 7168 3115 7170
rect 1301 7112 1306 7168
rect 1362 7112 3054 7168
rect 3110 7112 3115 7168
rect 1301 7110 3115 7112
rect 1301 7107 1367 7110
rect 3049 7107 3115 7110
rect 7005 7170 7071 7173
rect 7833 7170 7899 7173
rect 7005 7168 7899 7170
rect 7005 7112 7010 7168
rect 7066 7112 7838 7168
rect 7894 7112 7899 7168
rect 7005 7110 7899 7112
rect 7005 7107 7071 7110
rect 7833 7107 7899 7110
rect 28349 7170 28415 7173
rect 29200 7170 30000 7200
rect 28349 7168 30000 7170
rect 28349 7112 28354 7168
rect 28410 7112 30000 7168
rect 28349 7110 30000 7112
rect 28349 7107 28415 7110
rect 4419 7104 4735 7105
rect 4419 7040 4425 7104
rect 4489 7040 4505 7104
rect 4569 7040 4585 7104
rect 4649 7040 4665 7104
rect 4729 7040 4735 7104
rect 4419 7039 4735 7040
rect 11365 7104 11681 7105
rect 11365 7040 11371 7104
rect 11435 7040 11451 7104
rect 11515 7040 11531 7104
rect 11595 7040 11611 7104
rect 11675 7040 11681 7104
rect 11365 7039 11681 7040
rect 18311 7104 18627 7105
rect 18311 7040 18317 7104
rect 18381 7040 18397 7104
rect 18461 7040 18477 7104
rect 18541 7040 18557 7104
rect 18621 7040 18627 7104
rect 18311 7039 18627 7040
rect 25257 7104 25573 7105
rect 25257 7040 25263 7104
rect 25327 7040 25343 7104
rect 25407 7040 25423 7104
rect 25487 7040 25503 7104
rect 25567 7040 25573 7104
rect 29200 7080 30000 7110
rect 25257 7039 25573 7040
rect 0 6898 800 6928
rect 1485 6898 1551 6901
rect 0 6896 1551 6898
rect 0 6840 1490 6896
rect 1546 6840 1551 6896
rect 0 6838 1551 6840
rect 0 6808 800 6838
rect 1485 6835 1551 6838
rect 1761 6898 1827 6901
rect 6913 6898 6979 6901
rect 1761 6896 6979 6898
rect 1761 6840 1766 6896
rect 1822 6840 6918 6896
rect 6974 6840 6979 6896
rect 1761 6838 6979 6840
rect 1761 6835 1827 6838
rect 6913 6835 6979 6838
rect 8661 6898 8727 6901
rect 10777 6898 10843 6901
rect 8661 6896 10843 6898
rect 8661 6840 8666 6896
rect 8722 6840 10782 6896
rect 10838 6840 10843 6896
rect 8661 6838 10843 6840
rect 8661 6835 8727 6838
rect 10777 6835 10843 6838
rect 6269 6762 6335 6765
rect 8109 6762 8175 6765
rect 6269 6760 8175 6762
rect 6269 6704 6274 6760
rect 6330 6704 8114 6760
rect 8170 6704 8175 6760
rect 6269 6702 8175 6704
rect 6269 6699 6335 6702
rect 8109 6699 8175 6702
rect 0 6626 800 6656
rect 2037 6626 2103 6629
rect 0 6624 2103 6626
rect 0 6568 2042 6624
rect 2098 6568 2103 6624
rect 0 6566 2103 6568
rect 0 6536 800 6566
rect 2037 6563 2103 6566
rect 7892 6560 8208 6561
rect 7892 6496 7898 6560
rect 7962 6496 7978 6560
rect 8042 6496 8058 6560
rect 8122 6496 8138 6560
rect 8202 6496 8208 6560
rect 7892 6495 8208 6496
rect 14838 6560 15154 6561
rect 14838 6496 14844 6560
rect 14908 6496 14924 6560
rect 14988 6496 15004 6560
rect 15068 6496 15084 6560
rect 15148 6496 15154 6560
rect 14838 6495 15154 6496
rect 21784 6560 22100 6561
rect 21784 6496 21790 6560
rect 21854 6496 21870 6560
rect 21934 6496 21950 6560
rect 22014 6496 22030 6560
rect 22094 6496 22100 6560
rect 21784 6495 22100 6496
rect 28730 6560 29046 6561
rect 28730 6496 28736 6560
rect 28800 6496 28816 6560
rect 28880 6496 28896 6560
rect 28960 6496 28976 6560
rect 29040 6496 29046 6560
rect 28730 6495 29046 6496
rect 0 6354 800 6384
rect 1301 6354 1367 6357
rect 0 6352 1367 6354
rect 0 6296 1306 6352
rect 1362 6296 1367 6352
rect 0 6294 1367 6296
rect 0 6264 800 6294
rect 1301 6291 1367 6294
rect 28349 6354 28415 6357
rect 29200 6354 30000 6384
rect 28349 6352 30000 6354
rect 28349 6296 28354 6352
rect 28410 6296 30000 6352
rect 28349 6294 30000 6296
rect 28349 6291 28415 6294
rect 29200 6264 30000 6294
rect 5390 6156 5396 6220
rect 5460 6218 5466 6220
rect 24117 6218 24183 6221
rect 5460 6216 24183 6218
rect 5460 6160 24122 6216
rect 24178 6160 24183 6216
rect 5460 6158 24183 6160
rect 5460 6156 5466 6158
rect 24117 6155 24183 6158
rect 4419 6016 4735 6017
rect 4419 5952 4425 6016
rect 4489 5952 4505 6016
rect 4569 5952 4585 6016
rect 4649 5952 4665 6016
rect 4729 5952 4735 6016
rect 4419 5951 4735 5952
rect 11365 6016 11681 6017
rect 11365 5952 11371 6016
rect 11435 5952 11451 6016
rect 11515 5952 11531 6016
rect 11595 5952 11611 6016
rect 11675 5952 11681 6016
rect 11365 5951 11681 5952
rect 18311 6016 18627 6017
rect 18311 5952 18317 6016
rect 18381 5952 18397 6016
rect 18461 5952 18477 6016
rect 18541 5952 18557 6016
rect 18621 5952 18627 6016
rect 18311 5951 18627 5952
rect 25257 6016 25573 6017
rect 25257 5952 25263 6016
rect 25327 5952 25343 6016
rect 25407 5952 25423 6016
rect 25487 5952 25503 6016
rect 25567 5952 25573 6016
rect 25257 5951 25573 5952
rect 28809 5810 28875 5813
rect 28809 5808 29378 5810
rect 28809 5752 28814 5808
rect 28870 5752 29378 5808
rect 28809 5750 29378 5752
rect 28809 5747 28875 5750
rect 29318 5568 29378 5750
rect 1945 5538 2011 5541
rect 2957 5538 3023 5541
rect 1945 5536 3023 5538
rect 1945 5480 1950 5536
rect 2006 5480 2962 5536
rect 3018 5480 3023 5536
rect 1945 5478 3023 5480
rect 1945 5475 2011 5478
rect 2957 5475 3023 5478
rect 7892 5472 8208 5473
rect 7892 5408 7898 5472
rect 7962 5408 7978 5472
rect 8042 5408 8058 5472
rect 8122 5408 8138 5472
rect 8202 5408 8208 5472
rect 7892 5407 8208 5408
rect 14838 5472 15154 5473
rect 14838 5408 14844 5472
rect 14908 5408 14924 5472
rect 14988 5408 15004 5472
rect 15068 5408 15084 5472
rect 15148 5408 15154 5472
rect 14838 5407 15154 5408
rect 21784 5472 22100 5473
rect 21784 5408 21790 5472
rect 21854 5408 21870 5472
rect 21934 5408 21950 5472
rect 22014 5408 22030 5472
rect 22094 5408 22100 5472
rect 21784 5407 22100 5408
rect 28730 5472 29046 5473
rect 28730 5408 28736 5472
rect 28800 5408 28816 5472
rect 28880 5408 28896 5472
rect 28960 5408 28976 5472
rect 29040 5408 29046 5472
rect 29200 5448 30000 5568
rect 28730 5407 29046 5408
rect 2405 5266 2471 5269
rect 6085 5266 6151 5269
rect 8109 5266 8175 5269
rect 2405 5264 2514 5266
rect 2405 5208 2410 5264
rect 2466 5208 2514 5264
rect 2405 5203 2514 5208
rect 6085 5264 8175 5266
rect 6085 5208 6090 5264
rect 6146 5208 8114 5264
rect 8170 5208 8175 5264
rect 6085 5206 8175 5208
rect 6085 5203 6151 5206
rect 8109 5203 8175 5206
rect 2454 5130 2514 5203
rect 6545 5130 6611 5133
rect 2454 5128 6611 5130
rect 2454 5072 6550 5128
rect 6606 5072 6611 5128
rect 2454 5070 6611 5072
rect 6545 5067 6611 5070
rect 7373 4994 7439 4997
rect 8201 4994 8267 4997
rect 7373 4992 8267 4994
rect 7373 4936 7378 4992
rect 7434 4936 8206 4992
rect 8262 4936 8267 4992
rect 7373 4934 8267 4936
rect 7373 4931 7439 4934
rect 8201 4931 8267 4934
rect 4419 4928 4735 4929
rect 4419 4864 4425 4928
rect 4489 4864 4505 4928
rect 4569 4864 4585 4928
rect 4649 4864 4665 4928
rect 4729 4864 4735 4928
rect 4419 4863 4735 4864
rect 11365 4928 11681 4929
rect 11365 4864 11371 4928
rect 11435 4864 11451 4928
rect 11515 4864 11531 4928
rect 11595 4864 11611 4928
rect 11675 4864 11681 4928
rect 11365 4863 11681 4864
rect 18311 4928 18627 4929
rect 18311 4864 18317 4928
rect 18381 4864 18397 4928
rect 18461 4864 18477 4928
rect 18541 4864 18557 4928
rect 18621 4864 18627 4928
rect 18311 4863 18627 4864
rect 25257 4928 25573 4929
rect 25257 4864 25263 4928
rect 25327 4864 25343 4928
rect 25407 4864 25423 4928
rect 25487 4864 25503 4928
rect 25567 4864 25573 4928
rect 25257 4863 25573 4864
rect 4061 4722 4127 4725
rect 8109 4722 8175 4725
rect 4061 4720 8175 4722
rect 4061 4664 4066 4720
rect 4122 4664 8114 4720
rect 8170 4664 8175 4720
rect 4061 4662 8175 4664
rect 4061 4659 4127 4662
rect 8109 4659 8175 4662
rect 20897 4722 20963 4725
rect 25865 4722 25931 4725
rect 20897 4720 25931 4722
rect 20897 4664 20902 4720
rect 20958 4664 25870 4720
rect 25926 4664 25931 4720
rect 20897 4662 25931 4664
rect 20897 4659 20963 4662
rect 25865 4659 25931 4662
rect 28717 4722 28783 4725
rect 29200 4722 30000 4752
rect 28717 4720 30000 4722
rect 28717 4664 28722 4720
rect 28778 4664 30000 4720
rect 28717 4662 30000 4664
rect 28717 4659 28783 4662
rect 29200 4632 30000 4662
rect 7892 4384 8208 4385
rect 7892 4320 7898 4384
rect 7962 4320 7978 4384
rect 8042 4320 8058 4384
rect 8122 4320 8138 4384
rect 8202 4320 8208 4384
rect 7892 4319 8208 4320
rect 14838 4384 15154 4385
rect 14838 4320 14844 4384
rect 14908 4320 14924 4384
rect 14988 4320 15004 4384
rect 15068 4320 15084 4384
rect 15148 4320 15154 4384
rect 14838 4319 15154 4320
rect 21784 4384 22100 4385
rect 21784 4320 21790 4384
rect 21854 4320 21870 4384
rect 21934 4320 21950 4384
rect 22014 4320 22030 4384
rect 22094 4320 22100 4384
rect 21784 4319 22100 4320
rect 28730 4384 29046 4385
rect 28730 4320 28736 4384
rect 28800 4320 28816 4384
rect 28880 4320 28896 4384
rect 28960 4320 28976 4384
rect 29040 4320 29046 4384
rect 28730 4319 29046 4320
rect 8753 4314 8819 4317
rect 9857 4314 9923 4317
rect 8753 4312 9923 4314
rect 8753 4256 8758 4312
rect 8814 4256 9862 4312
rect 9918 4256 9923 4312
rect 8753 4254 9923 4256
rect 8753 4251 8819 4254
rect 9857 4251 9923 4254
rect 9305 4178 9371 4181
rect 11329 4178 11395 4181
rect 9305 4176 11395 4178
rect 9305 4120 9310 4176
rect 9366 4120 11334 4176
rect 11390 4120 11395 4176
rect 9305 4118 11395 4120
rect 9305 4115 9371 4118
rect 11329 4115 11395 4118
rect 4102 3980 4108 4044
rect 4172 4042 4178 4044
rect 4797 4042 4863 4045
rect 4172 4040 4863 4042
rect 4172 3984 4802 4040
rect 4858 3984 4863 4040
rect 4172 3982 4863 3984
rect 4172 3980 4178 3982
rect 4797 3979 4863 3982
rect 8569 4042 8635 4045
rect 10593 4042 10659 4045
rect 8569 4040 10659 4042
rect 8569 3984 8574 4040
rect 8630 3984 10598 4040
rect 10654 3984 10659 4040
rect 8569 3982 10659 3984
rect 8569 3979 8635 3982
rect 10593 3979 10659 3982
rect 26877 3906 26943 3909
rect 29200 3906 30000 3936
rect 26877 3904 30000 3906
rect 26877 3848 26882 3904
rect 26938 3848 30000 3904
rect 26877 3846 30000 3848
rect 26877 3843 26943 3846
rect 4419 3840 4735 3841
rect 4419 3776 4425 3840
rect 4489 3776 4505 3840
rect 4569 3776 4585 3840
rect 4649 3776 4665 3840
rect 4729 3776 4735 3840
rect 4419 3775 4735 3776
rect 11365 3840 11681 3841
rect 11365 3776 11371 3840
rect 11435 3776 11451 3840
rect 11515 3776 11531 3840
rect 11595 3776 11611 3840
rect 11675 3776 11681 3840
rect 11365 3775 11681 3776
rect 18311 3840 18627 3841
rect 18311 3776 18317 3840
rect 18381 3776 18397 3840
rect 18461 3776 18477 3840
rect 18541 3776 18557 3840
rect 18621 3776 18627 3840
rect 18311 3775 18627 3776
rect 25257 3840 25573 3841
rect 25257 3776 25263 3840
rect 25327 3776 25343 3840
rect 25407 3776 25423 3840
rect 25487 3776 25503 3840
rect 25567 3776 25573 3840
rect 29200 3816 30000 3846
rect 25257 3775 25573 3776
rect 10133 3770 10199 3773
rect 10777 3770 10843 3773
rect 10133 3768 10843 3770
rect 10133 3712 10138 3768
rect 10194 3712 10782 3768
rect 10838 3712 10843 3768
rect 10133 3710 10843 3712
rect 10133 3707 10199 3710
rect 10777 3707 10843 3710
rect 9581 3634 9647 3637
rect 12249 3634 12315 3637
rect 9581 3632 12315 3634
rect 9581 3576 9586 3632
rect 9642 3576 12254 3632
rect 12310 3576 12315 3632
rect 9581 3574 12315 3576
rect 9581 3571 9647 3574
rect 12249 3571 12315 3574
rect 2037 3498 2103 3501
rect 5073 3498 5139 3501
rect 15193 3498 15259 3501
rect 2037 3496 15259 3498
rect 2037 3440 2042 3496
rect 2098 3440 5078 3496
rect 5134 3440 15198 3496
rect 15254 3440 15259 3496
rect 2037 3438 15259 3440
rect 2037 3435 2103 3438
rect 5073 3435 5139 3438
rect 15193 3435 15259 3438
rect 2865 3362 2931 3365
rect 4521 3362 4587 3365
rect 2865 3360 4587 3362
rect 2865 3304 2870 3360
rect 2926 3304 4526 3360
rect 4582 3304 4587 3360
rect 2865 3302 4587 3304
rect 2865 3299 2931 3302
rect 4521 3299 4587 3302
rect 7892 3296 8208 3297
rect 7892 3232 7898 3296
rect 7962 3232 7978 3296
rect 8042 3232 8058 3296
rect 8122 3232 8138 3296
rect 8202 3232 8208 3296
rect 7892 3231 8208 3232
rect 14838 3296 15154 3297
rect 14838 3232 14844 3296
rect 14908 3232 14924 3296
rect 14988 3232 15004 3296
rect 15068 3232 15084 3296
rect 15148 3232 15154 3296
rect 14838 3231 15154 3232
rect 21784 3296 22100 3297
rect 21784 3232 21790 3296
rect 21854 3232 21870 3296
rect 21934 3232 21950 3296
rect 22014 3232 22030 3296
rect 22094 3232 22100 3296
rect 21784 3231 22100 3232
rect 28730 3296 29046 3297
rect 28730 3232 28736 3296
rect 28800 3232 28816 3296
rect 28880 3232 28896 3296
rect 28960 3232 28976 3296
rect 29040 3232 29046 3296
rect 28730 3231 29046 3232
rect 24669 3090 24735 3093
rect 29200 3090 30000 3120
rect 24669 3088 30000 3090
rect 24669 3032 24674 3088
rect 24730 3032 30000 3088
rect 24669 3030 30000 3032
rect 24669 3027 24735 3030
rect 29200 3000 30000 3030
rect 6729 2954 6795 2957
rect 21817 2954 21883 2957
rect 6729 2952 21883 2954
rect 6729 2896 6734 2952
rect 6790 2896 21822 2952
rect 21878 2896 21883 2952
rect 6729 2894 21883 2896
rect 6729 2891 6795 2894
rect 21817 2891 21883 2894
rect 23381 2954 23447 2957
rect 28625 2954 28691 2957
rect 23381 2952 28691 2954
rect 23381 2896 23386 2952
rect 23442 2896 28630 2952
rect 28686 2896 28691 2952
rect 23381 2894 28691 2896
rect 23381 2891 23447 2894
rect 28625 2891 28691 2894
rect 4419 2752 4735 2753
rect 4419 2688 4425 2752
rect 4489 2688 4505 2752
rect 4569 2688 4585 2752
rect 4649 2688 4665 2752
rect 4729 2688 4735 2752
rect 4419 2687 4735 2688
rect 11365 2752 11681 2753
rect 11365 2688 11371 2752
rect 11435 2688 11451 2752
rect 11515 2688 11531 2752
rect 11595 2688 11611 2752
rect 11675 2688 11681 2752
rect 11365 2687 11681 2688
rect 18311 2752 18627 2753
rect 18311 2688 18317 2752
rect 18381 2688 18397 2752
rect 18461 2688 18477 2752
rect 18541 2688 18557 2752
rect 18621 2688 18627 2752
rect 18311 2687 18627 2688
rect 25257 2752 25573 2753
rect 25257 2688 25263 2752
rect 25327 2688 25343 2752
rect 25407 2688 25423 2752
rect 25487 2688 25503 2752
rect 25567 2688 25573 2752
rect 25257 2687 25573 2688
rect 25589 2410 25655 2413
rect 25589 2408 29194 2410
rect 25589 2352 25594 2408
rect 25650 2352 29194 2408
rect 25589 2350 29194 2352
rect 25589 2347 25655 2350
rect 29134 2308 29194 2350
rect 29134 2304 29378 2308
rect 29134 2248 30000 2304
rect 7892 2208 8208 2209
rect 7892 2144 7898 2208
rect 7962 2144 7978 2208
rect 8042 2144 8058 2208
rect 8122 2144 8138 2208
rect 8202 2144 8208 2208
rect 7892 2143 8208 2144
rect 14838 2208 15154 2209
rect 14838 2144 14844 2208
rect 14908 2144 14924 2208
rect 14988 2144 15004 2208
rect 15068 2144 15084 2208
rect 15148 2144 15154 2208
rect 14838 2143 15154 2144
rect 21784 2208 22100 2209
rect 21784 2144 21790 2208
rect 21854 2144 21870 2208
rect 21934 2144 21950 2208
rect 22014 2144 22030 2208
rect 22094 2144 22100 2208
rect 21784 2143 22100 2144
rect 28730 2208 29046 2209
rect 28730 2144 28736 2208
rect 28800 2144 28816 2208
rect 28880 2144 28896 2208
rect 28960 2144 28976 2208
rect 29040 2144 29046 2208
rect 29200 2184 30000 2248
rect 28730 2143 29046 2144
<< via3 >>
rect 4425 27772 4489 27776
rect 4425 27716 4429 27772
rect 4429 27716 4485 27772
rect 4485 27716 4489 27772
rect 4425 27712 4489 27716
rect 4505 27772 4569 27776
rect 4505 27716 4509 27772
rect 4509 27716 4565 27772
rect 4565 27716 4569 27772
rect 4505 27712 4569 27716
rect 4585 27772 4649 27776
rect 4585 27716 4589 27772
rect 4589 27716 4645 27772
rect 4645 27716 4649 27772
rect 4585 27712 4649 27716
rect 4665 27772 4729 27776
rect 4665 27716 4669 27772
rect 4669 27716 4725 27772
rect 4725 27716 4729 27772
rect 4665 27712 4729 27716
rect 11371 27772 11435 27776
rect 11371 27716 11375 27772
rect 11375 27716 11431 27772
rect 11431 27716 11435 27772
rect 11371 27712 11435 27716
rect 11451 27772 11515 27776
rect 11451 27716 11455 27772
rect 11455 27716 11511 27772
rect 11511 27716 11515 27772
rect 11451 27712 11515 27716
rect 11531 27772 11595 27776
rect 11531 27716 11535 27772
rect 11535 27716 11591 27772
rect 11591 27716 11595 27772
rect 11531 27712 11595 27716
rect 11611 27772 11675 27776
rect 11611 27716 11615 27772
rect 11615 27716 11671 27772
rect 11671 27716 11675 27772
rect 11611 27712 11675 27716
rect 18317 27772 18381 27776
rect 18317 27716 18321 27772
rect 18321 27716 18377 27772
rect 18377 27716 18381 27772
rect 18317 27712 18381 27716
rect 18397 27772 18461 27776
rect 18397 27716 18401 27772
rect 18401 27716 18457 27772
rect 18457 27716 18461 27772
rect 18397 27712 18461 27716
rect 18477 27772 18541 27776
rect 18477 27716 18481 27772
rect 18481 27716 18537 27772
rect 18537 27716 18541 27772
rect 18477 27712 18541 27716
rect 18557 27772 18621 27776
rect 18557 27716 18561 27772
rect 18561 27716 18617 27772
rect 18617 27716 18621 27772
rect 18557 27712 18621 27716
rect 25263 27772 25327 27776
rect 25263 27716 25267 27772
rect 25267 27716 25323 27772
rect 25323 27716 25327 27772
rect 25263 27712 25327 27716
rect 25343 27772 25407 27776
rect 25343 27716 25347 27772
rect 25347 27716 25403 27772
rect 25403 27716 25407 27772
rect 25343 27712 25407 27716
rect 25423 27772 25487 27776
rect 25423 27716 25427 27772
rect 25427 27716 25483 27772
rect 25483 27716 25487 27772
rect 25423 27712 25487 27716
rect 25503 27772 25567 27776
rect 25503 27716 25507 27772
rect 25507 27716 25563 27772
rect 25563 27716 25567 27772
rect 25503 27712 25567 27716
rect 7898 27228 7962 27232
rect 7898 27172 7902 27228
rect 7902 27172 7958 27228
rect 7958 27172 7962 27228
rect 7898 27168 7962 27172
rect 7978 27228 8042 27232
rect 7978 27172 7982 27228
rect 7982 27172 8038 27228
rect 8038 27172 8042 27228
rect 7978 27168 8042 27172
rect 8058 27228 8122 27232
rect 8058 27172 8062 27228
rect 8062 27172 8118 27228
rect 8118 27172 8122 27228
rect 8058 27168 8122 27172
rect 8138 27228 8202 27232
rect 8138 27172 8142 27228
rect 8142 27172 8198 27228
rect 8198 27172 8202 27228
rect 8138 27168 8202 27172
rect 14844 27228 14908 27232
rect 14844 27172 14848 27228
rect 14848 27172 14904 27228
rect 14904 27172 14908 27228
rect 14844 27168 14908 27172
rect 14924 27228 14988 27232
rect 14924 27172 14928 27228
rect 14928 27172 14984 27228
rect 14984 27172 14988 27228
rect 14924 27168 14988 27172
rect 15004 27228 15068 27232
rect 15004 27172 15008 27228
rect 15008 27172 15064 27228
rect 15064 27172 15068 27228
rect 15004 27168 15068 27172
rect 15084 27228 15148 27232
rect 15084 27172 15088 27228
rect 15088 27172 15144 27228
rect 15144 27172 15148 27228
rect 15084 27168 15148 27172
rect 21790 27228 21854 27232
rect 21790 27172 21794 27228
rect 21794 27172 21850 27228
rect 21850 27172 21854 27228
rect 21790 27168 21854 27172
rect 21870 27228 21934 27232
rect 21870 27172 21874 27228
rect 21874 27172 21930 27228
rect 21930 27172 21934 27228
rect 21870 27168 21934 27172
rect 21950 27228 22014 27232
rect 21950 27172 21954 27228
rect 21954 27172 22010 27228
rect 22010 27172 22014 27228
rect 21950 27168 22014 27172
rect 22030 27228 22094 27232
rect 22030 27172 22034 27228
rect 22034 27172 22090 27228
rect 22090 27172 22094 27228
rect 22030 27168 22094 27172
rect 28736 27228 28800 27232
rect 28736 27172 28740 27228
rect 28740 27172 28796 27228
rect 28796 27172 28800 27228
rect 28736 27168 28800 27172
rect 28816 27228 28880 27232
rect 28816 27172 28820 27228
rect 28820 27172 28876 27228
rect 28876 27172 28880 27228
rect 28816 27168 28880 27172
rect 28896 27228 28960 27232
rect 28896 27172 28900 27228
rect 28900 27172 28956 27228
rect 28956 27172 28960 27228
rect 28896 27168 28960 27172
rect 28976 27228 29040 27232
rect 28976 27172 28980 27228
rect 28980 27172 29036 27228
rect 29036 27172 29040 27228
rect 28976 27168 29040 27172
rect 4425 26684 4489 26688
rect 4425 26628 4429 26684
rect 4429 26628 4485 26684
rect 4485 26628 4489 26684
rect 4425 26624 4489 26628
rect 4505 26684 4569 26688
rect 4505 26628 4509 26684
rect 4509 26628 4565 26684
rect 4565 26628 4569 26684
rect 4505 26624 4569 26628
rect 4585 26684 4649 26688
rect 4585 26628 4589 26684
rect 4589 26628 4645 26684
rect 4645 26628 4649 26684
rect 4585 26624 4649 26628
rect 4665 26684 4729 26688
rect 4665 26628 4669 26684
rect 4669 26628 4725 26684
rect 4725 26628 4729 26684
rect 4665 26624 4729 26628
rect 11371 26684 11435 26688
rect 11371 26628 11375 26684
rect 11375 26628 11431 26684
rect 11431 26628 11435 26684
rect 11371 26624 11435 26628
rect 11451 26684 11515 26688
rect 11451 26628 11455 26684
rect 11455 26628 11511 26684
rect 11511 26628 11515 26684
rect 11451 26624 11515 26628
rect 11531 26684 11595 26688
rect 11531 26628 11535 26684
rect 11535 26628 11591 26684
rect 11591 26628 11595 26684
rect 11531 26624 11595 26628
rect 11611 26684 11675 26688
rect 11611 26628 11615 26684
rect 11615 26628 11671 26684
rect 11671 26628 11675 26684
rect 11611 26624 11675 26628
rect 18317 26684 18381 26688
rect 18317 26628 18321 26684
rect 18321 26628 18377 26684
rect 18377 26628 18381 26684
rect 18317 26624 18381 26628
rect 18397 26684 18461 26688
rect 18397 26628 18401 26684
rect 18401 26628 18457 26684
rect 18457 26628 18461 26684
rect 18397 26624 18461 26628
rect 18477 26684 18541 26688
rect 18477 26628 18481 26684
rect 18481 26628 18537 26684
rect 18537 26628 18541 26684
rect 18477 26624 18541 26628
rect 18557 26684 18621 26688
rect 18557 26628 18561 26684
rect 18561 26628 18617 26684
rect 18617 26628 18621 26684
rect 18557 26624 18621 26628
rect 25263 26684 25327 26688
rect 25263 26628 25267 26684
rect 25267 26628 25323 26684
rect 25323 26628 25327 26684
rect 25263 26624 25327 26628
rect 25343 26684 25407 26688
rect 25343 26628 25347 26684
rect 25347 26628 25403 26684
rect 25403 26628 25407 26684
rect 25343 26624 25407 26628
rect 25423 26684 25487 26688
rect 25423 26628 25427 26684
rect 25427 26628 25483 26684
rect 25483 26628 25487 26684
rect 25423 26624 25487 26628
rect 25503 26684 25567 26688
rect 25503 26628 25507 26684
rect 25507 26628 25563 26684
rect 25563 26628 25567 26684
rect 25503 26624 25567 26628
rect 7898 26140 7962 26144
rect 7898 26084 7902 26140
rect 7902 26084 7958 26140
rect 7958 26084 7962 26140
rect 7898 26080 7962 26084
rect 7978 26140 8042 26144
rect 7978 26084 7982 26140
rect 7982 26084 8038 26140
rect 8038 26084 8042 26140
rect 7978 26080 8042 26084
rect 8058 26140 8122 26144
rect 8058 26084 8062 26140
rect 8062 26084 8118 26140
rect 8118 26084 8122 26140
rect 8058 26080 8122 26084
rect 8138 26140 8202 26144
rect 8138 26084 8142 26140
rect 8142 26084 8198 26140
rect 8198 26084 8202 26140
rect 8138 26080 8202 26084
rect 14844 26140 14908 26144
rect 14844 26084 14848 26140
rect 14848 26084 14904 26140
rect 14904 26084 14908 26140
rect 14844 26080 14908 26084
rect 14924 26140 14988 26144
rect 14924 26084 14928 26140
rect 14928 26084 14984 26140
rect 14984 26084 14988 26140
rect 14924 26080 14988 26084
rect 15004 26140 15068 26144
rect 15004 26084 15008 26140
rect 15008 26084 15064 26140
rect 15064 26084 15068 26140
rect 15004 26080 15068 26084
rect 15084 26140 15148 26144
rect 15084 26084 15088 26140
rect 15088 26084 15144 26140
rect 15144 26084 15148 26140
rect 15084 26080 15148 26084
rect 21790 26140 21854 26144
rect 21790 26084 21794 26140
rect 21794 26084 21850 26140
rect 21850 26084 21854 26140
rect 21790 26080 21854 26084
rect 21870 26140 21934 26144
rect 21870 26084 21874 26140
rect 21874 26084 21930 26140
rect 21930 26084 21934 26140
rect 21870 26080 21934 26084
rect 21950 26140 22014 26144
rect 21950 26084 21954 26140
rect 21954 26084 22010 26140
rect 22010 26084 22014 26140
rect 21950 26080 22014 26084
rect 22030 26140 22094 26144
rect 22030 26084 22034 26140
rect 22034 26084 22090 26140
rect 22090 26084 22094 26140
rect 22030 26080 22094 26084
rect 28736 26140 28800 26144
rect 28736 26084 28740 26140
rect 28740 26084 28796 26140
rect 28796 26084 28800 26140
rect 28736 26080 28800 26084
rect 28816 26140 28880 26144
rect 28816 26084 28820 26140
rect 28820 26084 28876 26140
rect 28876 26084 28880 26140
rect 28816 26080 28880 26084
rect 28896 26140 28960 26144
rect 28896 26084 28900 26140
rect 28900 26084 28956 26140
rect 28956 26084 28960 26140
rect 28896 26080 28960 26084
rect 28976 26140 29040 26144
rect 28976 26084 28980 26140
rect 28980 26084 29036 26140
rect 29036 26084 29040 26140
rect 28976 26080 29040 26084
rect 4425 25596 4489 25600
rect 4425 25540 4429 25596
rect 4429 25540 4485 25596
rect 4485 25540 4489 25596
rect 4425 25536 4489 25540
rect 4505 25596 4569 25600
rect 4505 25540 4509 25596
rect 4509 25540 4565 25596
rect 4565 25540 4569 25596
rect 4505 25536 4569 25540
rect 4585 25596 4649 25600
rect 4585 25540 4589 25596
rect 4589 25540 4645 25596
rect 4645 25540 4649 25596
rect 4585 25536 4649 25540
rect 4665 25596 4729 25600
rect 4665 25540 4669 25596
rect 4669 25540 4725 25596
rect 4725 25540 4729 25596
rect 4665 25536 4729 25540
rect 11371 25596 11435 25600
rect 11371 25540 11375 25596
rect 11375 25540 11431 25596
rect 11431 25540 11435 25596
rect 11371 25536 11435 25540
rect 11451 25596 11515 25600
rect 11451 25540 11455 25596
rect 11455 25540 11511 25596
rect 11511 25540 11515 25596
rect 11451 25536 11515 25540
rect 11531 25596 11595 25600
rect 11531 25540 11535 25596
rect 11535 25540 11591 25596
rect 11591 25540 11595 25596
rect 11531 25536 11595 25540
rect 11611 25596 11675 25600
rect 11611 25540 11615 25596
rect 11615 25540 11671 25596
rect 11671 25540 11675 25596
rect 11611 25536 11675 25540
rect 18317 25596 18381 25600
rect 18317 25540 18321 25596
rect 18321 25540 18377 25596
rect 18377 25540 18381 25596
rect 18317 25536 18381 25540
rect 18397 25596 18461 25600
rect 18397 25540 18401 25596
rect 18401 25540 18457 25596
rect 18457 25540 18461 25596
rect 18397 25536 18461 25540
rect 18477 25596 18541 25600
rect 18477 25540 18481 25596
rect 18481 25540 18537 25596
rect 18537 25540 18541 25596
rect 18477 25536 18541 25540
rect 18557 25596 18621 25600
rect 18557 25540 18561 25596
rect 18561 25540 18617 25596
rect 18617 25540 18621 25596
rect 18557 25536 18621 25540
rect 25263 25596 25327 25600
rect 25263 25540 25267 25596
rect 25267 25540 25323 25596
rect 25323 25540 25327 25596
rect 25263 25536 25327 25540
rect 25343 25596 25407 25600
rect 25343 25540 25347 25596
rect 25347 25540 25403 25596
rect 25403 25540 25407 25596
rect 25343 25536 25407 25540
rect 25423 25596 25487 25600
rect 25423 25540 25427 25596
rect 25427 25540 25483 25596
rect 25483 25540 25487 25596
rect 25423 25536 25487 25540
rect 25503 25596 25567 25600
rect 25503 25540 25507 25596
rect 25507 25540 25563 25596
rect 25563 25540 25567 25596
rect 25503 25536 25567 25540
rect 7898 25052 7962 25056
rect 7898 24996 7902 25052
rect 7902 24996 7958 25052
rect 7958 24996 7962 25052
rect 7898 24992 7962 24996
rect 7978 25052 8042 25056
rect 7978 24996 7982 25052
rect 7982 24996 8038 25052
rect 8038 24996 8042 25052
rect 7978 24992 8042 24996
rect 8058 25052 8122 25056
rect 8058 24996 8062 25052
rect 8062 24996 8118 25052
rect 8118 24996 8122 25052
rect 8058 24992 8122 24996
rect 8138 25052 8202 25056
rect 8138 24996 8142 25052
rect 8142 24996 8198 25052
rect 8198 24996 8202 25052
rect 8138 24992 8202 24996
rect 14844 25052 14908 25056
rect 14844 24996 14848 25052
rect 14848 24996 14904 25052
rect 14904 24996 14908 25052
rect 14844 24992 14908 24996
rect 14924 25052 14988 25056
rect 14924 24996 14928 25052
rect 14928 24996 14984 25052
rect 14984 24996 14988 25052
rect 14924 24992 14988 24996
rect 15004 25052 15068 25056
rect 15004 24996 15008 25052
rect 15008 24996 15064 25052
rect 15064 24996 15068 25052
rect 15004 24992 15068 24996
rect 15084 25052 15148 25056
rect 15084 24996 15088 25052
rect 15088 24996 15144 25052
rect 15144 24996 15148 25052
rect 15084 24992 15148 24996
rect 21790 25052 21854 25056
rect 21790 24996 21794 25052
rect 21794 24996 21850 25052
rect 21850 24996 21854 25052
rect 21790 24992 21854 24996
rect 21870 25052 21934 25056
rect 21870 24996 21874 25052
rect 21874 24996 21930 25052
rect 21930 24996 21934 25052
rect 21870 24992 21934 24996
rect 21950 25052 22014 25056
rect 21950 24996 21954 25052
rect 21954 24996 22010 25052
rect 22010 24996 22014 25052
rect 21950 24992 22014 24996
rect 22030 25052 22094 25056
rect 22030 24996 22034 25052
rect 22034 24996 22090 25052
rect 22090 24996 22094 25052
rect 22030 24992 22094 24996
rect 28736 25052 28800 25056
rect 28736 24996 28740 25052
rect 28740 24996 28796 25052
rect 28796 24996 28800 25052
rect 28736 24992 28800 24996
rect 28816 25052 28880 25056
rect 28816 24996 28820 25052
rect 28820 24996 28876 25052
rect 28876 24996 28880 25052
rect 28816 24992 28880 24996
rect 28896 25052 28960 25056
rect 28896 24996 28900 25052
rect 28900 24996 28956 25052
rect 28956 24996 28960 25052
rect 28896 24992 28960 24996
rect 28976 25052 29040 25056
rect 28976 24996 28980 25052
rect 28980 24996 29036 25052
rect 29036 24996 29040 25052
rect 28976 24992 29040 24996
rect 4425 24508 4489 24512
rect 4425 24452 4429 24508
rect 4429 24452 4485 24508
rect 4485 24452 4489 24508
rect 4425 24448 4489 24452
rect 4505 24508 4569 24512
rect 4505 24452 4509 24508
rect 4509 24452 4565 24508
rect 4565 24452 4569 24508
rect 4505 24448 4569 24452
rect 4585 24508 4649 24512
rect 4585 24452 4589 24508
rect 4589 24452 4645 24508
rect 4645 24452 4649 24508
rect 4585 24448 4649 24452
rect 4665 24508 4729 24512
rect 4665 24452 4669 24508
rect 4669 24452 4725 24508
rect 4725 24452 4729 24508
rect 4665 24448 4729 24452
rect 11371 24508 11435 24512
rect 11371 24452 11375 24508
rect 11375 24452 11431 24508
rect 11431 24452 11435 24508
rect 11371 24448 11435 24452
rect 11451 24508 11515 24512
rect 11451 24452 11455 24508
rect 11455 24452 11511 24508
rect 11511 24452 11515 24508
rect 11451 24448 11515 24452
rect 11531 24508 11595 24512
rect 11531 24452 11535 24508
rect 11535 24452 11591 24508
rect 11591 24452 11595 24508
rect 11531 24448 11595 24452
rect 11611 24508 11675 24512
rect 11611 24452 11615 24508
rect 11615 24452 11671 24508
rect 11671 24452 11675 24508
rect 11611 24448 11675 24452
rect 18317 24508 18381 24512
rect 18317 24452 18321 24508
rect 18321 24452 18377 24508
rect 18377 24452 18381 24508
rect 18317 24448 18381 24452
rect 18397 24508 18461 24512
rect 18397 24452 18401 24508
rect 18401 24452 18457 24508
rect 18457 24452 18461 24508
rect 18397 24448 18461 24452
rect 18477 24508 18541 24512
rect 18477 24452 18481 24508
rect 18481 24452 18537 24508
rect 18537 24452 18541 24508
rect 18477 24448 18541 24452
rect 18557 24508 18621 24512
rect 18557 24452 18561 24508
rect 18561 24452 18617 24508
rect 18617 24452 18621 24508
rect 18557 24448 18621 24452
rect 25263 24508 25327 24512
rect 25263 24452 25267 24508
rect 25267 24452 25323 24508
rect 25323 24452 25327 24508
rect 25263 24448 25327 24452
rect 25343 24508 25407 24512
rect 25343 24452 25347 24508
rect 25347 24452 25403 24508
rect 25403 24452 25407 24508
rect 25343 24448 25407 24452
rect 25423 24508 25487 24512
rect 25423 24452 25427 24508
rect 25427 24452 25483 24508
rect 25483 24452 25487 24508
rect 25423 24448 25487 24452
rect 25503 24508 25567 24512
rect 25503 24452 25507 24508
rect 25507 24452 25563 24508
rect 25563 24452 25567 24508
rect 25503 24448 25567 24452
rect 7898 23964 7962 23968
rect 7898 23908 7902 23964
rect 7902 23908 7958 23964
rect 7958 23908 7962 23964
rect 7898 23904 7962 23908
rect 7978 23964 8042 23968
rect 7978 23908 7982 23964
rect 7982 23908 8038 23964
rect 8038 23908 8042 23964
rect 7978 23904 8042 23908
rect 8058 23964 8122 23968
rect 8058 23908 8062 23964
rect 8062 23908 8118 23964
rect 8118 23908 8122 23964
rect 8058 23904 8122 23908
rect 8138 23964 8202 23968
rect 8138 23908 8142 23964
rect 8142 23908 8198 23964
rect 8198 23908 8202 23964
rect 8138 23904 8202 23908
rect 14844 23964 14908 23968
rect 14844 23908 14848 23964
rect 14848 23908 14904 23964
rect 14904 23908 14908 23964
rect 14844 23904 14908 23908
rect 14924 23964 14988 23968
rect 14924 23908 14928 23964
rect 14928 23908 14984 23964
rect 14984 23908 14988 23964
rect 14924 23904 14988 23908
rect 15004 23964 15068 23968
rect 15004 23908 15008 23964
rect 15008 23908 15064 23964
rect 15064 23908 15068 23964
rect 15004 23904 15068 23908
rect 15084 23964 15148 23968
rect 15084 23908 15088 23964
rect 15088 23908 15144 23964
rect 15144 23908 15148 23964
rect 15084 23904 15148 23908
rect 21790 23964 21854 23968
rect 21790 23908 21794 23964
rect 21794 23908 21850 23964
rect 21850 23908 21854 23964
rect 21790 23904 21854 23908
rect 21870 23964 21934 23968
rect 21870 23908 21874 23964
rect 21874 23908 21930 23964
rect 21930 23908 21934 23964
rect 21870 23904 21934 23908
rect 21950 23964 22014 23968
rect 21950 23908 21954 23964
rect 21954 23908 22010 23964
rect 22010 23908 22014 23964
rect 21950 23904 22014 23908
rect 22030 23964 22094 23968
rect 22030 23908 22034 23964
rect 22034 23908 22090 23964
rect 22090 23908 22094 23964
rect 22030 23904 22094 23908
rect 28736 23964 28800 23968
rect 28736 23908 28740 23964
rect 28740 23908 28796 23964
rect 28796 23908 28800 23964
rect 28736 23904 28800 23908
rect 28816 23964 28880 23968
rect 28816 23908 28820 23964
rect 28820 23908 28876 23964
rect 28876 23908 28880 23964
rect 28816 23904 28880 23908
rect 28896 23964 28960 23968
rect 28896 23908 28900 23964
rect 28900 23908 28956 23964
rect 28956 23908 28960 23964
rect 28896 23904 28960 23908
rect 28976 23964 29040 23968
rect 28976 23908 28980 23964
rect 28980 23908 29036 23964
rect 29036 23908 29040 23964
rect 28976 23904 29040 23908
rect 4425 23420 4489 23424
rect 4425 23364 4429 23420
rect 4429 23364 4485 23420
rect 4485 23364 4489 23420
rect 4425 23360 4489 23364
rect 4505 23420 4569 23424
rect 4505 23364 4509 23420
rect 4509 23364 4565 23420
rect 4565 23364 4569 23420
rect 4505 23360 4569 23364
rect 4585 23420 4649 23424
rect 4585 23364 4589 23420
rect 4589 23364 4645 23420
rect 4645 23364 4649 23420
rect 4585 23360 4649 23364
rect 4665 23420 4729 23424
rect 4665 23364 4669 23420
rect 4669 23364 4725 23420
rect 4725 23364 4729 23420
rect 4665 23360 4729 23364
rect 11371 23420 11435 23424
rect 11371 23364 11375 23420
rect 11375 23364 11431 23420
rect 11431 23364 11435 23420
rect 11371 23360 11435 23364
rect 11451 23420 11515 23424
rect 11451 23364 11455 23420
rect 11455 23364 11511 23420
rect 11511 23364 11515 23420
rect 11451 23360 11515 23364
rect 11531 23420 11595 23424
rect 11531 23364 11535 23420
rect 11535 23364 11591 23420
rect 11591 23364 11595 23420
rect 11531 23360 11595 23364
rect 11611 23420 11675 23424
rect 11611 23364 11615 23420
rect 11615 23364 11671 23420
rect 11671 23364 11675 23420
rect 11611 23360 11675 23364
rect 18317 23420 18381 23424
rect 18317 23364 18321 23420
rect 18321 23364 18377 23420
rect 18377 23364 18381 23420
rect 18317 23360 18381 23364
rect 18397 23420 18461 23424
rect 18397 23364 18401 23420
rect 18401 23364 18457 23420
rect 18457 23364 18461 23420
rect 18397 23360 18461 23364
rect 18477 23420 18541 23424
rect 18477 23364 18481 23420
rect 18481 23364 18537 23420
rect 18537 23364 18541 23420
rect 18477 23360 18541 23364
rect 18557 23420 18621 23424
rect 18557 23364 18561 23420
rect 18561 23364 18617 23420
rect 18617 23364 18621 23420
rect 18557 23360 18621 23364
rect 25263 23420 25327 23424
rect 25263 23364 25267 23420
rect 25267 23364 25323 23420
rect 25323 23364 25327 23420
rect 25263 23360 25327 23364
rect 25343 23420 25407 23424
rect 25343 23364 25347 23420
rect 25347 23364 25403 23420
rect 25403 23364 25407 23420
rect 25343 23360 25407 23364
rect 25423 23420 25487 23424
rect 25423 23364 25427 23420
rect 25427 23364 25483 23420
rect 25483 23364 25487 23420
rect 25423 23360 25487 23364
rect 25503 23420 25567 23424
rect 25503 23364 25507 23420
rect 25507 23364 25563 23420
rect 25563 23364 25567 23420
rect 25503 23360 25567 23364
rect 7898 22876 7962 22880
rect 7898 22820 7902 22876
rect 7902 22820 7958 22876
rect 7958 22820 7962 22876
rect 7898 22816 7962 22820
rect 7978 22876 8042 22880
rect 7978 22820 7982 22876
rect 7982 22820 8038 22876
rect 8038 22820 8042 22876
rect 7978 22816 8042 22820
rect 8058 22876 8122 22880
rect 8058 22820 8062 22876
rect 8062 22820 8118 22876
rect 8118 22820 8122 22876
rect 8058 22816 8122 22820
rect 8138 22876 8202 22880
rect 8138 22820 8142 22876
rect 8142 22820 8198 22876
rect 8198 22820 8202 22876
rect 8138 22816 8202 22820
rect 14844 22876 14908 22880
rect 14844 22820 14848 22876
rect 14848 22820 14904 22876
rect 14904 22820 14908 22876
rect 14844 22816 14908 22820
rect 14924 22876 14988 22880
rect 14924 22820 14928 22876
rect 14928 22820 14984 22876
rect 14984 22820 14988 22876
rect 14924 22816 14988 22820
rect 15004 22876 15068 22880
rect 15004 22820 15008 22876
rect 15008 22820 15064 22876
rect 15064 22820 15068 22876
rect 15004 22816 15068 22820
rect 15084 22876 15148 22880
rect 15084 22820 15088 22876
rect 15088 22820 15144 22876
rect 15144 22820 15148 22876
rect 15084 22816 15148 22820
rect 21790 22876 21854 22880
rect 21790 22820 21794 22876
rect 21794 22820 21850 22876
rect 21850 22820 21854 22876
rect 21790 22816 21854 22820
rect 21870 22876 21934 22880
rect 21870 22820 21874 22876
rect 21874 22820 21930 22876
rect 21930 22820 21934 22876
rect 21870 22816 21934 22820
rect 21950 22876 22014 22880
rect 21950 22820 21954 22876
rect 21954 22820 22010 22876
rect 22010 22820 22014 22876
rect 21950 22816 22014 22820
rect 22030 22876 22094 22880
rect 22030 22820 22034 22876
rect 22034 22820 22090 22876
rect 22090 22820 22094 22876
rect 22030 22816 22094 22820
rect 28736 22876 28800 22880
rect 28736 22820 28740 22876
rect 28740 22820 28796 22876
rect 28796 22820 28800 22876
rect 28736 22816 28800 22820
rect 28816 22876 28880 22880
rect 28816 22820 28820 22876
rect 28820 22820 28876 22876
rect 28876 22820 28880 22876
rect 28816 22816 28880 22820
rect 28896 22876 28960 22880
rect 28896 22820 28900 22876
rect 28900 22820 28956 22876
rect 28956 22820 28960 22876
rect 28896 22816 28960 22820
rect 28976 22876 29040 22880
rect 28976 22820 28980 22876
rect 28980 22820 29036 22876
rect 29036 22820 29040 22876
rect 28976 22816 29040 22820
rect 4425 22332 4489 22336
rect 4425 22276 4429 22332
rect 4429 22276 4485 22332
rect 4485 22276 4489 22332
rect 4425 22272 4489 22276
rect 4505 22332 4569 22336
rect 4505 22276 4509 22332
rect 4509 22276 4565 22332
rect 4565 22276 4569 22332
rect 4505 22272 4569 22276
rect 4585 22332 4649 22336
rect 4585 22276 4589 22332
rect 4589 22276 4645 22332
rect 4645 22276 4649 22332
rect 4585 22272 4649 22276
rect 4665 22332 4729 22336
rect 4665 22276 4669 22332
rect 4669 22276 4725 22332
rect 4725 22276 4729 22332
rect 4665 22272 4729 22276
rect 11371 22332 11435 22336
rect 11371 22276 11375 22332
rect 11375 22276 11431 22332
rect 11431 22276 11435 22332
rect 11371 22272 11435 22276
rect 11451 22332 11515 22336
rect 11451 22276 11455 22332
rect 11455 22276 11511 22332
rect 11511 22276 11515 22332
rect 11451 22272 11515 22276
rect 11531 22332 11595 22336
rect 11531 22276 11535 22332
rect 11535 22276 11591 22332
rect 11591 22276 11595 22332
rect 11531 22272 11595 22276
rect 11611 22332 11675 22336
rect 11611 22276 11615 22332
rect 11615 22276 11671 22332
rect 11671 22276 11675 22332
rect 11611 22272 11675 22276
rect 18317 22332 18381 22336
rect 18317 22276 18321 22332
rect 18321 22276 18377 22332
rect 18377 22276 18381 22332
rect 18317 22272 18381 22276
rect 18397 22332 18461 22336
rect 18397 22276 18401 22332
rect 18401 22276 18457 22332
rect 18457 22276 18461 22332
rect 18397 22272 18461 22276
rect 18477 22332 18541 22336
rect 18477 22276 18481 22332
rect 18481 22276 18537 22332
rect 18537 22276 18541 22332
rect 18477 22272 18541 22276
rect 18557 22332 18621 22336
rect 18557 22276 18561 22332
rect 18561 22276 18617 22332
rect 18617 22276 18621 22332
rect 18557 22272 18621 22276
rect 25263 22332 25327 22336
rect 25263 22276 25267 22332
rect 25267 22276 25323 22332
rect 25323 22276 25327 22332
rect 25263 22272 25327 22276
rect 25343 22332 25407 22336
rect 25343 22276 25347 22332
rect 25347 22276 25403 22332
rect 25403 22276 25407 22332
rect 25343 22272 25407 22276
rect 25423 22332 25487 22336
rect 25423 22276 25427 22332
rect 25427 22276 25483 22332
rect 25483 22276 25487 22332
rect 25423 22272 25487 22276
rect 25503 22332 25567 22336
rect 25503 22276 25507 22332
rect 25507 22276 25563 22332
rect 25563 22276 25567 22332
rect 25503 22272 25567 22276
rect 7898 21788 7962 21792
rect 7898 21732 7902 21788
rect 7902 21732 7958 21788
rect 7958 21732 7962 21788
rect 7898 21728 7962 21732
rect 7978 21788 8042 21792
rect 7978 21732 7982 21788
rect 7982 21732 8038 21788
rect 8038 21732 8042 21788
rect 7978 21728 8042 21732
rect 8058 21788 8122 21792
rect 8058 21732 8062 21788
rect 8062 21732 8118 21788
rect 8118 21732 8122 21788
rect 8058 21728 8122 21732
rect 8138 21788 8202 21792
rect 8138 21732 8142 21788
rect 8142 21732 8198 21788
rect 8198 21732 8202 21788
rect 8138 21728 8202 21732
rect 14844 21788 14908 21792
rect 14844 21732 14848 21788
rect 14848 21732 14904 21788
rect 14904 21732 14908 21788
rect 14844 21728 14908 21732
rect 14924 21788 14988 21792
rect 14924 21732 14928 21788
rect 14928 21732 14984 21788
rect 14984 21732 14988 21788
rect 14924 21728 14988 21732
rect 15004 21788 15068 21792
rect 15004 21732 15008 21788
rect 15008 21732 15064 21788
rect 15064 21732 15068 21788
rect 15004 21728 15068 21732
rect 15084 21788 15148 21792
rect 15084 21732 15088 21788
rect 15088 21732 15144 21788
rect 15144 21732 15148 21788
rect 15084 21728 15148 21732
rect 21790 21788 21854 21792
rect 21790 21732 21794 21788
rect 21794 21732 21850 21788
rect 21850 21732 21854 21788
rect 21790 21728 21854 21732
rect 21870 21788 21934 21792
rect 21870 21732 21874 21788
rect 21874 21732 21930 21788
rect 21930 21732 21934 21788
rect 21870 21728 21934 21732
rect 21950 21788 22014 21792
rect 21950 21732 21954 21788
rect 21954 21732 22010 21788
rect 22010 21732 22014 21788
rect 21950 21728 22014 21732
rect 22030 21788 22094 21792
rect 22030 21732 22034 21788
rect 22034 21732 22090 21788
rect 22090 21732 22094 21788
rect 22030 21728 22094 21732
rect 28736 21788 28800 21792
rect 28736 21732 28740 21788
rect 28740 21732 28796 21788
rect 28796 21732 28800 21788
rect 28736 21728 28800 21732
rect 28816 21788 28880 21792
rect 28816 21732 28820 21788
rect 28820 21732 28876 21788
rect 28876 21732 28880 21788
rect 28816 21728 28880 21732
rect 28896 21788 28960 21792
rect 28896 21732 28900 21788
rect 28900 21732 28956 21788
rect 28956 21732 28960 21788
rect 28896 21728 28960 21732
rect 28976 21788 29040 21792
rect 28976 21732 28980 21788
rect 28980 21732 29036 21788
rect 29036 21732 29040 21788
rect 28976 21728 29040 21732
rect 4425 21244 4489 21248
rect 4425 21188 4429 21244
rect 4429 21188 4485 21244
rect 4485 21188 4489 21244
rect 4425 21184 4489 21188
rect 4505 21244 4569 21248
rect 4505 21188 4509 21244
rect 4509 21188 4565 21244
rect 4565 21188 4569 21244
rect 4505 21184 4569 21188
rect 4585 21244 4649 21248
rect 4585 21188 4589 21244
rect 4589 21188 4645 21244
rect 4645 21188 4649 21244
rect 4585 21184 4649 21188
rect 4665 21244 4729 21248
rect 4665 21188 4669 21244
rect 4669 21188 4725 21244
rect 4725 21188 4729 21244
rect 4665 21184 4729 21188
rect 11371 21244 11435 21248
rect 11371 21188 11375 21244
rect 11375 21188 11431 21244
rect 11431 21188 11435 21244
rect 11371 21184 11435 21188
rect 11451 21244 11515 21248
rect 11451 21188 11455 21244
rect 11455 21188 11511 21244
rect 11511 21188 11515 21244
rect 11451 21184 11515 21188
rect 11531 21244 11595 21248
rect 11531 21188 11535 21244
rect 11535 21188 11591 21244
rect 11591 21188 11595 21244
rect 11531 21184 11595 21188
rect 11611 21244 11675 21248
rect 11611 21188 11615 21244
rect 11615 21188 11671 21244
rect 11671 21188 11675 21244
rect 11611 21184 11675 21188
rect 18317 21244 18381 21248
rect 18317 21188 18321 21244
rect 18321 21188 18377 21244
rect 18377 21188 18381 21244
rect 18317 21184 18381 21188
rect 18397 21244 18461 21248
rect 18397 21188 18401 21244
rect 18401 21188 18457 21244
rect 18457 21188 18461 21244
rect 18397 21184 18461 21188
rect 18477 21244 18541 21248
rect 18477 21188 18481 21244
rect 18481 21188 18537 21244
rect 18537 21188 18541 21244
rect 18477 21184 18541 21188
rect 18557 21244 18621 21248
rect 18557 21188 18561 21244
rect 18561 21188 18617 21244
rect 18617 21188 18621 21244
rect 18557 21184 18621 21188
rect 25263 21244 25327 21248
rect 25263 21188 25267 21244
rect 25267 21188 25323 21244
rect 25323 21188 25327 21244
rect 25263 21184 25327 21188
rect 25343 21244 25407 21248
rect 25343 21188 25347 21244
rect 25347 21188 25403 21244
rect 25403 21188 25407 21244
rect 25343 21184 25407 21188
rect 25423 21244 25487 21248
rect 25423 21188 25427 21244
rect 25427 21188 25483 21244
rect 25483 21188 25487 21244
rect 25423 21184 25487 21188
rect 25503 21244 25567 21248
rect 25503 21188 25507 21244
rect 25507 21188 25563 21244
rect 25563 21188 25567 21244
rect 25503 21184 25567 21188
rect 7898 20700 7962 20704
rect 7898 20644 7902 20700
rect 7902 20644 7958 20700
rect 7958 20644 7962 20700
rect 7898 20640 7962 20644
rect 7978 20700 8042 20704
rect 7978 20644 7982 20700
rect 7982 20644 8038 20700
rect 8038 20644 8042 20700
rect 7978 20640 8042 20644
rect 8058 20700 8122 20704
rect 8058 20644 8062 20700
rect 8062 20644 8118 20700
rect 8118 20644 8122 20700
rect 8058 20640 8122 20644
rect 8138 20700 8202 20704
rect 8138 20644 8142 20700
rect 8142 20644 8198 20700
rect 8198 20644 8202 20700
rect 8138 20640 8202 20644
rect 14844 20700 14908 20704
rect 14844 20644 14848 20700
rect 14848 20644 14904 20700
rect 14904 20644 14908 20700
rect 14844 20640 14908 20644
rect 14924 20700 14988 20704
rect 14924 20644 14928 20700
rect 14928 20644 14984 20700
rect 14984 20644 14988 20700
rect 14924 20640 14988 20644
rect 15004 20700 15068 20704
rect 15004 20644 15008 20700
rect 15008 20644 15064 20700
rect 15064 20644 15068 20700
rect 15004 20640 15068 20644
rect 15084 20700 15148 20704
rect 15084 20644 15088 20700
rect 15088 20644 15144 20700
rect 15144 20644 15148 20700
rect 15084 20640 15148 20644
rect 21790 20700 21854 20704
rect 21790 20644 21794 20700
rect 21794 20644 21850 20700
rect 21850 20644 21854 20700
rect 21790 20640 21854 20644
rect 21870 20700 21934 20704
rect 21870 20644 21874 20700
rect 21874 20644 21930 20700
rect 21930 20644 21934 20700
rect 21870 20640 21934 20644
rect 21950 20700 22014 20704
rect 21950 20644 21954 20700
rect 21954 20644 22010 20700
rect 22010 20644 22014 20700
rect 21950 20640 22014 20644
rect 22030 20700 22094 20704
rect 22030 20644 22034 20700
rect 22034 20644 22090 20700
rect 22090 20644 22094 20700
rect 22030 20640 22094 20644
rect 28736 20700 28800 20704
rect 28736 20644 28740 20700
rect 28740 20644 28796 20700
rect 28796 20644 28800 20700
rect 28736 20640 28800 20644
rect 28816 20700 28880 20704
rect 28816 20644 28820 20700
rect 28820 20644 28876 20700
rect 28876 20644 28880 20700
rect 28816 20640 28880 20644
rect 28896 20700 28960 20704
rect 28896 20644 28900 20700
rect 28900 20644 28956 20700
rect 28956 20644 28960 20700
rect 28896 20640 28960 20644
rect 28976 20700 29040 20704
rect 28976 20644 28980 20700
rect 28980 20644 29036 20700
rect 29036 20644 29040 20700
rect 28976 20640 29040 20644
rect 4425 20156 4489 20160
rect 4425 20100 4429 20156
rect 4429 20100 4485 20156
rect 4485 20100 4489 20156
rect 4425 20096 4489 20100
rect 4505 20156 4569 20160
rect 4505 20100 4509 20156
rect 4509 20100 4565 20156
rect 4565 20100 4569 20156
rect 4505 20096 4569 20100
rect 4585 20156 4649 20160
rect 4585 20100 4589 20156
rect 4589 20100 4645 20156
rect 4645 20100 4649 20156
rect 4585 20096 4649 20100
rect 4665 20156 4729 20160
rect 4665 20100 4669 20156
rect 4669 20100 4725 20156
rect 4725 20100 4729 20156
rect 4665 20096 4729 20100
rect 11371 20156 11435 20160
rect 11371 20100 11375 20156
rect 11375 20100 11431 20156
rect 11431 20100 11435 20156
rect 11371 20096 11435 20100
rect 11451 20156 11515 20160
rect 11451 20100 11455 20156
rect 11455 20100 11511 20156
rect 11511 20100 11515 20156
rect 11451 20096 11515 20100
rect 11531 20156 11595 20160
rect 11531 20100 11535 20156
rect 11535 20100 11591 20156
rect 11591 20100 11595 20156
rect 11531 20096 11595 20100
rect 11611 20156 11675 20160
rect 11611 20100 11615 20156
rect 11615 20100 11671 20156
rect 11671 20100 11675 20156
rect 11611 20096 11675 20100
rect 18317 20156 18381 20160
rect 18317 20100 18321 20156
rect 18321 20100 18377 20156
rect 18377 20100 18381 20156
rect 18317 20096 18381 20100
rect 18397 20156 18461 20160
rect 18397 20100 18401 20156
rect 18401 20100 18457 20156
rect 18457 20100 18461 20156
rect 18397 20096 18461 20100
rect 18477 20156 18541 20160
rect 18477 20100 18481 20156
rect 18481 20100 18537 20156
rect 18537 20100 18541 20156
rect 18477 20096 18541 20100
rect 18557 20156 18621 20160
rect 18557 20100 18561 20156
rect 18561 20100 18617 20156
rect 18617 20100 18621 20156
rect 18557 20096 18621 20100
rect 25263 20156 25327 20160
rect 25263 20100 25267 20156
rect 25267 20100 25323 20156
rect 25323 20100 25327 20156
rect 25263 20096 25327 20100
rect 25343 20156 25407 20160
rect 25343 20100 25347 20156
rect 25347 20100 25403 20156
rect 25403 20100 25407 20156
rect 25343 20096 25407 20100
rect 25423 20156 25487 20160
rect 25423 20100 25427 20156
rect 25427 20100 25483 20156
rect 25483 20100 25487 20156
rect 25423 20096 25487 20100
rect 25503 20156 25567 20160
rect 25503 20100 25507 20156
rect 25507 20100 25563 20156
rect 25563 20100 25567 20156
rect 25503 20096 25567 20100
rect 7898 19612 7962 19616
rect 7898 19556 7902 19612
rect 7902 19556 7958 19612
rect 7958 19556 7962 19612
rect 7898 19552 7962 19556
rect 7978 19612 8042 19616
rect 7978 19556 7982 19612
rect 7982 19556 8038 19612
rect 8038 19556 8042 19612
rect 7978 19552 8042 19556
rect 8058 19612 8122 19616
rect 8058 19556 8062 19612
rect 8062 19556 8118 19612
rect 8118 19556 8122 19612
rect 8058 19552 8122 19556
rect 8138 19612 8202 19616
rect 8138 19556 8142 19612
rect 8142 19556 8198 19612
rect 8198 19556 8202 19612
rect 8138 19552 8202 19556
rect 14844 19612 14908 19616
rect 14844 19556 14848 19612
rect 14848 19556 14904 19612
rect 14904 19556 14908 19612
rect 14844 19552 14908 19556
rect 14924 19612 14988 19616
rect 14924 19556 14928 19612
rect 14928 19556 14984 19612
rect 14984 19556 14988 19612
rect 14924 19552 14988 19556
rect 15004 19612 15068 19616
rect 15004 19556 15008 19612
rect 15008 19556 15064 19612
rect 15064 19556 15068 19612
rect 15004 19552 15068 19556
rect 15084 19612 15148 19616
rect 15084 19556 15088 19612
rect 15088 19556 15144 19612
rect 15144 19556 15148 19612
rect 15084 19552 15148 19556
rect 21790 19612 21854 19616
rect 21790 19556 21794 19612
rect 21794 19556 21850 19612
rect 21850 19556 21854 19612
rect 21790 19552 21854 19556
rect 21870 19612 21934 19616
rect 21870 19556 21874 19612
rect 21874 19556 21930 19612
rect 21930 19556 21934 19612
rect 21870 19552 21934 19556
rect 21950 19612 22014 19616
rect 21950 19556 21954 19612
rect 21954 19556 22010 19612
rect 22010 19556 22014 19612
rect 21950 19552 22014 19556
rect 22030 19612 22094 19616
rect 22030 19556 22034 19612
rect 22034 19556 22090 19612
rect 22090 19556 22094 19612
rect 22030 19552 22094 19556
rect 28736 19612 28800 19616
rect 28736 19556 28740 19612
rect 28740 19556 28796 19612
rect 28796 19556 28800 19612
rect 28736 19552 28800 19556
rect 28816 19612 28880 19616
rect 28816 19556 28820 19612
rect 28820 19556 28876 19612
rect 28876 19556 28880 19612
rect 28816 19552 28880 19556
rect 28896 19612 28960 19616
rect 28896 19556 28900 19612
rect 28900 19556 28956 19612
rect 28956 19556 28960 19612
rect 28896 19552 28960 19556
rect 28976 19612 29040 19616
rect 28976 19556 28980 19612
rect 28980 19556 29036 19612
rect 29036 19556 29040 19612
rect 28976 19552 29040 19556
rect 4425 19068 4489 19072
rect 4425 19012 4429 19068
rect 4429 19012 4485 19068
rect 4485 19012 4489 19068
rect 4425 19008 4489 19012
rect 4505 19068 4569 19072
rect 4505 19012 4509 19068
rect 4509 19012 4565 19068
rect 4565 19012 4569 19068
rect 4505 19008 4569 19012
rect 4585 19068 4649 19072
rect 4585 19012 4589 19068
rect 4589 19012 4645 19068
rect 4645 19012 4649 19068
rect 4585 19008 4649 19012
rect 4665 19068 4729 19072
rect 4665 19012 4669 19068
rect 4669 19012 4725 19068
rect 4725 19012 4729 19068
rect 4665 19008 4729 19012
rect 11371 19068 11435 19072
rect 11371 19012 11375 19068
rect 11375 19012 11431 19068
rect 11431 19012 11435 19068
rect 11371 19008 11435 19012
rect 11451 19068 11515 19072
rect 11451 19012 11455 19068
rect 11455 19012 11511 19068
rect 11511 19012 11515 19068
rect 11451 19008 11515 19012
rect 11531 19068 11595 19072
rect 11531 19012 11535 19068
rect 11535 19012 11591 19068
rect 11591 19012 11595 19068
rect 11531 19008 11595 19012
rect 11611 19068 11675 19072
rect 11611 19012 11615 19068
rect 11615 19012 11671 19068
rect 11671 19012 11675 19068
rect 11611 19008 11675 19012
rect 18317 19068 18381 19072
rect 18317 19012 18321 19068
rect 18321 19012 18377 19068
rect 18377 19012 18381 19068
rect 18317 19008 18381 19012
rect 18397 19068 18461 19072
rect 18397 19012 18401 19068
rect 18401 19012 18457 19068
rect 18457 19012 18461 19068
rect 18397 19008 18461 19012
rect 18477 19068 18541 19072
rect 18477 19012 18481 19068
rect 18481 19012 18537 19068
rect 18537 19012 18541 19068
rect 18477 19008 18541 19012
rect 18557 19068 18621 19072
rect 18557 19012 18561 19068
rect 18561 19012 18617 19068
rect 18617 19012 18621 19068
rect 18557 19008 18621 19012
rect 25263 19068 25327 19072
rect 25263 19012 25267 19068
rect 25267 19012 25323 19068
rect 25323 19012 25327 19068
rect 25263 19008 25327 19012
rect 25343 19068 25407 19072
rect 25343 19012 25347 19068
rect 25347 19012 25403 19068
rect 25403 19012 25407 19068
rect 25343 19008 25407 19012
rect 25423 19068 25487 19072
rect 25423 19012 25427 19068
rect 25427 19012 25483 19068
rect 25483 19012 25487 19068
rect 25423 19008 25487 19012
rect 25503 19068 25567 19072
rect 25503 19012 25507 19068
rect 25507 19012 25563 19068
rect 25563 19012 25567 19068
rect 25503 19008 25567 19012
rect 8340 18804 8404 18868
rect 7898 18524 7962 18528
rect 7898 18468 7902 18524
rect 7902 18468 7958 18524
rect 7958 18468 7962 18524
rect 7898 18464 7962 18468
rect 7978 18524 8042 18528
rect 7978 18468 7982 18524
rect 7982 18468 8038 18524
rect 8038 18468 8042 18524
rect 7978 18464 8042 18468
rect 8058 18524 8122 18528
rect 8058 18468 8062 18524
rect 8062 18468 8118 18524
rect 8118 18468 8122 18524
rect 8058 18464 8122 18468
rect 8138 18524 8202 18528
rect 8138 18468 8142 18524
rect 8142 18468 8198 18524
rect 8198 18468 8202 18524
rect 8138 18464 8202 18468
rect 14844 18524 14908 18528
rect 14844 18468 14848 18524
rect 14848 18468 14904 18524
rect 14904 18468 14908 18524
rect 14844 18464 14908 18468
rect 14924 18524 14988 18528
rect 14924 18468 14928 18524
rect 14928 18468 14984 18524
rect 14984 18468 14988 18524
rect 14924 18464 14988 18468
rect 15004 18524 15068 18528
rect 15004 18468 15008 18524
rect 15008 18468 15064 18524
rect 15064 18468 15068 18524
rect 15004 18464 15068 18468
rect 15084 18524 15148 18528
rect 15084 18468 15088 18524
rect 15088 18468 15144 18524
rect 15144 18468 15148 18524
rect 15084 18464 15148 18468
rect 21790 18524 21854 18528
rect 21790 18468 21794 18524
rect 21794 18468 21850 18524
rect 21850 18468 21854 18524
rect 21790 18464 21854 18468
rect 21870 18524 21934 18528
rect 21870 18468 21874 18524
rect 21874 18468 21930 18524
rect 21930 18468 21934 18524
rect 21870 18464 21934 18468
rect 21950 18524 22014 18528
rect 21950 18468 21954 18524
rect 21954 18468 22010 18524
rect 22010 18468 22014 18524
rect 21950 18464 22014 18468
rect 22030 18524 22094 18528
rect 22030 18468 22034 18524
rect 22034 18468 22090 18524
rect 22090 18468 22094 18524
rect 22030 18464 22094 18468
rect 28736 18524 28800 18528
rect 28736 18468 28740 18524
rect 28740 18468 28796 18524
rect 28796 18468 28800 18524
rect 28736 18464 28800 18468
rect 28816 18524 28880 18528
rect 28816 18468 28820 18524
rect 28820 18468 28876 18524
rect 28876 18468 28880 18524
rect 28816 18464 28880 18468
rect 28896 18524 28960 18528
rect 28896 18468 28900 18524
rect 28900 18468 28956 18524
rect 28956 18468 28960 18524
rect 28896 18464 28960 18468
rect 28976 18524 29040 18528
rect 28976 18468 28980 18524
rect 28980 18468 29036 18524
rect 29036 18468 29040 18524
rect 28976 18464 29040 18468
rect 4425 17980 4489 17984
rect 4425 17924 4429 17980
rect 4429 17924 4485 17980
rect 4485 17924 4489 17980
rect 4425 17920 4489 17924
rect 4505 17980 4569 17984
rect 4505 17924 4509 17980
rect 4509 17924 4565 17980
rect 4565 17924 4569 17980
rect 4505 17920 4569 17924
rect 4585 17980 4649 17984
rect 4585 17924 4589 17980
rect 4589 17924 4645 17980
rect 4645 17924 4649 17980
rect 4585 17920 4649 17924
rect 4665 17980 4729 17984
rect 4665 17924 4669 17980
rect 4669 17924 4725 17980
rect 4725 17924 4729 17980
rect 4665 17920 4729 17924
rect 11371 17980 11435 17984
rect 11371 17924 11375 17980
rect 11375 17924 11431 17980
rect 11431 17924 11435 17980
rect 11371 17920 11435 17924
rect 11451 17980 11515 17984
rect 11451 17924 11455 17980
rect 11455 17924 11511 17980
rect 11511 17924 11515 17980
rect 11451 17920 11515 17924
rect 11531 17980 11595 17984
rect 11531 17924 11535 17980
rect 11535 17924 11591 17980
rect 11591 17924 11595 17980
rect 11531 17920 11595 17924
rect 11611 17980 11675 17984
rect 11611 17924 11615 17980
rect 11615 17924 11671 17980
rect 11671 17924 11675 17980
rect 11611 17920 11675 17924
rect 18317 17980 18381 17984
rect 18317 17924 18321 17980
rect 18321 17924 18377 17980
rect 18377 17924 18381 17980
rect 18317 17920 18381 17924
rect 18397 17980 18461 17984
rect 18397 17924 18401 17980
rect 18401 17924 18457 17980
rect 18457 17924 18461 17980
rect 18397 17920 18461 17924
rect 18477 17980 18541 17984
rect 18477 17924 18481 17980
rect 18481 17924 18537 17980
rect 18537 17924 18541 17980
rect 18477 17920 18541 17924
rect 18557 17980 18621 17984
rect 18557 17924 18561 17980
rect 18561 17924 18617 17980
rect 18617 17924 18621 17980
rect 18557 17920 18621 17924
rect 25263 17980 25327 17984
rect 25263 17924 25267 17980
rect 25267 17924 25323 17980
rect 25323 17924 25327 17980
rect 25263 17920 25327 17924
rect 25343 17980 25407 17984
rect 25343 17924 25347 17980
rect 25347 17924 25403 17980
rect 25403 17924 25407 17980
rect 25343 17920 25407 17924
rect 25423 17980 25487 17984
rect 25423 17924 25427 17980
rect 25427 17924 25483 17980
rect 25483 17924 25487 17980
rect 25423 17920 25487 17924
rect 25503 17980 25567 17984
rect 25503 17924 25507 17980
rect 25507 17924 25563 17980
rect 25563 17924 25567 17980
rect 25503 17920 25567 17924
rect 7898 17436 7962 17440
rect 7898 17380 7902 17436
rect 7902 17380 7958 17436
rect 7958 17380 7962 17436
rect 7898 17376 7962 17380
rect 7978 17436 8042 17440
rect 7978 17380 7982 17436
rect 7982 17380 8038 17436
rect 8038 17380 8042 17436
rect 7978 17376 8042 17380
rect 8058 17436 8122 17440
rect 8058 17380 8062 17436
rect 8062 17380 8118 17436
rect 8118 17380 8122 17436
rect 8058 17376 8122 17380
rect 8138 17436 8202 17440
rect 8138 17380 8142 17436
rect 8142 17380 8198 17436
rect 8198 17380 8202 17436
rect 8138 17376 8202 17380
rect 14844 17436 14908 17440
rect 14844 17380 14848 17436
rect 14848 17380 14904 17436
rect 14904 17380 14908 17436
rect 14844 17376 14908 17380
rect 14924 17436 14988 17440
rect 14924 17380 14928 17436
rect 14928 17380 14984 17436
rect 14984 17380 14988 17436
rect 14924 17376 14988 17380
rect 15004 17436 15068 17440
rect 15004 17380 15008 17436
rect 15008 17380 15064 17436
rect 15064 17380 15068 17436
rect 15004 17376 15068 17380
rect 15084 17436 15148 17440
rect 15084 17380 15088 17436
rect 15088 17380 15144 17436
rect 15144 17380 15148 17436
rect 15084 17376 15148 17380
rect 21790 17436 21854 17440
rect 21790 17380 21794 17436
rect 21794 17380 21850 17436
rect 21850 17380 21854 17436
rect 21790 17376 21854 17380
rect 21870 17436 21934 17440
rect 21870 17380 21874 17436
rect 21874 17380 21930 17436
rect 21930 17380 21934 17436
rect 21870 17376 21934 17380
rect 21950 17436 22014 17440
rect 21950 17380 21954 17436
rect 21954 17380 22010 17436
rect 22010 17380 22014 17436
rect 21950 17376 22014 17380
rect 22030 17436 22094 17440
rect 22030 17380 22034 17436
rect 22034 17380 22090 17436
rect 22090 17380 22094 17436
rect 22030 17376 22094 17380
rect 28736 17436 28800 17440
rect 28736 17380 28740 17436
rect 28740 17380 28796 17436
rect 28796 17380 28800 17436
rect 28736 17376 28800 17380
rect 28816 17436 28880 17440
rect 28816 17380 28820 17436
rect 28820 17380 28876 17436
rect 28876 17380 28880 17436
rect 28816 17376 28880 17380
rect 28896 17436 28960 17440
rect 28896 17380 28900 17436
rect 28900 17380 28956 17436
rect 28956 17380 28960 17436
rect 28896 17376 28960 17380
rect 28976 17436 29040 17440
rect 28976 17380 28980 17436
rect 28980 17380 29036 17436
rect 29036 17380 29040 17436
rect 28976 17376 29040 17380
rect 4425 16892 4489 16896
rect 4425 16836 4429 16892
rect 4429 16836 4485 16892
rect 4485 16836 4489 16892
rect 4425 16832 4489 16836
rect 4505 16892 4569 16896
rect 4505 16836 4509 16892
rect 4509 16836 4565 16892
rect 4565 16836 4569 16892
rect 4505 16832 4569 16836
rect 4585 16892 4649 16896
rect 4585 16836 4589 16892
rect 4589 16836 4645 16892
rect 4645 16836 4649 16892
rect 4585 16832 4649 16836
rect 4665 16892 4729 16896
rect 4665 16836 4669 16892
rect 4669 16836 4725 16892
rect 4725 16836 4729 16892
rect 4665 16832 4729 16836
rect 11371 16892 11435 16896
rect 11371 16836 11375 16892
rect 11375 16836 11431 16892
rect 11431 16836 11435 16892
rect 11371 16832 11435 16836
rect 11451 16892 11515 16896
rect 11451 16836 11455 16892
rect 11455 16836 11511 16892
rect 11511 16836 11515 16892
rect 11451 16832 11515 16836
rect 11531 16892 11595 16896
rect 11531 16836 11535 16892
rect 11535 16836 11591 16892
rect 11591 16836 11595 16892
rect 11531 16832 11595 16836
rect 11611 16892 11675 16896
rect 11611 16836 11615 16892
rect 11615 16836 11671 16892
rect 11671 16836 11675 16892
rect 11611 16832 11675 16836
rect 18317 16892 18381 16896
rect 18317 16836 18321 16892
rect 18321 16836 18377 16892
rect 18377 16836 18381 16892
rect 18317 16832 18381 16836
rect 18397 16892 18461 16896
rect 18397 16836 18401 16892
rect 18401 16836 18457 16892
rect 18457 16836 18461 16892
rect 18397 16832 18461 16836
rect 18477 16892 18541 16896
rect 18477 16836 18481 16892
rect 18481 16836 18537 16892
rect 18537 16836 18541 16892
rect 18477 16832 18541 16836
rect 18557 16892 18621 16896
rect 18557 16836 18561 16892
rect 18561 16836 18617 16892
rect 18617 16836 18621 16892
rect 18557 16832 18621 16836
rect 25263 16892 25327 16896
rect 25263 16836 25267 16892
rect 25267 16836 25323 16892
rect 25323 16836 25327 16892
rect 25263 16832 25327 16836
rect 25343 16892 25407 16896
rect 25343 16836 25347 16892
rect 25347 16836 25403 16892
rect 25403 16836 25407 16892
rect 25343 16832 25407 16836
rect 25423 16892 25487 16896
rect 25423 16836 25427 16892
rect 25427 16836 25483 16892
rect 25483 16836 25487 16892
rect 25423 16832 25487 16836
rect 25503 16892 25567 16896
rect 25503 16836 25507 16892
rect 25507 16836 25563 16892
rect 25563 16836 25567 16892
rect 25503 16832 25567 16836
rect 7898 16348 7962 16352
rect 7898 16292 7902 16348
rect 7902 16292 7958 16348
rect 7958 16292 7962 16348
rect 7898 16288 7962 16292
rect 7978 16348 8042 16352
rect 7978 16292 7982 16348
rect 7982 16292 8038 16348
rect 8038 16292 8042 16348
rect 7978 16288 8042 16292
rect 8058 16348 8122 16352
rect 8058 16292 8062 16348
rect 8062 16292 8118 16348
rect 8118 16292 8122 16348
rect 8058 16288 8122 16292
rect 8138 16348 8202 16352
rect 8138 16292 8142 16348
rect 8142 16292 8198 16348
rect 8198 16292 8202 16348
rect 8138 16288 8202 16292
rect 14844 16348 14908 16352
rect 14844 16292 14848 16348
rect 14848 16292 14904 16348
rect 14904 16292 14908 16348
rect 14844 16288 14908 16292
rect 14924 16348 14988 16352
rect 14924 16292 14928 16348
rect 14928 16292 14984 16348
rect 14984 16292 14988 16348
rect 14924 16288 14988 16292
rect 15004 16348 15068 16352
rect 15004 16292 15008 16348
rect 15008 16292 15064 16348
rect 15064 16292 15068 16348
rect 15004 16288 15068 16292
rect 15084 16348 15148 16352
rect 15084 16292 15088 16348
rect 15088 16292 15144 16348
rect 15144 16292 15148 16348
rect 15084 16288 15148 16292
rect 21790 16348 21854 16352
rect 21790 16292 21794 16348
rect 21794 16292 21850 16348
rect 21850 16292 21854 16348
rect 21790 16288 21854 16292
rect 21870 16348 21934 16352
rect 21870 16292 21874 16348
rect 21874 16292 21930 16348
rect 21930 16292 21934 16348
rect 21870 16288 21934 16292
rect 21950 16348 22014 16352
rect 21950 16292 21954 16348
rect 21954 16292 22010 16348
rect 22010 16292 22014 16348
rect 21950 16288 22014 16292
rect 22030 16348 22094 16352
rect 22030 16292 22034 16348
rect 22034 16292 22090 16348
rect 22090 16292 22094 16348
rect 22030 16288 22094 16292
rect 28736 16348 28800 16352
rect 28736 16292 28740 16348
rect 28740 16292 28796 16348
rect 28796 16292 28800 16348
rect 28736 16288 28800 16292
rect 28816 16348 28880 16352
rect 28816 16292 28820 16348
rect 28820 16292 28876 16348
rect 28876 16292 28880 16348
rect 28816 16288 28880 16292
rect 28896 16348 28960 16352
rect 28896 16292 28900 16348
rect 28900 16292 28956 16348
rect 28956 16292 28960 16348
rect 28896 16288 28960 16292
rect 28976 16348 29040 16352
rect 28976 16292 28980 16348
rect 28980 16292 29036 16348
rect 29036 16292 29040 16348
rect 28976 16288 29040 16292
rect 4425 15804 4489 15808
rect 4425 15748 4429 15804
rect 4429 15748 4485 15804
rect 4485 15748 4489 15804
rect 4425 15744 4489 15748
rect 4505 15804 4569 15808
rect 4505 15748 4509 15804
rect 4509 15748 4565 15804
rect 4565 15748 4569 15804
rect 4505 15744 4569 15748
rect 4585 15804 4649 15808
rect 4585 15748 4589 15804
rect 4589 15748 4645 15804
rect 4645 15748 4649 15804
rect 4585 15744 4649 15748
rect 4665 15804 4729 15808
rect 4665 15748 4669 15804
rect 4669 15748 4725 15804
rect 4725 15748 4729 15804
rect 4665 15744 4729 15748
rect 11371 15804 11435 15808
rect 11371 15748 11375 15804
rect 11375 15748 11431 15804
rect 11431 15748 11435 15804
rect 11371 15744 11435 15748
rect 11451 15804 11515 15808
rect 11451 15748 11455 15804
rect 11455 15748 11511 15804
rect 11511 15748 11515 15804
rect 11451 15744 11515 15748
rect 11531 15804 11595 15808
rect 11531 15748 11535 15804
rect 11535 15748 11591 15804
rect 11591 15748 11595 15804
rect 11531 15744 11595 15748
rect 11611 15804 11675 15808
rect 11611 15748 11615 15804
rect 11615 15748 11671 15804
rect 11671 15748 11675 15804
rect 11611 15744 11675 15748
rect 18317 15804 18381 15808
rect 18317 15748 18321 15804
rect 18321 15748 18377 15804
rect 18377 15748 18381 15804
rect 18317 15744 18381 15748
rect 18397 15804 18461 15808
rect 18397 15748 18401 15804
rect 18401 15748 18457 15804
rect 18457 15748 18461 15804
rect 18397 15744 18461 15748
rect 18477 15804 18541 15808
rect 18477 15748 18481 15804
rect 18481 15748 18537 15804
rect 18537 15748 18541 15804
rect 18477 15744 18541 15748
rect 18557 15804 18621 15808
rect 18557 15748 18561 15804
rect 18561 15748 18617 15804
rect 18617 15748 18621 15804
rect 18557 15744 18621 15748
rect 25263 15804 25327 15808
rect 25263 15748 25267 15804
rect 25267 15748 25323 15804
rect 25323 15748 25327 15804
rect 25263 15744 25327 15748
rect 25343 15804 25407 15808
rect 25343 15748 25347 15804
rect 25347 15748 25403 15804
rect 25403 15748 25407 15804
rect 25343 15744 25407 15748
rect 25423 15804 25487 15808
rect 25423 15748 25427 15804
rect 25427 15748 25483 15804
rect 25483 15748 25487 15804
rect 25423 15744 25487 15748
rect 25503 15804 25567 15808
rect 25503 15748 25507 15804
rect 25507 15748 25563 15804
rect 25563 15748 25567 15804
rect 25503 15744 25567 15748
rect 4108 15268 4172 15332
rect 7898 15260 7962 15264
rect 7898 15204 7902 15260
rect 7902 15204 7958 15260
rect 7958 15204 7962 15260
rect 7898 15200 7962 15204
rect 7978 15260 8042 15264
rect 7978 15204 7982 15260
rect 7982 15204 8038 15260
rect 8038 15204 8042 15260
rect 7978 15200 8042 15204
rect 8058 15260 8122 15264
rect 8058 15204 8062 15260
rect 8062 15204 8118 15260
rect 8118 15204 8122 15260
rect 8058 15200 8122 15204
rect 8138 15260 8202 15264
rect 8138 15204 8142 15260
rect 8142 15204 8198 15260
rect 8198 15204 8202 15260
rect 8138 15200 8202 15204
rect 14844 15260 14908 15264
rect 14844 15204 14848 15260
rect 14848 15204 14904 15260
rect 14904 15204 14908 15260
rect 14844 15200 14908 15204
rect 14924 15260 14988 15264
rect 14924 15204 14928 15260
rect 14928 15204 14984 15260
rect 14984 15204 14988 15260
rect 14924 15200 14988 15204
rect 15004 15260 15068 15264
rect 15004 15204 15008 15260
rect 15008 15204 15064 15260
rect 15064 15204 15068 15260
rect 15004 15200 15068 15204
rect 15084 15260 15148 15264
rect 15084 15204 15088 15260
rect 15088 15204 15144 15260
rect 15144 15204 15148 15260
rect 15084 15200 15148 15204
rect 21790 15260 21854 15264
rect 21790 15204 21794 15260
rect 21794 15204 21850 15260
rect 21850 15204 21854 15260
rect 21790 15200 21854 15204
rect 21870 15260 21934 15264
rect 21870 15204 21874 15260
rect 21874 15204 21930 15260
rect 21930 15204 21934 15260
rect 21870 15200 21934 15204
rect 21950 15260 22014 15264
rect 21950 15204 21954 15260
rect 21954 15204 22010 15260
rect 22010 15204 22014 15260
rect 21950 15200 22014 15204
rect 22030 15260 22094 15264
rect 22030 15204 22034 15260
rect 22034 15204 22090 15260
rect 22090 15204 22094 15260
rect 22030 15200 22094 15204
rect 28736 15260 28800 15264
rect 28736 15204 28740 15260
rect 28740 15204 28796 15260
rect 28796 15204 28800 15260
rect 28736 15200 28800 15204
rect 28816 15260 28880 15264
rect 28816 15204 28820 15260
rect 28820 15204 28876 15260
rect 28876 15204 28880 15260
rect 28816 15200 28880 15204
rect 28896 15260 28960 15264
rect 28896 15204 28900 15260
rect 28900 15204 28956 15260
rect 28956 15204 28960 15260
rect 28896 15200 28960 15204
rect 28976 15260 29040 15264
rect 28976 15204 28980 15260
rect 28980 15204 29036 15260
rect 29036 15204 29040 15260
rect 28976 15200 29040 15204
rect 4425 14716 4489 14720
rect 4425 14660 4429 14716
rect 4429 14660 4485 14716
rect 4485 14660 4489 14716
rect 4425 14656 4489 14660
rect 4505 14716 4569 14720
rect 4505 14660 4509 14716
rect 4509 14660 4565 14716
rect 4565 14660 4569 14716
rect 4505 14656 4569 14660
rect 4585 14716 4649 14720
rect 4585 14660 4589 14716
rect 4589 14660 4645 14716
rect 4645 14660 4649 14716
rect 4585 14656 4649 14660
rect 4665 14716 4729 14720
rect 4665 14660 4669 14716
rect 4669 14660 4725 14716
rect 4725 14660 4729 14716
rect 4665 14656 4729 14660
rect 11371 14716 11435 14720
rect 11371 14660 11375 14716
rect 11375 14660 11431 14716
rect 11431 14660 11435 14716
rect 11371 14656 11435 14660
rect 11451 14716 11515 14720
rect 11451 14660 11455 14716
rect 11455 14660 11511 14716
rect 11511 14660 11515 14716
rect 11451 14656 11515 14660
rect 11531 14716 11595 14720
rect 11531 14660 11535 14716
rect 11535 14660 11591 14716
rect 11591 14660 11595 14716
rect 11531 14656 11595 14660
rect 11611 14716 11675 14720
rect 11611 14660 11615 14716
rect 11615 14660 11671 14716
rect 11671 14660 11675 14716
rect 11611 14656 11675 14660
rect 18317 14716 18381 14720
rect 18317 14660 18321 14716
rect 18321 14660 18377 14716
rect 18377 14660 18381 14716
rect 18317 14656 18381 14660
rect 18397 14716 18461 14720
rect 18397 14660 18401 14716
rect 18401 14660 18457 14716
rect 18457 14660 18461 14716
rect 18397 14656 18461 14660
rect 18477 14716 18541 14720
rect 18477 14660 18481 14716
rect 18481 14660 18537 14716
rect 18537 14660 18541 14716
rect 18477 14656 18541 14660
rect 18557 14716 18621 14720
rect 18557 14660 18561 14716
rect 18561 14660 18617 14716
rect 18617 14660 18621 14716
rect 18557 14656 18621 14660
rect 25263 14716 25327 14720
rect 25263 14660 25267 14716
rect 25267 14660 25323 14716
rect 25323 14660 25327 14716
rect 25263 14656 25327 14660
rect 25343 14716 25407 14720
rect 25343 14660 25347 14716
rect 25347 14660 25403 14716
rect 25403 14660 25407 14716
rect 25343 14656 25407 14660
rect 25423 14716 25487 14720
rect 25423 14660 25427 14716
rect 25427 14660 25483 14716
rect 25483 14660 25487 14716
rect 25423 14656 25487 14660
rect 25503 14716 25567 14720
rect 25503 14660 25507 14716
rect 25507 14660 25563 14716
rect 25563 14660 25567 14716
rect 25503 14656 25567 14660
rect 7898 14172 7962 14176
rect 7898 14116 7902 14172
rect 7902 14116 7958 14172
rect 7958 14116 7962 14172
rect 7898 14112 7962 14116
rect 7978 14172 8042 14176
rect 7978 14116 7982 14172
rect 7982 14116 8038 14172
rect 8038 14116 8042 14172
rect 7978 14112 8042 14116
rect 8058 14172 8122 14176
rect 8058 14116 8062 14172
rect 8062 14116 8118 14172
rect 8118 14116 8122 14172
rect 8058 14112 8122 14116
rect 8138 14172 8202 14176
rect 8138 14116 8142 14172
rect 8142 14116 8198 14172
rect 8198 14116 8202 14172
rect 8138 14112 8202 14116
rect 14844 14172 14908 14176
rect 14844 14116 14848 14172
rect 14848 14116 14904 14172
rect 14904 14116 14908 14172
rect 14844 14112 14908 14116
rect 14924 14172 14988 14176
rect 14924 14116 14928 14172
rect 14928 14116 14984 14172
rect 14984 14116 14988 14172
rect 14924 14112 14988 14116
rect 15004 14172 15068 14176
rect 15004 14116 15008 14172
rect 15008 14116 15064 14172
rect 15064 14116 15068 14172
rect 15004 14112 15068 14116
rect 15084 14172 15148 14176
rect 15084 14116 15088 14172
rect 15088 14116 15144 14172
rect 15144 14116 15148 14172
rect 15084 14112 15148 14116
rect 21790 14172 21854 14176
rect 21790 14116 21794 14172
rect 21794 14116 21850 14172
rect 21850 14116 21854 14172
rect 21790 14112 21854 14116
rect 21870 14172 21934 14176
rect 21870 14116 21874 14172
rect 21874 14116 21930 14172
rect 21930 14116 21934 14172
rect 21870 14112 21934 14116
rect 21950 14172 22014 14176
rect 21950 14116 21954 14172
rect 21954 14116 22010 14172
rect 22010 14116 22014 14172
rect 21950 14112 22014 14116
rect 22030 14172 22094 14176
rect 22030 14116 22034 14172
rect 22034 14116 22090 14172
rect 22090 14116 22094 14172
rect 22030 14112 22094 14116
rect 28736 14172 28800 14176
rect 28736 14116 28740 14172
rect 28740 14116 28796 14172
rect 28796 14116 28800 14172
rect 28736 14112 28800 14116
rect 28816 14172 28880 14176
rect 28816 14116 28820 14172
rect 28820 14116 28876 14172
rect 28876 14116 28880 14172
rect 28816 14112 28880 14116
rect 28896 14172 28960 14176
rect 28896 14116 28900 14172
rect 28900 14116 28956 14172
rect 28956 14116 28960 14172
rect 28896 14112 28960 14116
rect 28976 14172 29040 14176
rect 28976 14116 28980 14172
rect 28980 14116 29036 14172
rect 29036 14116 29040 14172
rect 28976 14112 29040 14116
rect 8340 13696 8404 13700
rect 8340 13640 8390 13696
rect 8390 13640 8404 13696
rect 8340 13636 8404 13640
rect 4425 13628 4489 13632
rect 4425 13572 4429 13628
rect 4429 13572 4485 13628
rect 4485 13572 4489 13628
rect 4425 13568 4489 13572
rect 4505 13628 4569 13632
rect 4505 13572 4509 13628
rect 4509 13572 4565 13628
rect 4565 13572 4569 13628
rect 4505 13568 4569 13572
rect 4585 13628 4649 13632
rect 4585 13572 4589 13628
rect 4589 13572 4645 13628
rect 4645 13572 4649 13628
rect 4585 13568 4649 13572
rect 4665 13628 4729 13632
rect 4665 13572 4669 13628
rect 4669 13572 4725 13628
rect 4725 13572 4729 13628
rect 4665 13568 4729 13572
rect 11371 13628 11435 13632
rect 11371 13572 11375 13628
rect 11375 13572 11431 13628
rect 11431 13572 11435 13628
rect 11371 13568 11435 13572
rect 11451 13628 11515 13632
rect 11451 13572 11455 13628
rect 11455 13572 11511 13628
rect 11511 13572 11515 13628
rect 11451 13568 11515 13572
rect 11531 13628 11595 13632
rect 11531 13572 11535 13628
rect 11535 13572 11591 13628
rect 11591 13572 11595 13628
rect 11531 13568 11595 13572
rect 11611 13628 11675 13632
rect 11611 13572 11615 13628
rect 11615 13572 11671 13628
rect 11671 13572 11675 13628
rect 11611 13568 11675 13572
rect 18317 13628 18381 13632
rect 18317 13572 18321 13628
rect 18321 13572 18377 13628
rect 18377 13572 18381 13628
rect 18317 13568 18381 13572
rect 18397 13628 18461 13632
rect 18397 13572 18401 13628
rect 18401 13572 18457 13628
rect 18457 13572 18461 13628
rect 18397 13568 18461 13572
rect 18477 13628 18541 13632
rect 18477 13572 18481 13628
rect 18481 13572 18537 13628
rect 18537 13572 18541 13628
rect 18477 13568 18541 13572
rect 18557 13628 18621 13632
rect 18557 13572 18561 13628
rect 18561 13572 18617 13628
rect 18617 13572 18621 13628
rect 18557 13568 18621 13572
rect 25263 13628 25327 13632
rect 25263 13572 25267 13628
rect 25267 13572 25323 13628
rect 25323 13572 25327 13628
rect 25263 13568 25327 13572
rect 25343 13628 25407 13632
rect 25343 13572 25347 13628
rect 25347 13572 25403 13628
rect 25403 13572 25407 13628
rect 25343 13568 25407 13572
rect 25423 13628 25487 13632
rect 25423 13572 25427 13628
rect 25427 13572 25483 13628
rect 25483 13572 25487 13628
rect 25423 13568 25487 13572
rect 25503 13628 25567 13632
rect 25503 13572 25507 13628
rect 25507 13572 25563 13628
rect 25563 13572 25567 13628
rect 25503 13568 25567 13572
rect 7898 13084 7962 13088
rect 7898 13028 7902 13084
rect 7902 13028 7958 13084
rect 7958 13028 7962 13084
rect 7898 13024 7962 13028
rect 7978 13084 8042 13088
rect 7978 13028 7982 13084
rect 7982 13028 8038 13084
rect 8038 13028 8042 13084
rect 7978 13024 8042 13028
rect 8058 13084 8122 13088
rect 8058 13028 8062 13084
rect 8062 13028 8118 13084
rect 8118 13028 8122 13084
rect 8058 13024 8122 13028
rect 8138 13084 8202 13088
rect 8138 13028 8142 13084
rect 8142 13028 8198 13084
rect 8198 13028 8202 13084
rect 8138 13024 8202 13028
rect 14844 13084 14908 13088
rect 14844 13028 14848 13084
rect 14848 13028 14904 13084
rect 14904 13028 14908 13084
rect 14844 13024 14908 13028
rect 14924 13084 14988 13088
rect 14924 13028 14928 13084
rect 14928 13028 14984 13084
rect 14984 13028 14988 13084
rect 14924 13024 14988 13028
rect 15004 13084 15068 13088
rect 15004 13028 15008 13084
rect 15008 13028 15064 13084
rect 15064 13028 15068 13084
rect 15004 13024 15068 13028
rect 15084 13084 15148 13088
rect 15084 13028 15088 13084
rect 15088 13028 15144 13084
rect 15144 13028 15148 13084
rect 15084 13024 15148 13028
rect 21790 13084 21854 13088
rect 21790 13028 21794 13084
rect 21794 13028 21850 13084
rect 21850 13028 21854 13084
rect 21790 13024 21854 13028
rect 21870 13084 21934 13088
rect 21870 13028 21874 13084
rect 21874 13028 21930 13084
rect 21930 13028 21934 13084
rect 21870 13024 21934 13028
rect 21950 13084 22014 13088
rect 21950 13028 21954 13084
rect 21954 13028 22010 13084
rect 22010 13028 22014 13084
rect 21950 13024 22014 13028
rect 22030 13084 22094 13088
rect 22030 13028 22034 13084
rect 22034 13028 22090 13084
rect 22090 13028 22094 13084
rect 22030 13024 22094 13028
rect 28736 13084 28800 13088
rect 28736 13028 28740 13084
rect 28740 13028 28796 13084
rect 28796 13028 28800 13084
rect 28736 13024 28800 13028
rect 28816 13084 28880 13088
rect 28816 13028 28820 13084
rect 28820 13028 28876 13084
rect 28876 13028 28880 13084
rect 28816 13024 28880 13028
rect 28896 13084 28960 13088
rect 28896 13028 28900 13084
rect 28900 13028 28956 13084
rect 28956 13028 28960 13084
rect 28896 13024 28960 13028
rect 28976 13084 29040 13088
rect 28976 13028 28980 13084
rect 28980 13028 29036 13084
rect 29036 13028 29040 13084
rect 28976 13024 29040 13028
rect 4425 12540 4489 12544
rect 4425 12484 4429 12540
rect 4429 12484 4485 12540
rect 4485 12484 4489 12540
rect 4425 12480 4489 12484
rect 4505 12540 4569 12544
rect 4505 12484 4509 12540
rect 4509 12484 4565 12540
rect 4565 12484 4569 12540
rect 4505 12480 4569 12484
rect 4585 12540 4649 12544
rect 4585 12484 4589 12540
rect 4589 12484 4645 12540
rect 4645 12484 4649 12540
rect 4585 12480 4649 12484
rect 4665 12540 4729 12544
rect 4665 12484 4669 12540
rect 4669 12484 4725 12540
rect 4725 12484 4729 12540
rect 4665 12480 4729 12484
rect 11371 12540 11435 12544
rect 11371 12484 11375 12540
rect 11375 12484 11431 12540
rect 11431 12484 11435 12540
rect 11371 12480 11435 12484
rect 11451 12540 11515 12544
rect 11451 12484 11455 12540
rect 11455 12484 11511 12540
rect 11511 12484 11515 12540
rect 11451 12480 11515 12484
rect 11531 12540 11595 12544
rect 11531 12484 11535 12540
rect 11535 12484 11591 12540
rect 11591 12484 11595 12540
rect 11531 12480 11595 12484
rect 11611 12540 11675 12544
rect 11611 12484 11615 12540
rect 11615 12484 11671 12540
rect 11671 12484 11675 12540
rect 11611 12480 11675 12484
rect 18317 12540 18381 12544
rect 18317 12484 18321 12540
rect 18321 12484 18377 12540
rect 18377 12484 18381 12540
rect 18317 12480 18381 12484
rect 18397 12540 18461 12544
rect 18397 12484 18401 12540
rect 18401 12484 18457 12540
rect 18457 12484 18461 12540
rect 18397 12480 18461 12484
rect 18477 12540 18541 12544
rect 18477 12484 18481 12540
rect 18481 12484 18537 12540
rect 18537 12484 18541 12540
rect 18477 12480 18541 12484
rect 18557 12540 18621 12544
rect 18557 12484 18561 12540
rect 18561 12484 18617 12540
rect 18617 12484 18621 12540
rect 18557 12480 18621 12484
rect 25263 12540 25327 12544
rect 25263 12484 25267 12540
rect 25267 12484 25323 12540
rect 25323 12484 25327 12540
rect 25263 12480 25327 12484
rect 25343 12540 25407 12544
rect 25343 12484 25347 12540
rect 25347 12484 25403 12540
rect 25403 12484 25407 12540
rect 25343 12480 25407 12484
rect 25423 12540 25487 12544
rect 25423 12484 25427 12540
rect 25427 12484 25483 12540
rect 25483 12484 25487 12540
rect 25423 12480 25487 12484
rect 25503 12540 25567 12544
rect 25503 12484 25507 12540
rect 25507 12484 25563 12540
rect 25563 12484 25567 12540
rect 25503 12480 25567 12484
rect 7898 11996 7962 12000
rect 7898 11940 7902 11996
rect 7902 11940 7958 11996
rect 7958 11940 7962 11996
rect 7898 11936 7962 11940
rect 7978 11996 8042 12000
rect 7978 11940 7982 11996
rect 7982 11940 8038 11996
rect 8038 11940 8042 11996
rect 7978 11936 8042 11940
rect 8058 11996 8122 12000
rect 8058 11940 8062 11996
rect 8062 11940 8118 11996
rect 8118 11940 8122 11996
rect 8058 11936 8122 11940
rect 8138 11996 8202 12000
rect 8138 11940 8142 11996
rect 8142 11940 8198 11996
rect 8198 11940 8202 11996
rect 8138 11936 8202 11940
rect 14844 11996 14908 12000
rect 14844 11940 14848 11996
rect 14848 11940 14904 11996
rect 14904 11940 14908 11996
rect 14844 11936 14908 11940
rect 14924 11996 14988 12000
rect 14924 11940 14928 11996
rect 14928 11940 14984 11996
rect 14984 11940 14988 11996
rect 14924 11936 14988 11940
rect 15004 11996 15068 12000
rect 15004 11940 15008 11996
rect 15008 11940 15064 11996
rect 15064 11940 15068 11996
rect 15004 11936 15068 11940
rect 15084 11996 15148 12000
rect 15084 11940 15088 11996
rect 15088 11940 15144 11996
rect 15144 11940 15148 11996
rect 15084 11936 15148 11940
rect 21790 11996 21854 12000
rect 21790 11940 21794 11996
rect 21794 11940 21850 11996
rect 21850 11940 21854 11996
rect 21790 11936 21854 11940
rect 21870 11996 21934 12000
rect 21870 11940 21874 11996
rect 21874 11940 21930 11996
rect 21930 11940 21934 11996
rect 21870 11936 21934 11940
rect 21950 11996 22014 12000
rect 21950 11940 21954 11996
rect 21954 11940 22010 11996
rect 22010 11940 22014 11996
rect 21950 11936 22014 11940
rect 22030 11996 22094 12000
rect 22030 11940 22034 11996
rect 22034 11940 22090 11996
rect 22090 11940 22094 11996
rect 22030 11936 22094 11940
rect 28736 11996 28800 12000
rect 28736 11940 28740 11996
rect 28740 11940 28796 11996
rect 28796 11940 28800 11996
rect 28736 11936 28800 11940
rect 28816 11996 28880 12000
rect 28816 11940 28820 11996
rect 28820 11940 28876 11996
rect 28876 11940 28880 11996
rect 28816 11936 28880 11940
rect 28896 11996 28960 12000
rect 28896 11940 28900 11996
rect 28900 11940 28956 11996
rect 28956 11940 28960 11996
rect 28896 11936 28960 11940
rect 28976 11996 29040 12000
rect 28976 11940 28980 11996
rect 28980 11940 29036 11996
rect 29036 11940 29040 11996
rect 28976 11936 29040 11940
rect 4425 11452 4489 11456
rect 4425 11396 4429 11452
rect 4429 11396 4485 11452
rect 4485 11396 4489 11452
rect 4425 11392 4489 11396
rect 4505 11452 4569 11456
rect 4505 11396 4509 11452
rect 4509 11396 4565 11452
rect 4565 11396 4569 11452
rect 4505 11392 4569 11396
rect 4585 11452 4649 11456
rect 4585 11396 4589 11452
rect 4589 11396 4645 11452
rect 4645 11396 4649 11452
rect 4585 11392 4649 11396
rect 4665 11452 4729 11456
rect 4665 11396 4669 11452
rect 4669 11396 4725 11452
rect 4725 11396 4729 11452
rect 4665 11392 4729 11396
rect 11371 11452 11435 11456
rect 11371 11396 11375 11452
rect 11375 11396 11431 11452
rect 11431 11396 11435 11452
rect 11371 11392 11435 11396
rect 11451 11452 11515 11456
rect 11451 11396 11455 11452
rect 11455 11396 11511 11452
rect 11511 11396 11515 11452
rect 11451 11392 11515 11396
rect 11531 11452 11595 11456
rect 11531 11396 11535 11452
rect 11535 11396 11591 11452
rect 11591 11396 11595 11452
rect 11531 11392 11595 11396
rect 11611 11452 11675 11456
rect 11611 11396 11615 11452
rect 11615 11396 11671 11452
rect 11671 11396 11675 11452
rect 11611 11392 11675 11396
rect 18317 11452 18381 11456
rect 18317 11396 18321 11452
rect 18321 11396 18377 11452
rect 18377 11396 18381 11452
rect 18317 11392 18381 11396
rect 18397 11452 18461 11456
rect 18397 11396 18401 11452
rect 18401 11396 18457 11452
rect 18457 11396 18461 11452
rect 18397 11392 18461 11396
rect 18477 11452 18541 11456
rect 18477 11396 18481 11452
rect 18481 11396 18537 11452
rect 18537 11396 18541 11452
rect 18477 11392 18541 11396
rect 18557 11452 18621 11456
rect 18557 11396 18561 11452
rect 18561 11396 18617 11452
rect 18617 11396 18621 11452
rect 18557 11392 18621 11396
rect 25263 11452 25327 11456
rect 25263 11396 25267 11452
rect 25267 11396 25323 11452
rect 25323 11396 25327 11452
rect 25263 11392 25327 11396
rect 25343 11452 25407 11456
rect 25343 11396 25347 11452
rect 25347 11396 25403 11452
rect 25403 11396 25407 11452
rect 25343 11392 25407 11396
rect 25423 11452 25487 11456
rect 25423 11396 25427 11452
rect 25427 11396 25483 11452
rect 25483 11396 25487 11452
rect 25423 11392 25487 11396
rect 25503 11452 25567 11456
rect 25503 11396 25507 11452
rect 25507 11396 25563 11452
rect 25563 11396 25567 11452
rect 25503 11392 25567 11396
rect 7898 10908 7962 10912
rect 7898 10852 7902 10908
rect 7902 10852 7958 10908
rect 7958 10852 7962 10908
rect 7898 10848 7962 10852
rect 7978 10908 8042 10912
rect 7978 10852 7982 10908
rect 7982 10852 8038 10908
rect 8038 10852 8042 10908
rect 7978 10848 8042 10852
rect 8058 10908 8122 10912
rect 8058 10852 8062 10908
rect 8062 10852 8118 10908
rect 8118 10852 8122 10908
rect 8058 10848 8122 10852
rect 8138 10908 8202 10912
rect 8138 10852 8142 10908
rect 8142 10852 8198 10908
rect 8198 10852 8202 10908
rect 8138 10848 8202 10852
rect 14844 10908 14908 10912
rect 14844 10852 14848 10908
rect 14848 10852 14904 10908
rect 14904 10852 14908 10908
rect 14844 10848 14908 10852
rect 14924 10908 14988 10912
rect 14924 10852 14928 10908
rect 14928 10852 14984 10908
rect 14984 10852 14988 10908
rect 14924 10848 14988 10852
rect 15004 10908 15068 10912
rect 15004 10852 15008 10908
rect 15008 10852 15064 10908
rect 15064 10852 15068 10908
rect 15004 10848 15068 10852
rect 15084 10908 15148 10912
rect 15084 10852 15088 10908
rect 15088 10852 15144 10908
rect 15144 10852 15148 10908
rect 15084 10848 15148 10852
rect 21790 10908 21854 10912
rect 21790 10852 21794 10908
rect 21794 10852 21850 10908
rect 21850 10852 21854 10908
rect 21790 10848 21854 10852
rect 21870 10908 21934 10912
rect 21870 10852 21874 10908
rect 21874 10852 21930 10908
rect 21930 10852 21934 10908
rect 21870 10848 21934 10852
rect 21950 10908 22014 10912
rect 21950 10852 21954 10908
rect 21954 10852 22010 10908
rect 22010 10852 22014 10908
rect 21950 10848 22014 10852
rect 22030 10908 22094 10912
rect 22030 10852 22034 10908
rect 22034 10852 22090 10908
rect 22090 10852 22094 10908
rect 22030 10848 22094 10852
rect 28736 10908 28800 10912
rect 28736 10852 28740 10908
rect 28740 10852 28796 10908
rect 28796 10852 28800 10908
rect 28736 10848 28800 10852
rect 28816 10908 28880 10912
rect 28816 10852 28820 10908
rect 28820 10852 28876 10908
rect 28876 10852 28880 10908
rect 28816 10848 28880 10852
rect 28896 10908 28960 10912
rect 28896 10852 28900 10908
rect 28900 10852 28956 10908
rect 28956 10852 28960 10908
rect 28896 10848 28960 10852
rect 28976 10908 29040 10912
rect 28976 10852 28980 10908
rect 28980 10852 29036 10908
rect 29036 10852 29040 10908
rect 28976 10848 29040 10852
rect 4425 10364 4489 10368
rect 4425 10308 4429 10364
rect 4429 10308 4485 10364
rect 4485 10308 4489 10364
rect 4425 10304 4489 10308
rect 4505 10364 4569 10368
rect 4505 10308 4509 10364
rect 4509 10308 4565 10364
rect 4565 10308 4569 10364
rect 4505 10304 4569 10308
rect 4585 10364 4649 10368
rect 4585 10308 4589 10364
rect 4589 10308 4645 10364
rect 4645 10308 4649 10364
rect 4585 10304 4649 10308
rect 4665 10364 4729 10368
rect 4665 10308 4669 10364
rect 4669 10308 4725 10364
rect 4725 10308 4729 10364
rect 4665 10304 4729 10308
rect 11371 10364 11435 10368
rect 11371 10308 11375 10364
rect 11375 10308 11431 10364
rect 11431 10308 11435 10364
rect 11371 10304 11435 10308
rect 11451 10364 11515 10368
rect 11451 10308 11455 10364
rect 11455 10308 11511 10364
rect 11511 10308 11515 10364
rect 11451 10304 11515 10308
rect 11531 10364 11595 10368
rect 11531 10308 11535 10364
rect 11535 10308 11591 10364
rect 11591 10308 11595 10364
rect 11531 10304 11595 10308
rect 11611 10364 11675 10368
rect 11611 10308 11615 10364
rect 11615 10308 11671 10364
rect 11671 10308 11675 10364
rect 11611 10304 11675 10308
rect 18317 10364 18381 10368
rect 18317 10308 18321 10364
rect 18321 10308 18377 10364
rect 18377 10308 18381 10364
rect 18317 10304 18381 10308
rect 18397 10364 18461 10368
rect 18397 10308 18401 10364
rect 18401 10308 18457 10364
rect 18457 10308 18461 10364
rect 18397 10304 18461 10308
rect 18477 10364 18541 10368
rect 18477 10308 18481 10364
rect 18481 10308 18537 10364
rect 18537 10308 18541 10364
rect 18477 10304 18541 10308
rect 18557 10364 18621 10368
rect 18557 10308 18561 10364
rect 18561 10308 18617 10364
rect 18617 10308 18621 10364
rect 18557 10304 18621 10308
rect 25263 10364 25327 10368
rect 25263 10308 25267 10364
rect 25267 10308 25323 10364
rect 25323 10308 25327 10364
rect 25263 10304 25327 10308
rect 25343 10364 25407 10368
rect 25343 10308 25347 10364
rect 25347 10308 25403 10364
rect 25403 10308 25407 10364
rect 25343 10304 25407 10308
rect 25423 10364 25487 10368
rect 25423 10308 25427 10364
rect 25427 10308 25483 10364
rect 25483 10308 25487 10364
rect 25423 10304 25487 10308
rect 25503 10364 25567 10368
rect 25503 10308 25507 10364
rect 25507 10308 25563 10364
rect 25563 10308 25567 10364
rect 25503 10304 25567 10308
rect 7898 9820 7962 9824
rect 7898 9764 7902 9820
rect 7902 9764 7958 9820
rect 7958 9764 7962 9820
rect 7898 9760 7962 9764
rect 7978 9820 8042 9824
rect 7978 9764 7982 9820
rect 7982 9764 8038 9820
rect 8038 9764 8042 9820
rect 7978 9760 8042 9764
rect 8058 9820 8122 9824
rect 8058 9764 8062 9820
rect 8062 9764 8118 9820
rect 8118 9764 8122 9820
rect 8058 9760 8122 9764
rect 8138 9820 8202 9824
rect 8138 9764 8142 9820
rect 8142 9764 8198 9820
rect 8198 9764 8202 9820
rect 8138 9760 8202 9764
rect 14844 9820 14908 9824
rect 14844 9764 14848 9820
rect 14848 9764 14904 9820
rect 14904 9764 14908 9820
rect 14844 9760 14908 9764
rect 14924 9820 14988 9824
rect 14924 9764 14928 9820
rect 14928 9764 14984 9820
rect 14984 9764 14988 9820
rect 14924 9760 14988 9764
rect 15004 9820 15068 9824
rect 15004 9764 15008 9820
rect 15008 9764 15064 9820
rect 15064 9764 15068 9820
rect 15004 9760 15068 9764
rect 15084 9820 15148 9824
rect 15084 9764 15088 9820
rect 15088 9764 15144 9820
rect 15144 9764 15148 9820
rect 15084 9760 15148 9764
rect 21790 9820 21854 9824
rect 21790 9764 21794 9820
rect 21794 9764 21850 9820
rect 21850 9764 21854 9820
rect 21790 9760 21854 9764
rect 21870 9820 21934 9824
rect 21870 9764 21874 9820
rect 21874 9764 21930 9820
rect 21930 9764 21934 9820
rect 21870 9760 21934 9764
rect 21950 9820 22014 9824
rect 21950 9764 21954 9820
rect 21954 9764 22010 9820
rect 22010 9764 22014 9820
rect 21950 9760 22014 9764
rect 22030 9820 22094 9824
rect 22030 9764 22034 9820
rect 22034 9764 22090 9820
rect 22090 9764 22094 9820
rect 22030 9760 22094 9764
rect 28736 9820 28800 9824
rect 28736 9764 28740 9820
rect 28740 9764 28796 9820
rect 28796 9764 28800 9820
rect 28736 9760 28800 9764
rect 28816 9820 28880 9824
rect 28816 9764 28820 9820
rect 28820 9764 28876 9820
rect 28876 9764 28880 9820
rect 28816 9760 28880 9764
rect 28896 9820 28960 9824
rect 28896 9764 28900 9820
rect 28900 9764 28956 9820
rect 28956 9764 28960 9820
rect 28896 9760 28960 9764
rect 28976 9820 29040 9824
rect 28976 9764 28980 9820
rect 28980 9764 29036 9820
rect 29036 9764 29040 9820
rect 28976 9760 29040 9764
rect 4425 9276 4489 9280
rect 4425 9220 4429 9276
rect 4429 9220 4485 9276
rect 4485 9220 4489 9276
rect 4425 9216 4489 9220
rect 4505 9276 4569 9280
rect 4505 9220 4509 9276
rect 4509 9220 4565 9276
rect 4565 9220 4569 9276
rect 4505 9216 4569 9220
rect 4585 9276 4649 9280
rect 4585 9220 4589 9276
rect 4589 9220 4645 9276
rect 4645 9220 4649 9276
rect 4585 9216 4649 9220
rect 4665 9276 4729 9280
rect 4665 9220 4669 9276
rect 4669 9220 4725 9276
rect 4725 9220 4729 9276
rect 4665 9216 4729 9220
rect 11371 9276 11435 9280
rect 11371 9220 11375 9276
rect 11375 9220 11431 9276
rect 11431 9220 11435 9276
rect 11371 9216 11435 9220
rect 11451 9276 11515 9280
rect 11451 9220 11455 9276
rect 11455 9220 11511 9276
rect 11511 9220 11515 9276
rect 11451 9216 11515 9220
rect 11531 9276 11595 9280
rect 11531 9220 11535 9276
rect 11535 9220 11591 9276
rect 11591 9220 11595 9276
rect 11531 9216 11595 9220
rect 11611 9276 11675 9280
rect 11611 9220 11615 9276
rect 11615 9220 11671 9276
rect 11671 9220 11675 9276
rect 11611 9216 11675 9220
rect 18317 9276 18381 9280
rect 18317 9220 18321 9276
rect 18321 9220 18377 9276
rect 18377 9220 18381 9276
rect 18317 9216 18381 9220
rect 18397 9276 18461 9280
rect 18397 9220 18401 9276
rect 18401 9220 18457 9276
rect 18457 9220 18461 9276
rect 18397 9216 18461 9220
rect 18477 9276 18541 9280
rect 18477 9220 18481 9276
rect 18481 9220 18537 9276
rect 18537 9220 18541 9276
rect 18477 9216 18541 9220
rect 18557 9276 18621 9280
rect 18557 9220 18561 9276
rect 18561 9220 18617 9276
rect 18617 9220 18621 9276
rect 18557 9216 18621 9220
rect 25263 9276 25327 9280
rect 25263 9220 25267 9276
rect 25267 9220 25323 9276
rect 25323 9220 25327 9276
rect 25263 9216 25327 9220
rect 25343 9276 25407 9280
rect 25343 9220 25347 9276
rect 25347 9220 25403 9276
rect 25403 9220 25407 9276
rect 25343 9216 25407 9220
rect 25423 9276 25487 9280
rect 25423 9220 25427 9276
rect 25427 9220 25483 9276
rect 25483 9220 25487 9276
rect 25423 9216 25487 9220
rect 25503 9276 25567 9280
rect 25503 9220 25507 9276
rect 25507 9220 25563 9276
rect 25563 9220 25567 9276
rect 25503 9216 25567 9220
rect 5396 9208 5460 9212
rect 5396 9152 5410 9208
rect 5410 9152 5460 9208
rect 5396 9148 5460 9152
rect 7898 8732 7962 8736
rect 7898 8676 7902 8732
rect 7902 8676 7958 8732
rect 7958 8676 7962 8732
rect 7898 8672 7962 8676
rect 7978 8732 8042 8736
rect 7978 8676 7982 8732
rect 7982 8676 8038 8732
rect 8038 8676 8042 8732
rect 7978 8672 8042 8676
rect 8058 8732 8122 8736
rect 8058 8676 8062 8732
rect 8062 8676 8118 8732
rect 8118 8676 8122 8732
rect 8058 8672 8122 8676
rect 8138 8732 8202 8736
rect 8138 8676 8142 8732
rect 8142 8676 8198 8732
rect 8198 8676 8202 8732
rect 8138 8672 8202 8676
rect 14844 8732 14908 8736
rect 14844 8676 14848 8732
rect 14848 8676 14904 8732
rect 14904 8676 14908 8732
rect 14844 8672 14908 8676
rect 14924 8732 14988 8736
rect 14924 8676 14928 8732
rect 14928 8676 14984 8732
rect 14984 8676 14988 8732
rect 14924 8672 14988 8676
rect 15004 8732 15068 8736
rect 15004 8676 15008 8732
rect 15008 8676 15064 8732
rect 15064 8676 15068 8732
rect 15004 8672 15068 8676
rect 15084 8732 15148 8736
rect 15084 8676 15088 8732
rect 15088 8676 15144 8732
rect 15144 8676 15148 8732
rect 15084 8672 15148 8676
rect 21790 8732 21854 8736
rect 21790 8676 21794 8732
rect 21794 8676 21850 8732
rect 21850 8676 21854 8732
rect 21790 8672 21854 8676
rect 21870 8732 21934 8736
rect 21870 8676 21874 8732
rect 21874 8676 21930 8732
rect 21930 8676 21934 8732
rect 21870 8672 21934 8676
rect 21950 8732 22014 8736
rect 21950 8676 21954 8732
rect 21954 8676 22010 8732
rect 22010 8676 22014 8732
rect 21950 8672 22014 8676
rect 22030 8732 22094 8736
rect 22030 8676 22034 8732
rect 22034 8676 22090 8732
rect 22090 8676 22094 8732
rect 22030 8672 22094 8676
rect 28736 8732 28800 8736
rect 28736 8676 28740 8732
rect 28740 8676 28796 8732
rect 28796 8676 28800 8732
rect 28736 8672 28800 8676
rect 28816 8732 28880 8736
rect 28816 8676 28820 8732
rect 28820 8676 28876 8732
rect 28876 8676 28880 8732
rect 28816 8672 28880 8676
rect 28896 8732 28960 8736
rect 28896 8676 28900 8732
rect 28900 8676 28956 8732
rect 28956 8676 28960 8732
rect 28896 8672 28960 8676
rect 28976 8732 29040 8736
rect 28976 8676 28980 8732
rect 28980 8676 29036 8732
rect 29036 8676 29040 8732
rect 28976 8672 29040 8676
rect 4425 8188 4489 8192
rect 4425 8132 4429 8188
rect 4429 8132 4485 8188
rect 4485 8132 4489 8188
rect 4425 8128 4489 8132
rect 4505 8188 4569 8192
rect 4505 8132 4509 8188
rect 4509 8132 4565 8188
rect 4565 8132 4569 8188
rect 4505 8128 4569 8132
rect 4585 8188 4649 8192
rect 4585 8132 4589 8188
rect 4589 8132 4645 8188
rect 4645 8132 4649 8188
rect 4585 8128 4649 8132
rect 4665 8188 4729 8192
rect 4665 8132 4669 8188
rect 4669 8132 4725 8188
rect 4725 8132 4729 8188
rect 4665 8128 4729 8132
rect 11371 8188 11435 8192
rect 11371 8132 11375 8188
rect 11375 8132 11431 8188
rect 11431 8132 11435 8188
rect 11371 8128 11435 8132
rect 11451 8188 11515 8192
rect 11451 8132 11455 8188
rect 11455 8132 11511 8188
rect 11511 8132 11515 8188
rect 11451 8128 11515 8132
rect 11531 8188 11595 8192
rect 11531 8132 11535 8188
rect 11535 8132 11591 8188
rect 11591 8132 11595 8188
rect 11531 8128 11595 8132
rect 11611 8188 11675 8192
rect 11611 8132 11615 8188
rect 11615 8132 11671 8188
rect 11671 8132 11675 8188
rect 11611 8128 11675 8132
rect 18317 8188 18381 8192
rect 18317 8132 18321 8188
rect 18321 8132 18377 8188
rect 18377 8132 18381 8188
rect 18317 8128 18381 8132
rect 18397 8188 18461 8192
rect 18397 8132 18401 8188
rect 18401 8132 18457 8188
rect 18457 8132 18461 8188
rect 18397 8128 18461 8132
rect 18477 8188 18541 8192
rect 18477 8132 18481 8188
rect 18481 8132 18537 8188
rect 18537 8132 18541 8188
rect 18477 8128 18541 8132
rect 18557 8188 18621 8192
rect 18557 8132 18561 8188
rect 18561 8132 18617 8188
rect 18617 8132 18621 8188
rect 18557 8128 18621 8132
rect 25263 8188 25327 8192
rect 25263 8132 25267 8188
rect 25267 8132 25323 8188
rect 25323 8132 25327 8188
rect 25263 8128 25327 8132
rect 25343 8188 25407 8192
rect 25343 8132 25347 8188
rect 25347 8132 25403 8188
rect 25403 8132 25407 8188
rect 25343 8128 25407 8132
rect 25423 8188 25487 8192
rect 25423 8132 25427 8188
rect 25427 8132 25483 8188
rect 25483 8132 25487 8188
rect 25423 8128 25487 8132
rect 25503 8188 25567 8192
rect 25503 8132 25507 8188
rect 25507 8132 25563 8188
rect 25563 8132 25567 8188
rect 25503 8128 25567 8132
rect 7898 7644 7962 7648
rect 7898 7588 7902 7644
rect 7902 7588 7958 7644
rect 7958 7588 7962 7644
rect 7898 7584 7962 7588
rect 7978 7644 8042 7648
rect 7978 7588 7982 7644
rect 7982 7588 8038 7644
rect 8038 7588 8042 7644
rect 7978 7584 8042 7588
rect 8058 7644 8122 7648
rect 8058 7588 8062 7644
rect 8062 7588 8118 7644
rect 8118 7588 8122 7644
rect 8058 7584 8122 7588
rect 8138 7644 8202 7648
rect 8138 7588 8142 7644
rect 8142 7588 8198 7644
rect 8198 7588 8202 7644
rect 8138 7584 8202 7588
rect 14844 7644 14908 7648
rect 14844 7588 14848 7644
rect 14848 7588 14904 7644
rect 14904 7588 14908 7644
rect 14844 7584 14908 7588
rect 14924 7644 14988 7648
rect 14924 7588 14928 7644
rect 14928 7588 14984 7644
rect 14984 7588 14988 7644
rect 14924 7584 14988 7588
rect 15004 7644 15068 7648
rect 15004 7588 15008 7644
rect 15008 7588 15064 7644
rect 15064 7588 15068 7644
rect 15004 7584 15068 7588
rect 15084 7644 15148 7648
rect 15084 7588 15088 7644
rect 15088 7588 15144 7644
rect 15144 7588 15148 7644
rect 15084 7584 15148 7588
rect 21790 7644 21854 7648
rect 21790 7588 21794 7644
rect 21794 7588 21850 7644
rect 21850 7588 21854 7644
rect 21790 7584 21854 7588
rect 21870 7644 21934 7648
rect 21870 7588 21874 7644
rect 21874 7588 21930 7644
rect 21930 7588 21934 7644
rect 21870 7584 21934 7588
rect 21950 7644 22014 7648
rect 21950 7588 21954 7644
rect 21954 7588 22010 7644
rect 22010 7588 22014 7644
rect 21950 7584 22014 7588
rect 22030 7644 22094 7648
rect 22030 7588 22034 7644
rect 22034 7588 22090 7644
rect 22090 7588 22094 7644
rect 22030 7584 22094 7588
rect 28736 7644 28800 7648
rect 28736 7588 28740 7644
rect 28740 7588 28796 7644
rect 28796 7588 28800 7644
rect 28736 7584 28800 7588
rect 28816 7644 28880 7648
rect 28816 7588 28820 7644
rect 28820 7588 28876 7644
rect 28876 7588 28880 7644
rect 28816 7584 28880 7588
rect 28896 7644 28960 7648
rect 28896 7588 28900 7644
rect 28900 7588 28956 7644
rect 28956 7588 28960 7644
rect 28896 7584 28960 7588
rect 28976 7644 29040 7648
rect 28976 7588 28980 7644
rect 28980 7588 29036 7644
rect 29036 7588 29040 7644
rect 28976 7584 29040 7588
rect 4425 7100 4489 7104
rect 4425 7044 4429 7100
rect 4429 7044 4485 7100
rect 4485 7044 4489 7100
rect 4425 7040 4489 7044
rect 4505 7100 4569 7104
rect 4505 7044 4509 7100
rect 4509 7044 4565 7100
rect 4565 7044 4569 7100
rect 4505 7040 4569 7044
rect 4585 7100 4649 7104
rect 4585 7044 4589 7100
rect 4589 7044 4645 7100
rect 4645 7044 4649 7100
rect 4585 7040 4649 7044
rect 4665 7100 4729 7104
rect 4665 7044 4669 7100
rect 4669 7044 4725 7100
rect 4725 7044 4729 7100
rect 4665 7040 4729 7044
rect 11371 7100 11435 7104
rect 11371 7044 11375 7100
rect 11375 7044 11431 7100
rect 11431 7044 11435 7100
rect 11371 7040 11435 7044
rect 11451 7100 11515 7104
rect 11451 7044 11455 7100
rect 11455 7044 11511 7100
rect 11511 7044 11515 7100
rect 11451 7040 11515 7044
rect 11531 7100 11595 7104
rect 11531 7044 11535 7100
rect 11535 7044 11591 7100
rect 11591 7044 11595 7100
rect 11531 7040 11595 7044
rect 11611 7100 11675 7104
rect 11611 7044 11615 7100
rect 11615 7044 11671 7100
rect 11671 7044 11675 7100
rect 11611 7040 11675 7044
rect 18317 7100 18381 7104
rect 18317 7044 18321 7100
rect 18321 7044 18377 7100
rect 18377 7044 18381 7100
rect 18317 7040 18381 7044
rect 18397 7100 18461 7104
rect 18397 7044 18401 7100
rect 18401 7044 18457 7100
rect 18457 7044 18461 7100
rect 18397 7040 18461 7044
rect 18477 7100 18541 7104
rect 18477 7044 18481 7100
rect 18481 7044 18537 7100
rect 18537 7044 18541 7100
rect 18477 7040 18541 7044
rect 18557 7100 18621 7104
rect 18557 7044 18561 7100
rect 18561 7044 18617 7100
rect 18617 7044 18621 7100
rect 18557 7040 18621 7044
rect 25263 7100 25327 7104
rect 25263 7044 25267 7100
rect 25267 7044 25323 7100
rect 25323 7044 25327 7100
rect 25263 7040 25327 7044
rect 25343 7100 25407 7104
rect 25343 7044 25347 7100
rect 25347 7044 25403 7100
rect 25403 7044 25407 7100
rect 25343 7040 25407 7044
rect 25423 7100 25487 7104
rect 25423 7044 25427 7100
rect 25427 7044 25483 7100
rect 25483 7044 25487 7100
rect 25423 7040 25487 7044
rect 25503 7100 25567 7104
rect 25503 7044 25507 7100
rect 25507 7044 25563 7100
rect 25563 7044 25567 7100
rect 25503 7040 25567 7044
rect 7898 6556 7962 6560
rect 7898 6500 7902 6556
rect 7902 6500 7958 6556
rect 7958 6500 7962 6556
rect 7898 6496 7962 6500
rect 7978 6556 8042 6560
rect 7978 6500 7982 6556
rect 7982 6500 8038 6556
rect 8038 6500 8042 6556
rect 7978 6496 8042 6500
rect 8058 6556 8122 6560
rect 8058 6500 8062 6556
rect 8062 6500 8118 6556
rect 8118 6500 8122 6556
rect 8058 6496 8122 6500
rect 8138 6556 8202 6560
rect 8138 6500 8142 6556
rect 8142 6500 8198 6556
rect 8198 6500 8202 6556
rect 8138 6496 8202 6500
rect 14844 6556 14908 6560
rect 14844 6500 14848 6556
rect 14848 6500 14904 6556
rect 14904 6500 14908 6556
rect 14844 6496 14908 6500
rect 14924 6556 14988 6560
rect 14924 6500 14928 6556
rect 14928 6500 14984 6556
rect 14984 6500 14988 6556
rect 14924 6496 14988 6500
rect 15004 6556 15068 6560
rect 15004 6500 15008 6556
rect 15008 6500 15064 6556
rect 15064 6500 15068 6556
rect 15004 6496 15068 6500
rect 15084 6556 15148 6560
rect 15084 6500 15088 6556
rect 15088 6500 15144 6556
rect 15144 6500 15148 6556
rect 15084 6496 15148 6500
rect 21790 6556 21854 6560
rect 21790 6500 21794 6556
rect 21794 6500 21850 6556
rect 21850 6500 21854 6556
rect 21790 6496 21854 6500
rect 21870 6556 21934 6560
rect 21870 6500 21874 6556
rect 21874 6500 21930 6556
rect 21930 6500 21934 6556
rect 21870 6496 21934 6500
rect 21950 6556 22014 6560
rect 21950 6500 21954 6556
rect 21954 6500 22010 6556
rect 22010 6500 22014 6556
rect 21950 6496 22014 6500
rect 22030 6556 22094 6560
rect 22030 6500 22034 6556
rect 22034 6500 22090 6556
rect 22090 6500 22094 6556
rect 22030 6496 22094 6500
rect 28736 6556 28800 6560
rect 28736 6500 28740 6556
rect 28740 6500 28796 6556
rect 28796 6500 28800 6556
rect 28736 6496 28800 6500
rect 28816 6556 28880 6560
rect 28816 6500 28820 6556
rect 28820 6500 28876 6556
rect 28876 6500 28880 6556
rect 28816 6496 28880 6500
rect 28896 6556 28960 6560
rect 28896 6500 28900 6556
rect 28900 6500 28956 6556
rect 28956 6500 28960 6556
rect 28896 6496 28960 6500
rect 28976 6556 29040 6560
rect 28976 6500 28980 6556
rect 28980 6500 29036 6556
rect 29036 6500 29040 6556
rect 28976 6496 29040 6500
rect 5396 6156 5460 6220
rect 4425 6012 4489 6016
rect 4425 5956 4429 6012
rect 4429 5956 4485 6012
rect 4485 5956 4489 6012
rect 4425 5952 4489 5956
rect 4505 6012 4569 6016
rect 4505 5956 4509 6012
rect 4509 5956 4565 6012
rect 4565 5956 4569 6012
rect 4505 5952 4569 5956
rect 4585 6012 4649 6016
rect 4585 5956 4589 6012
rect 4589 5956 4645 6012
rect 4645 5956 4649 6012
rect 4585 5952 4649 5956
rect 4665 6012 4729 6016
rect 4665 5956 4669 6012
rect 4669 5956 4725 6012
rect 4725 5956 4729 6012
rect 4665 5952 4729 5956
rect 11371 6012 11435 6016
rect 11371 5956 11375 6012
rect 11375 5956 11431 6012
rect 11431 5956 11435 6012
rect 11371 5952 11435 5956
rect 11451 6012 11515 6016
rect 11451 5956 11455 6012
rect 11455 5956 11511 6012
rect 11511 5956 11515 6012
rect 11451 5952 11515 5956
rect 11531 6012 11595 6016
rect 11531 5956 11535 6012
rect 11535 5956 11591 6012
rect 11591 5956 11595 6012
rect 11531 5952 11595 5956
rect 11611 6012 11675 6016
rect 11611 5956 11615 6012
rect 11615 5956 11671 6012
rect 11671 5956 11675 6012
rect 11611 5952 11675 5956
rect 18317 6012 18381 6016
rect 18317 5956 18321 6012
rect 18321 5956 18377 6012
rect 18377 5956 18381 6012
rect 18317 5952 18381 5956
rect 18397 6012 18461 6016
rect 18397 5956 18401 6012
rect 18401 5956 18457 6012
rect 18457 5956 18461 6012
rect 18397 5952 18461 5956
rect 18477 6012 18541 6016
rect 18477 5956 18481 6012
rect 18481 5956 18537 6012
rect 18537 5956 18541 6012
rect 18477 5952 18541 5956
rect 18557 6012 18621 6016
rect 18557 5956 18561 6012
rect 18561 5956 18617 6012
rect 18617 5956 18621 6012
rect 18557 5952 18621 5956
rect 25263 6012 25327 6016
rect 25263 5956 25267 6012
rect 25267 5956 25323 6012
rect 25323 5956 25327 6012
rect 25263 5952 25327 5956
rect 25343 6012 25407 6016
rect 25343 5956 25347 6012
rect 25347 5956 25403 6012
rect 25403 5956 25407 6012
rect 25343 5952 25407 5956
rect 25423 6012 25487 6016
rect 25423 5956 25427 6012
rect 25427 5956 25483 6012
rect 25483 5956 25487 6012
rect 25423 5952 25487 5956
rect 25503 6012 25567 6016
rect 25503 5956 25507 6012
rect 25507 5956 25563 6012
rect 25563 5956 25567 6012
rect 25503 5952 25567 5956
rect 7898 5468 7962 5472
rect 7898 5412 7902 5468
rect 7902 5412 7958 5468
rect 7958 5412 7962 5468
rect 7898 5408 7962 5412
rect 7978 5468 8042 5472
rect 7978 5412 7982 5468
rect 7982 5412 8038 5468
rect 8038 5412 8042 5468
rect 7978 5408 8042 5412
rect 8058 5468 8122 5472
rect 8058 5412 8062 5468
rect 8062 5412 8118 5468
rect 8118 5412 8122 5468
rect 8058 5408 8122 5412
rect 8138 5468 8202 5472
rect 8138 5412 8142 5468
rect 8142 5412 8198 5468
rect 8198 5412 8202 5468
rect 8138 5408 8202 5412
rect 14844 5468 14908 5472
rect 14844 5412 14848 5468
rect 14848 5412 14904 5468
rect 14904 5412 14908 5468
rect 14844 5408 14908 5412
rect 14924 5468 14988 5472
rect 14924 5412 14928 5468
rect 14928 5412 14984 5468
rect 14984 5412 14988 5468
rect 14924 5408 14988 5412
rect 15004 5468 15068 5472
rect 15004 5412 15008 5468
rect 15008 5412 15064 5468
rect 15064 5412 15068 5468
rect 15004 5408 15068 5412
rect 15084 5468 15148 5472
rect 15084 5412 15088 5468
rect 15088 5412 15144 5468
rect 15144 5412 15148 5468
rect 15084 5408 15148 5412
rect 21790 5468 21854 5472
rect 21790 5412 21794 5468
rect 21794 5412 21850 5468
rect 21850 5412 21854 5468
rect 21790 5408 21854 5412
rect 21870 5468 21934 5472
rect 21870 5412 21874 5468
rect 21874 5412 21930 5468
rect 21930 5412 21934 5468
rect 21870 5408 21934 5412
rect 21950 5468 22014 5472
rect 21950 5412 21954 5468
rect 21954 5412 22010 5468
rect 22010 5412 22014 5468
rect 21950 5408 22014 5412
rect 22030 5468 22094 5472
rect 22030 5412 22034 5468
rect 22034 5412 22090 5468
rect 22090 5412 22094 5468
rect 22030 5408 22094 5412
rect 28736 5468 28800 5472
rect 28736 5412 28740 5468
rect 28740 5412 28796 5468
rect 28796 5412 28800 5468
rect 28736 5408 28800 5412
rect 28816 5468 28880 5472
rect 28816 5412 28820 5468
rect 28820 5412 28876 5468
rect 28876 5412 28880 5468
rect 28816 5408 28880 5412
rect 28896 5468 28960 5472
rect 28896 5412 28900 5468
rect 28900 5412 28956 5468
rect 28956 5412 28960 5468
rect 28896 5408 28960 5412
rect 28976 5468 29040 5472
rect 28976 5412 28980 5468
rect 28980 5412 29036 5468
rect 29036 5412 29040 5468
rect 28976 5408 29040 5412
rect 4425 4924 4489 4928
rect 4425 4868 4429 4924
rect 4429 4868 4485 4924
rect 4485 4868 4489 4924
rect 4425 4864 4489 4868
rect 4505 4924 4569 4928
rect 4505 4868 4509 4924
rect 4509 4868 4565 4924
rect 4565 4868 4569 4924
rect 4505 4864 4569 4868
rect 4585 4924 4649 4928
rect 4585 4868 4589 4924
rect 4589 4868 4645 4924
rect 4645 4868 4649 4924
rect 4585 4864 4649 4868
rect 4665 4924 4729 4928
rect 4665 4868 4669 4924
rect 4669 4868 4725 4924
rect 4725 4868 4729 4924
rect 4665 4864 4729 4868
rect 11371 4924 11435 4928
rect 11371 4868 11375 4924
rect 11375 4868 11431 4924
rect 11431 4868 11435 4924
rect 11371 4864 11435 4868
rect 11451 4924 11515 4928
rect 11451 4868 11455 4924
rect 11455 4868 11511 4924
rect 11511 4868 11515 4924
rect 11451 4864 11515 4868
rect 11531 4924 11595 4928
rect 11531 4868 11535 4924
rect 11535 4868 11591 4924
rect 11591 4868 11595 4924
rect 11531 4864 11595 4868
rect 11611 4924 11675 4928
rect 11611 4868 11615 4924
rect 11615 4868 11671 4924
rect 11671 4868 11675 4924
rect 11611 4864 11675 4868
rect 18317 4924 18381 4928
rect 18317 4868 18321 4924
rect 18321 4868 18377 4924
rect 18377 4868 18381 4924
rect 18317 4864 18381 4868
rect 18397 4924 18461 4928
rect 18397 4868 18401 4924
rect 18401 4868 18457 4924
rect 18457 4868 18461 4924
rect 18397 4864 18461 4868
rect 18477 4924 18541 4928
rect 18477 4868 18481 4924
rect 18481 4868 18537 4924
rect 18537 4868 18541 4924
rect 18477 4864 18541 4868
rect 18557 4924 18621 4928
rect 18557 4868 18561 4924
rect 18561 4868 18617 4924
rect 18617 4868 18621 4924
rect 18557 4864 18621 4868
rect 25263 4924 25327 4928
rect 25263 4868 25267 4924
rect 25267 4868 25323 4924
rect 25323 4868 25327 4924
rect 25263 4864 25327 4868
rect 25343 4924 25407 4928
rect 25343 4868 25347 4924
rect 25347 4868 25403 4924
rect 25403 4868 25407 4924
rect 25343 4864 25407 4868
rect 25423 4924 25487 4928
rect 25423 4868 25427 4924
rect 25427 4868 25483 4924
rect 25483 4868 25487 4924
rect 25423 4864 25487 4868
rect 25503 4924 25567 4928
rect 25503 4868 25507 4924
rect 25507 4868 25563 4924
rect 25563 4868 25567 4924
rect 25503 4864 25567 4868
rect 7898 4380 7962 4384
rect 7898 4324 7902 4380
rect 7902 4324 7958 4380
rect 7958 4324 7962 4380
rect 7898 4320 7962 4324
rect 7978 4380 8042 4384
rect 7978 4324 7982 4380
rect 7982 4324 8038 4380
rect 8038 4324 8042 4380
rect 7978 4320 8042 4324
rect 8058 4380 8122 4384
rect 8058 4324 8062 4380
rect 8062 4324 8118 4380
rect 8118 4324 8122 4380
rect 8058 4320 8122 4324
rect 8138 4380 8202 4384
rect 8138 4324 8142 4380
rect 8142 4324 8198 4380
rect 8198 4324 8202 4380
rect 8138 4320 8202 4324
rect 14844 4380 14908 4384
rect 14844 4324 14848 4380
rect 14848 4324 14904 4380
rect 14904 4324 14908 4380
rect 14844 4320 14908 4324
rect 14924 4380 14988 4384
rect 14924 4324 14928 4380
rect 14928 4324 14984 4380
rect 14984 4324 14988 4380
rect 14924 4320 14988 4324
rect 15004 4380 15068 4384
rect 15004 4324 15008 4380
rect 15008 4324 15064 4380
rect 15064 4324 15068 4380
rect 15004 4320 15068 4324
rect 15084 4380 15148 4384
rect 15084 4324 15088 4380
rect 15088 4324 15144 4380
rect 15144 4324 15148 4380
rect 15084 4320 15148 4324
rect 21790 4380 21854 4384
rect 21790 4324 21794 4380
rect 21794 4324 21850 4380
rect 21850 4324 21854 4380
rect 21790 4320 21854 4324
rect 21870 4380 21934 4384
rect 21870 4324 21874 4380
rect 21874 4324 21930 4380
rect 21930 4324 21934 4380
rect 21870 4320 21934 4324
rect 21950 4380 22014 4384
rect 21950 4324 21954 4380
rect 21954 4324 22010 4380
rect 22010 4324 22014 4380
rect 21950 4320 22014 4324
rect 22030 4380 22094 4384
rect 22030 4324 22034 4380
rect 22034 4324 22090 4380
rect 22090 4324 22094 4380
rect 22030 4320 22094 4324
rect 28736 4380 28800 4384
rect 28736 4324 28740 4380
rect 28740 4324 28796 4380
rect 28796 4324 28800 4380
rect 28736 4320 28800 4324
rect 28816 4380 28880 4384
rect 28816 4324 28820 4380
rect 28820 4324 28876 4380
rect 28876 4324 28880 4380
rect 28816 4320 28880 4324
rect 28896 4380 28960 4384
rect 28896 4324 28900 4380
rect 28900 4324 28956 4380
rect 28956 4324 28960 4380
rect 28896 4320 28960 4324
rect 28976 4380 29040 4384
rect 28976 4324 28980 4380
rect 28980 4324 29036 4380
rect 29036 4324 29040 4380
rect 28976 4320 29040 4324
rect 4108 3980 4172 4044
rect 4425 3836 4489 3840
rect 4425 3780 4429 3836
rect 4429 3780 4485 3836
rect 4485 3780 4489 3836
rect 4425 3776 4489 3780
rect 4505 3836 4569 3840
rect 4505 3780 4509 3836
rect 4509 3780 4565 3836
rect 4565 3780 4569 3836
rect 4505 3776 4569 3780
rect 4585 3836 4649 3840
rect 4585 3780 4589 3836
rect 4589 3780 4645 3836
rect 4645 3780 4649 3836
rect 4585 3776 4649 3780
rect 4665 3836 4729 3840
rect 4665 3780 4669 3836
rect 4669 3780 4725 3836
rect 4725 3780 4729 3836
rect 4665 3776 4729 3780
rect 11371 3836 11435 3840
rect 11371 3780 11375 3836
rect 11375 3780 11431 3836
rect 11431 3780 11435 3836
rect 11371 3776 11435 3780
rect 11451 3836 11515 3840
rect 11451 3780 11455 3836
rect 11455 3780 11511 3836
rect 11511 3780 11515 3836
rect 11451 3776 11515 3780
rect 11531 3836 11595 3840
rect 11531 3780 11535 3836
rect 11535 3780 11591 3836
rect 11591 3780 11595 3836
rect 11531 3776 11595 3780
rect 11611 3836 11675 3840
rect 11611 3780 11615 3836
rect 11615 3780 11671 3836
rect 11671 3780 11675 3836
rect 11611 3776 11675 3780
rect 18317 3836 18381 3840
rect 18317 3780 18321 3836
rect 18321 3780 18377 3836
rect 18377 3780 18381 3836
rect 18317 3776 18381 3780
rect 18397 3836 18461 3840
rect 18397 3780 18401 3836
rect 18401 3780 18457 3836
rect 18457 3780 18461 3836
rect 18397 3776 18461 3780
rect 18477 3836 18541 3840
rect 18477 3780 18481 3836
rect 18481 3780 18537 3836
rect 18537 3780 18541 3836
rect 18477 3776 18541 3780
rect 18557 3836 18621 3840
rect 18557 3780 18561 3836
rect 18561 3780 18617 3836
rect 18617 3780 18621 3836
rect 18557 3776 18621 3780
rect 25263 3836 25327 3840
rect 25263 3780 25267 3836
rect 25267 3780 25323 3836
rect 25323 3780 25327 3836
rect 25263 3776 25327 3780
rect 25343 3836 25407 3840
rect 25343 3780 25347 3836
rect 25347 3780 25403 3836
rect 25403 3780 25407 3836
rect 25343 3776 25407 3780
rect 25423 3836 25487 3840
rect 25423 3780 25427 3836
rect 25427 3780 25483 3836
rect 25483 3780 25487 3836
rect 25423 3776 25487 3780
rect 25503 3836 25567 3840
rect 25503 3780 25507 3836
rect 25507 3780 25563 3836
rect 25563 3780 25567 3836
rect 25503 3776 25567 3780
rect 7898 3292 7962 3296
rect 7898 3236 7902 3292
rect 7902 3236 7958 3292
rect 7958 3236 7962 3292
rect 7898 3232 7962 3236
rect 7978 3292 8042 3296
rect 7978 3236 7982 3292
rect 7982 3236 8038 3292
rect 8038 3236 8042 3292
rect 7978 3232 8042 3236
rect 8058 3292 8122 3296
rect 8058 3236 8062 3292
rect 8062 3236 8118 3292
rect 8118 3236 8122 3292
rect 8058 3232 8122 3236
rect 8138 3292 8202 3296
rect 8138 3236 8142 3292
rect 8142 3236 8198 3292
rect 8198 3236 8202 3292
rect 8138 3232 8202 3236
rect 14844 3292 14908 3296
rect 14844 3236 14848 3292
rect 14848 3236 14904 3292
rect 14904 3236 14908 3292
rect 14844 3232 14908 3236
rect 14924 3292 14988 3296
rect 14924 3236 14928 3292
rect 14928 3236 14984 3292
rect 14984 3236 14988 3292
rect 14924 3232 14988 3236
rect 15004 3292 15068 3296
rect 15004 3236 15008 3292
rect 15008 3236 15064 3292
rect 15064 3236 15068 3292
rect 15004 3232 15068 3236
rect 15084 3292 15148 3296
rect 15084 3236 15088 3292
rect 15088 3236 15144 3292
rect 15144 3236 15148 3292
rect 15084 3232 15148 3236
rect 21790 3292 21854 3296
rect 21790 3236 21794 3292
rect 21794 3236 21850 3292
rect 21850 3236 21854 3292
rect 21790 3232 21854 3236
rect 21870 3292 21934 3296
rect 21870 3236 21874 3292
rect 21874 3236 21930 3292
rect 21930 3236 21934 3292
rect 21870 3232 21934 3236
rect 21950 3292 22014 3296
rect 21950 3236 21954 3292
rect 21954 3236 22010 3292
rect 22010 3236 22014 3292
rect 21950 3232 22014 3236
rect 22030 3292 22094 3296
rect 22030 3236 22034 3292
rect 22034 3236 22090 3292
rect 22090 3236 22094 3292
rect 22030 3232 22094 3236
rect 28736 3292 28800 3296
rect 28736 3236 28740 3292
rect 28740 3236 28796 3292
rect 28796 3236 28800 3292
rect 28736 3232 28800 3236
rect 28816 3292 28880 3296
rect 28816 3236 28820 3292
rect 28820 3236 28876 3292
rect 28876 3236 28880 3292
rect 28816 3232 28880 3236
rect 28896 3292 28960 3296
rect 28896 3236 28900 3292
rect 28900 3236 28956 3292
rect 28956 3236 28960 3292
rect 28896 3232 28960 3236
rect 28976 3292 29040 3296
rect 28976 3236 28980 3292
rect 28980 3236 29036 3292
rect 29036 3236 29040 3292
rect 28976 3232 29040 3236
rect 4425 2748 4489 2752
rect 4425 2692 4429 2748
rect 4429 2692 4485 2748
rect 4485 2692 4489 2748
rect 4425 2688 4489 2692
rect 4505 2748 4569 2752
rect 4505 2692 4509 2748
rect 4509 2692 4565 2748
rect 4565 2692 4569 2748
rect 4505 2688 4569 2692
rect 4585 2748 4649 2752
rect 4585 2692 4589 2748
rect 4589 2692 4645 2748
rect 4645 2692 4649 2748
rect 4585 2688 4649 2692
rect 4665 2748 4729 2752
rect 4665 2692 4669 2748
rect 4669 2692 4725 2748
rect 4725 2692 4729 2748
rect 4665 2688 4729 2692
rect 11371 2748 11435 2752
rect 11371 2692 11375 2748
rect 11375 2692 11431 2748
rect 11431 2692 11435 2748
rect 11371 2688 11435 2692
rect 11451 2748 11515 2752
rect 11451 2692 11455 2748
rect 11455 2692 11511 2748
rect 11511 2692 11515 2748
rect 11451 2688 11515 2692
rect 11531 2748 11595 2752
rect 11531 2692 11535 2748
rect 11535 2692 11591 2748
rect 11591 2692 11595 2748
rect 11531 2688 11595 2692
rect 11611 2748 11675 2752
rect 11611 2692 11615 2748
rect 11615 2692 11671 2748
rect 11671 2692 11675 2748
rect 11611 2688 11675 2692
rect 18317 2748 18381 2752
rect 18317 2692 18321 2748
rect 18321 2692 18377 2748
rect 18377 2692 18381 2748
rect 18317 2688 18381 2692
rect 18397 2748 18461 2752
rect 18397 2692 18401 2748
rect 18401 2692 18457 2748
rect 18457 2692 18461 2748
rect 18397 2688 18461 2692
rect 18477 2748 18541 2752
rect 18477 2692 18481 2748
rect 18481 2692 18537 2748
rect 18537 2692 18541 2748
rect 18477 2688 18541 2692
rect 18557 2748 18621 2752
rect 18557 2692 18561 2748
rect 18561 2692 18617 2748
rect 18617 2692 18621 2748
rect 18557 2688 18621 2692
rect 25263 2748 25327 2752
rect 25263 2692 25267 2748
rect 25267 2692 25323 2748
rect 25323 2692 25327 2748
rect 25263 2688 25327 2692
rect 25343 2748 25407 2752
rect 25343 2692 25347 2748
rect 25347 2692 25403 2748
rect 25403 2692 25407 2748
rect 25343 2688 25407 2692
rect 25423 2748 25487 2752
rect 25423 2692 25427 2748
rect 25427 2692 25483 2748
rect 25483 2692 25487 2748
rect 25423 2688 25487 2692
rect 25503 2748 25567 2752
rect 25503 2692 25507 2748
rect 25507 2692 25563 2748
rect 25563 2692 25567 2748
rect 25503 2688 25567 2692
rect 7898 2204 7962 2208
rect 7898 2148 7902 2204
rect 7902 2148 7958 2204
rect 7958 2148 7962 2204
rect 7898 2144 7962 2148
rect 7978 2204 8042 2208
rect 7978 2148 7982 2204
rect 7982 2148 8038 2204
rect 8038 2148 8042 2204
rect 7978 2144 8042 2148
rect 8058 2204 8122 2208
rect 8058 2148 8062 2204
rect 8062 2148 8118 2204
rect 8118 2148 8122 2204
rect 8058 2144 8122 2148
rect 8138 2204 8202 2208
rect 8138 2148 8142 2204
rect 8142 2148 8198 2204
rect 8198 2148 8202 2204
rect 8138 2144 8202 2148
rect 14844 2204 14908 2208
rect 14844 2148 14848 2204
rect 14848 2148 14904 2204
rect 14904 2148 14908 2204
rect 14844 2144 14908 2148
rect 14924 2204 14988 2208
rect 14924 2148 14928 2204
rect 14928 2148 14984 2204
rect 14984 2148 14988 2204
rect 14924 2144 14988 2148
rect 15004 2204 15068 2208
rect 15004 2148 15008 2204
rect 15008 2148 15064 2204
rect 15064 2148 15068 2204
rect 15004 2144 15068 2148
rect 15084 2204 15148 2208
rect 15084 2148 15088 2204
rect 15088 2148 15144 2204
rect 15144 2148 15148 2204
rect 15084 2144 15148 2148
rect 21790 2204 21854 2208
rect 21790 2148 21794 2204
rect 21794 2148 21850 2204
rect 21850 2148 21854 2204
rect 21790 2144 21854 2148
rect 21870 2204 21934 2208
rect 21870 2148 21874 2204
rect 21874 2148 21930 2204
rect 21930 2148 21934 2204
rect 21870 2144 21934 2148
rect 21950 2204 22014 2208
rect 21950 2148 21954 2204
rect 21954 2148 22010 2204
rect 22010 2148 22014 2204
rect 21950 2144 22014 2148
rect 22030 2204 22094 2208
rect 22030 2148 22034 2204
rect 22034 2148 22090 2204
rect 22090 2148 22094 2204
rect 22030 2144 22094 2148
rect 28736 2204 28800 2208
rect 28736 2148 28740 2204
rect 28740 2148 28796 2204
rect 28796 2148 28800 2204
rect 28736 2144 28800 2148
rect 28816 2204 28880 2208
rect 28816 2148 28820 2204
rect 28820 2148 28876 2204
rect 28876 2148 28880 2204
rect 28816 2144 28880 2148
rect 28896 2204 28960 2208
rect 28896 2148 28900 2204
rect 28900 2148 28956 2204
rect 28956 2148 28960 2204
rect 28896 2144 28960 2148
rect 28976 2204 29040 2208
rect 28976 2148 28980 2204
rect 28980 2148 29036 2204
rect 29036 2148 29040 2204
rect 28976 2144 29040 2148
<< metal4 >>
rect 4417 27776 4737 27792
rect 4417 27712 4425 27776
rect 4489 27712 4505 27776
rect 4569 27712 4585 27776
rect 4649 27712 4665 27776
rect 4729 27712 4737 27776
rect 4417 26688 4737 27712
rect 4417 26624 4425 26688
rect 4489 26624 4505 26688
rect 4569 26624 4585 26688
rect 4649 26624 4665 26688
rect 4729 26624 4737 26688
rect 4417 25600 4737 26624
rect 4417 25536 4425 25600
rect 4489 25536 4505 25600
rect 4569 25536 4585 25600
rect 4649 25536 4665 25600
rect 4729 25536 4737 25600
rect 4417 24512 4737 25536
rect 4417 24448 4425 24512
rect 4489 24448 4505 24512
rect 4569 24448 4585 24512
rect 4649 24448 4665 24512
rect 4729 24448 4737 24512
rect 4417 23424 4737 24448
rect 4417 23360 4425 23424
rect 4489 23360 4505 23424
rect 4569 23360 4585 23424
rect 4649 23360 4665 23424
rect 4729 23360 4737 23424
rect 4417 22336 4737 23360
rect 4417 22272 4425 22336
rect 4489 22272 4505 22336
rect 4569 22272 4585 22336
rect 4649 22272 4665 22336
rect 4729 22272 4737 22336
rect 4417 21248 4737 22272
rect 4417 21184 4425 21248
rect 4489 21184 4505 21248
rect 4569 21184 4585 21248
rect 4649 21184 4665 21248
rect 4729 21184 4737 21248
rect 4417 20160 4737 21184
rect 4417 20096 4425 20160
rect 4489 20096 4505 20160
rect 4569 20096 4585 20160
rect 4649 20096 4665 20160
rect 4729 20096 4737 20160
rect 4417 19072 4737 20096
rect 4417 19008 4425 19072
rect 4489 19008 4505 19072
rect 4569 19008 4585 19072
rect 4649 19008 4665 19072
rect 4729 19008 4737 19072
rect 4417 17984 4737 19008
rect 4417 17920 4425 17984
rect 4489 17920 4505 17984
rect 4569 17920 4585 17984
rect 4649 17920 4665 17984
rect 4729 17920 4737 17984
rect 4417 16896 4737 17920
rect 4417 16832 4425 16896
rect 4489 16832 4505 16896
rect 4569 16832 4585 16896
rect 4649 16832 4665 16896
rect 4729 16832 4737 16896
rect 4417 15808 4737 16832
rect 4417 15744 4425 15808
rect 4489 15744 4505 15808
rect 4569 15744 4585 15808
rect 4649 15744 4665 15808
rect 4729 15744 4737 15808
rect 4107 15332 4173 15333
rect 4107 15268 4108 15332
rect 4172 15268 4173 15332
rect 4107 15267 4173 15268
rect 4110 4045 4170 15267
rect 4417 14720 4737 15744
rect 4417 14656 4425 14720
rect 4489 14656 4505 14720
rect 4569 14656 4585 14720
rect 4649 14656 4665 14720
rect 4729 14656 4737 14720
rect 4417 13632 4737 14656
rect 4417 13568 4425 13632
rect 4489 13568 4505 13632
rect 4569 13568 4585 13632
rect 4649 13568 4665 13632
rect 4729 13568 4737 13632
rect 4417 12544 4737 13568
rect 4417 12480 4425 12544
rect 4489 12480 4505 12544
rect 4569 12480 4585 12544
rect 4649 12480 4665 12544
rect 4729 12480 4737 12544
rect 4417 11456 4737 12480
rect 4417 11392 4425 11456
rect 4489 11392 4505 11456
rect 4569 11392 4585 11456
rect 4649 11392 4665 11456
rect 4729 11392 4737 11456
rect 4417 10368 4737 11392
rect 4417 10304 4425 10368
rect 4489 10304 4505 10368
rect 4569 10304 4585 10368
rect 4649 10304 4665 10368
rect 4729 10304 4737 10368
rect 4417 9280 4737 10304
rect 4417 9216 4425 9280
rect 4489 9216 4505 9280
rect 4569 9216 4585 9280
rect 4649 9216 4665 9280
rect 4729 9216 4737 9280
rect 4417 8192 4737 9216
rect 7890 27232 8210 27792
rect 7890 27168 7898 27232
rect 7962 27168 7978 27232
rect 8042 27168 8058 27232
rect 8122 27168 8138 27232
rect 8202 27168 8210 27232
rect 7890 26144 8210 27168
rect 7890 26080 7898 26144
rect 7962 26080 7978 26144
rect 8042 26080 8058 26144
rect 8122 26080 8138 26144
rect 8202 26080 8210 26144
rect 7890 25056 8210 26080
rect 7890 24992 7898 25056
rect 7962 24992 7978 25056
rect 8042 24992 8058 25056
rect 8122 24992 8138 25056
rect 8202 24992 8210 25056
rect 7890 23968 8210 24992
rect 7890 23904 7898 23968
rect 7962 23904 7978 23968
rect 8042 23904 8058 23968
rect 8122 23904 8138 23968
rect 8202 23904 8210 23968
rect 7890 22880 8210 23904
rect 7890 22816 7898 22880
rect 7962 22816 7978 22880
rect 8042 22816 8058 22880
rect 8122 22816 8138 22880
rect 8202 22816 8210 22880
rect 7890 21792 8210 22816
rect 7890 21728 7898 21792
rect 7962 21728 7978 21792
rect 8042 21728 8058 21792
rect 8122 21728 8138 21792
rect 8202 21728 8210 21792
rect 7890 20704 8210 21728
rect 7890 20640 7898 20704
rect 7962 20640 7978 20704
rect 8042 20640 8058 20704
rect 8122 20640 8138 20704
rect 8202 20640 8210 20704
rect 7890 19616 8210 20640
rect 7890 19552 7898 19616
rect 7962 19552 7978 19616
rect 8042 19552 8058 19616
rect 8122 19552 8138 19616
rect 8202 19552 8210 19616
rect 7890 18528 8210 19552
rect 11363 27776 11683 27792
rect 11363 27712 11371 27776
rect 11435 27712 11451 27776
rect 11515 27712 11531 27776
rect 11595 27712 11611 27776
rect 11675 27712 11683 27776
rect 11363 26688 11683 27712
rect 11363 26624 11371 26688
rect 11435 26624 11451 26688
rect 11515 26624 11531 26688
rect 11595 26624 11611 26688
rect 11675 26624 11683 26688
rect 11363 25600 11683 26624
rect 11363 25536 11371 25600
rect 11435 25536 11451 25600
rect 11515 25536 11531 25600
rect 11595 25536 11611 25600
rect 11675 25536 11683 25600
rect 11363 24512 11683 25536
rect 11363 24448 11371 24512
rect 11435 24448 11451 24512
rect 11515 24448 11531 24512
rect 11595 24448 11611 24512
rect 11675 24448 11683 24512
rect 11363 23424 11683 24448
rect 11363 23360 11371 23424
rect 11435 23360 11451 23424
rect 11515 23360 11531 23424
rect 11595 23360 11611 23424
rect 11675 23360 11683 23424
rect 11363 22336 11683 23360
rect 11363 22272 11371 22336
rect 11435 22272 11451 22336
rect 11515 22272 11531 22336
rect 11595 22272 11611 22336
rect 11675 22272 11683 22336
rect 11363 21248 11683 22272
rect 11363 21184 11371 21248
rect 11435 21184 11451 21248
rect 11515 21184 11531 21248
rect 11595 21184 11611 21248
rect 11675 21184 11683 21248
rect 11363 20160 11683 21184
rect 11363 20096 11371 20160
rect 11435 20096 11451 20160
rect 11515 20096 11531 20160
rect 11595 20096 11611 20160
rect 11675 20096 11683 20160
rect 11363 19072 11683 20096
rect 11363 19008 11371 19072
rect 11435 19008 11451 19072
rect 11515 19008 11531 19072
rect 11595 19008 11611 19072
rect 11675 19008 11683 19072
rect 8339 18868 8405 18869
rect 8339 18804 8340 18868
rect 8404 18804 8405 18868
rect 8339 18803 8405 18804
rect 7890 18464 7898 18528
rect 7962 18464 7978 18528
rect 8042 18464 8058 18528
rect 8122 18464 8138 18528
rect 8202 18464 8210 18528
rect 7890 17440 8210 18464
rect 7890 17376 7898 17440
rect 7962 17376 7978 17440
rect 8042 17376 8058 17440
rect 8122 17376 8138 17440
rect 8202 17376 8210 17440
rect 7890 16352 8210 17376
rect 7890 16288 7898 16352
rect 7962 16288 7978 16352
rect 8042 16288 8058 16352
rect 8122 16288 8138 16352
rect 8202 16288 8210 16352
rect 7890 15264 8210 16288
rect 7890 15200 7898 15264
rect 7962 15200 7978 15264
rect 8042 15200 8058 15264
rect 8122 15200 8138 15264
rect 8202 15200 8210 15264
rect 7890 14176 8210 15200
rect 7890 14112 7898 14176
rect 7962 14112 7978 14176
rect 8042 14112 8058 14176
rect 8122 14112 8138 14176
rect 8202 14112 8210 14176
rect 7890 13088 8210 14112
rect 8342 13701 8402 18803
rect 11363 17984 11683 19008
rect 11363 17920 11371 17984
rect 11435 17920 11451 17984
rect 11515 17920 11531 17984
rect 11595 17920 11611 17984
rect 11675 17920 11683 17984
rect 11363 16896 11683 17920
rect 11363 16832 11371 16896
rect 11435 16832 11451 16896
rect 11515 16832 11531 16896
rect 11595 16832 11611 16896
rect 11675 16832 11683 16896
rect 11363 15808 11683 16832
rect 11363 15744 11371 15808
rect 11435 15744 11451 15808
rect 11515 15744 11531 15808
rect 11595 15744 11611 15808
rect 11675 15744 11683 15808
rect 11363 14720 11683 15744
rect 11363 14656 11371 14720
rect 11435 14656 11451 14720
rect 11515 14656 11531 14720
rect 11595 14656 11611 14720
rect 11675 14656 11683 14720
rect 8339 13700 8405 13701
rect 8339 13636 8340 13700
rect 8404 13636 8405 13700
rect 8339 13635 8405 13636
rect 7890 13024 7898 13088
rect 7962 13024 7978 13088
rect 8042 13024 8058 13088
rect 8122 13024 8138 13088
rect 8202 13024 8210 13088
rect 7890 12000 8210 13024
rect 7890 11936 7898 12000
rect 7962 11936 7978 12000
rect 8042 11936 8058 12000
rect 8122 11936 8138 12000
rect 8202 11936 8210 12000
rect 7890 10912 8210 11936
rect 7890 10848 7898 10912
rect 7962 10848 7978 10912
rect 8042 10848 8058 10912
rect 8122 10848 8138 10912
rect 8202 10848 8210 10912
rect 7890 9824 8210 10848
rect 7890 9760 7898 9824
rect 7962 9760 7978 9824
rect 8042 9760 8058 9824
rect 8122 9760 8138 9824
rect 8202 9760 8210 9824
rect 5395 9212 5461 9213
rect 5395 9148 5396 9212
rect 5460 9148 5461 9212
rect 5395 9147 5461 9148
rect 4417 8128 4425 8192
rect 4489 8128 4505 8192
rect 4569 8128 4585 8192
rect 4649 8128 4665 8192
rect 4729 8128 4737 8192
rect 4417 7104 4737 8128
rect 4417 7040 4425 7104
rect 4489 7040 4505 7104
rect 4569 7040 4585 7104
rect 4649 7040 4665 7104
rect 4729 7040 4737 7104
rect 4417 6016 4737 7040
rect 5398 6221 5458 9147
rect 7890 8736 8210 9760
rect 7890 8672 7898 8736
rect 7962 8672 7978 8736
rect 8042 8672 8058 8736
rect 8122 8672 8138 8736
rect 8202 8672 8210 8736
rect 7890 7648 8210 8672
rect 7890 7584 7898 7648
rect 7962 7584 7978 7648
rect 8042 7584 8058 7648
rect 8122 7584 8138 7648
rect 8202 7584 8210 7648
rect 7890 6560 8210 7584
rect 7890 6496 7898 6560
rect 7962 6496 7978 6560
rect 8042 6496 8058 6560
rect 8122 6496 8138 6560
rect 8202 6496 8210 6560
rect 5395 6220 5461 6221
rect 5395 6156 5396 6220
rect 5460 6156 5461 6220
rect 5395 6155 5461 6156
rect 4417 5952 4425 6016
rect 4489 5952 4505 6016
rect 4569 5952 4585 6016
rect 4649 5952 4665 6016
rect 4729 5952 4737 6016
rect 4417 4928 4737 5952
rect 4417 4864 4425 4928
rect 4489 4864 4505 4928
rect 4569 4864 4585 4928
rect 4649 4864 4665 4928
rect 4729 4864 4737 4928
rect 4107 4044 4173 4045
rect 4107 3980 4108 4044
rect 4172 3980 4173 4044
rect 4107 3979 4173 3980
rect 4417 3840 4737 4864
rect 4417 3776 4425 3840
rect 4489 3776 4505 3840
rect 4569 3776 4585 3840
rect 4649 3776 4665 3840
rect 4729 3776 4737 3840
rect 4417 2752 4737 3776
rect 4417 2688 4425 2752
rect 4489 2688 4505 2752
rect 4569 2688 4585 2752
rect 4649 2688 4665 2752
rect 4729 2688 4737 2752
rect 4417 2128 4737 2688
rect 7890 5472 8210 6496
rect 7890 5408 7898 5472
rect 7962 5408 7978 5472
rect 8042 5408 8058 5472
rect 8122 5408 8138 5472
rect 8202 5408 8210 5472
rect 7890 4384 8210 5408
rect 7890 4320 7898 4384
rect 7962 4320 7978 4384
rect 8042 4320 8058 4384
rect 8122 4320 8138 4384
rect 8202 4320 8210 4384
rect 7890 3296 8210 4320
rect 7890 3232 7898 3296
rect 7962 3232 7978 3296
rect 8042 3232 8058 3296
rect 8122 3232 8138 3296
rect 8202 3232 8210 3296
rect 7890 2208 8210 3232
rect 7890 2144 7898 2208
rect 7962 2144 7978 2208
rect 8042 2144 8058 2208
rect 8122 2144 8138 2208
rect 8202 2144 8210 2208
rect 7890 2128 8210 2144
rect 11363 13632 11683 14656
rect 11363 13568 11371 13632
rect 11435 13568 11451 13632
rect 11515 13568 11531 13632
rect 11595 13568 11611 13632
rect 11675 13568 11683 13632
rect 11363 12544 11683 13568
rect 11363 12480 11371 12544
rect 11435 12480 11451 12544
rect 11515 12480 11531 12544
rect 11595 12480 11611 12544
rect 11675 12480 11683 12544
rect 11363 11456 11683 12480
rect 11363 11392 11371 11456
rect 11435 11392 11451 11456
rect 11515 11392 11531 11456
rect 11595 11392 11611 11456
rect 11675 11392 11683 11456
rect 11363 10368 11683 11392
rect 11363 10304 11371 10368
rect 11435 10304 11451 10368
rect 11515 10304 11531 10368
rect 11595 10304 11611 10368
rect 11675 10304 11683 10368
rect 11363 9280 11683 10304
rect 11363 9216 11371 9280
rect 11435 9216 11451 9280
rect 11515 9216 11531 9280
rect 11595 9216 11611 9280
rect 11675 9216 11683 9280
rect 11363 8192 11683 9216
rect 11363 8128 11371 8192
rect 11435 8128 11451 8192
rect 11515 8128 11531 8192
rect 11595 8128 11611 8192
rect 11675 8128 11683 8192
rect 11363 7104 11683 8128
rect 11363 7040 11371 7104
rect 11435 7040 11451 7104
rect 11515 7040 11531 7104
rect 11595 7040 11611 7104
rect 11675 7040 11683 7104
rect 11363 6016 11683 7040
rect 11363 5952 11371 6016
rect 11435 5952 11451 6016
rect 11515 5952 11531 6016
rect 11595 5952 11611 6016
rect 11675 5952 11683 6016
rect 11363 4928 11683 5952
rect 11363 4864 11371 4928
rect 11435 4864 11451 4928
rect 11515 4864 11531 4928
rect 11595 4864 11611 4928
rect 11675 4864 11683 4928
rect 11363 3840 11683 4864
rect 11363 3776 11371 3840
rect 11435 3776 11451 3840
rect 11515 3776 11531 3840
rect 11595 3776 11611 3840
rect 11675 3776 11683 3840
rect 11363 2752 11683 3776
rect 11363 2688 11371 2752
rect 11435 2688 11451 2752
rect 11515 2688 11531 2752
rect 11595 2688 11611 2752
rect 11675 2688 11683 2752
rect 11363 2128 11683 2688
rect 14836 27232 15156 27792
rect 14836 27168 14844 27232
rect 14908 27168 14924 27232
rect 14988 27168 15004 27232
rect 15068 27168 15084 27232
rect 15148 27168 15156 27232
rect 14836 26144 15156 27168
rect 14836 26080 14844 26144
rect 14908 26080 14924 26144
rect 14988 26080 15004 26144
rect 15068 26080 15084 26144
rect 15148 26080 15156 26144
rect 14836 25056 15156 26080
rect 14836 24992 14844 25056
rect 14908 24992 14924 25056
rect 14988 24992 15004 25056
rect 15068 24992 15084 25056
rect 15148 24992 15156 25056
rect 14836 23968 15156 24992
rect 14836 23904 14844 23968
rect 14908 23904 14924 23968
rect 14988 23904 15004 23968
rect 15068 23904 15084 23968
rect 15148 23904 15156 23968
rect 14836 22880 15156 23904
rect 14836 22816 14844 22880
rect 14908 22816 14924 22880
rect 14988 22816 15004 22880
rect 15068 22816 15084 22880
rect 15148 22816 15156 22880
rect 14836 21792 15156 22816
rect 14836 21728 14844 21792
rect 14908 21728 14924 21792
rect 14988 21728 15004 21792
rect 15068 21728 15084 21792
rect 15148 21728 15156 21792
rect 14836 20704 15156 21728
rect 14836 20640 14844 20704
rect 14908 20640 14924 20704
rect 14988 20640 15004 20704
rect 15068 20640 15084 20704
rect 15148 20640 15156 20704
rect 14836 19616 15156 20640
rect 14836 19552 14844 19616
rect 14908 19552 14924 19616
rect 14988 19552 15004 19616
rect 15068 19552 15084 19616
rect 15148 19552 15156 19616
rect 14836 18528 15156 19552
rect 14836 18464 14844 18528
rect 14908 18464 14924 18528
rect 14988 18464 15004 18528
rect 15068 18464 15084 18528
rect 15148 18464 15156 18528
rect 14836 17440 15156 18464
rect 14836 17376 14844 17440
rect 14908 17376 14924 17440
rect 14988 17376 15004 17440
rect 15068 17376 15084 17440
rect 15148 17376 15156 17440
rect 14836 16352 15156 17376
rect 14836 16288 14844 16352
rect 14908 16288 14924 16352
rect 14988 16288 15004 16352
rect 15068 16288 15084 16352
rect 15148 16288 15156 16352
rect 14836 15264 15156 16288
rect 14836 15200 14844 15264
rect 14908 15200 14924 15264
rect 14988 15200 15004 15264
rect 15068 15200 15084 15264
rect 15148 15200 15156 15264
rect 14836 14176 15156 15200
rect 14836 14112 14844 14176
rect 14908 14112 14924 14176
rect 14988 14112 15004 14176
rect 15068 14112 15084 14176
rect 15148 14112 15156 14176
rect 14836 13088 15156 14112
rect 14836 13024 14844 13088
rect 14908 13024 14924 13088
rect 14988 13024 15004 13088
rect 15068 13024 15084 13088
rect 15148 13024 15156 13088
rect 14836 12000 15156 13024
rect 14836 11936 14844 12000
rect 14908 11936 14924 12000
rect 14988 11936 15004 12000
rect 15068 11936 15084 12000
rect 15148 11936 15156 12000
rect 14836 10912 15156 11936
rect 14836 10848 14844 10912
rect 14908 10848 14924 10912
rect 14988 10848 15004 10912
rect 15068 10848 15084 10912
rect 15148 10848 15156 10912
rect 14836 9824 15156 10848
rect 14836 9760 14844 9824
rect 14908 9760 14924 9824
rect 14988 9760 15004 9824
rect 15068 9760 15084 9824
rect 15148 9760 15156 9824
rect 14836 8736 15156 9760
rect 14836 8672 14844 8736
rect 14908 8672 14924 8736
rect 14988 8672 15004 8736
rect 15068 8672 15084 8736
rect 15148 8672 15156 8736
rect 14836 7648 15156 8672
rect 14836 7584 14844 7648
rect 14908 7584 14924 7648
rect 14988 7584 15004 7648
rect 15068 7584 15084 7648
rect 15148 7584 15156 7648
rect 14836 6560 15156 7584
rect 14836 6496 14844 6560
rect 14908 6496 14924 6560
rect 14988 6496 15004 6560
rect 15068 6496 15084 6560
rect 15148 6496 15156 6560
rect 14836 5472 15156 6496
rect 14836 5408 14844 5472
rect 14908 5408 14924 5472
rect 14988 5408 15004 5472
rect 15068 5408 15084 5472
rect 15148 5408 15156 5472
rect 14836 4384 15156 5408
rect 14836 4320 14844 4384
rect 14908 4320 14924 4384
rect 14988 4320 15004 4384
rect 15068 4320 15084 4384
rect 15148 4320 15156 4384
rect 14836 3296 15156 4320
rect 14836 3232 14844 3296
rect 14908 3232 14924 3296
rect 14988 3232 15004 3296
rect 15068 3232 15084 3296
rect 15148 3232 15156 3296
rect 14836 2208 15156 3232
rect 14836 2144 14844 2208
rect 14908 2144 14924 2208
rect 14988 2144 15004 2208
rect 15068 2144 15084 2208
rect 15148 2144 15156 2208
rect 14836 2128 15156 2144
rect 18309 27776 18629 27792
rect 18309 27712 18317 27776
rect 18381 27712 18397 27776
rect 18461 27712 18477 27776
rect 18541 27712 18557 27776
rect 18621 27712 18629 27776
rect 18309 26688 18629 27712
rect 18309 26624 18317 26688
rect 18381 26624 18397 26688
rect 18461 26624 18477 26688
rect 18541 26624 18557 26688
rect 18621 26624 18629 26688
rect 18309 25600 18629 26624
rect 18309 25536 18317 25600
rect 18381 25536 18397 25600
rect 18461 25536 18477 25600
rect 18541 25536 18557 25600
rect 18621 25536 18629 25600
rect 18309 24512 18629 25536
rect 18309 24448 18317 24512
rect 18381 24448 18397 24512
rect 18461 24448 18477 24512
rect 18541 24448 18557 24512
rect 18621 24448 18629 24512
rect 18309 23424 18629 24448
rect 18309 23360 18317 23424
rect 18381 23360 18397 23424
rect 18461 23360 18477 23424
rect 18541 23360 18557 23424
rect 18621 23360 18629 23424
rect 18309 22336 18629 23360
rect 18309 22272 18317 22336
rect 18381 22272 18397 22336
rect 18461 22272 18477 22336
rect 18541 22272 18557 22336
rect 18621 22272 18629 22336
rect 18309 21248 18629 22272
rect 18309 21184 18317 21248
rect 18381 21184 18397 21248
rect 18461 21184 18477 21248
rect 18541 21184 18557 21248
rect 18621 21184 18629 21248
rect 18309 20160 18629 21184
rect 18309 20096 18317 20160
rect 18381 20096 18397 20160
rect 18461 20096 18477 20160
rect 18541 20096 18557 20160
rect 18621 20096 18629 20160
rect 18309 19072 18629 20096
rect 18309 19008 18317 19072
rect 18381 19008 18397 19072
rect 18461 19008 18477 19072
rect 18541 19008 18557 19072
rect 18621 19008 18629 19072
rect 18309 17984 18629 19008
rect 18309 17920 18317 17984
rect 18381 17920 18397 17984
rect 18461 17920 18477 17984
rect 18541 17920 18557 17984
rect 18621 17920 18629 17984
rect 18309 16896 18629 17920
rect 18309 16832 18317 16896
rect 18381 16832 18397 16896
rect 18461 16832 18477 16896
rect 18541 16832 18557 16896
rect 18621 16832 18629 16896
rect 18309 15808 18629 16832
rect 18309 15744 18317 15808
rect 18381 15744 18397 15808
rect 18461 15744 18477 15808
rect 18541 15744 18557 15808
rect 18621 15744 18629 15808
rect 18309 14720 18629 15744
rect 18309 14656 18317 14720
rect 18381 14656 18397 14720
rect 18461 14656 18477 14720
rect 18541 14656 18557 14720
rect 18621 14656 18629 14720
rect 18309 13632 18629 14656
rect 18309 13568 18317 13632
rect 18381 13568 18397 13632
rect 18461 13568 18477 13632
rect 18541 13568 18557 13632
rect 18621 13568 18629 13632
rect 18309 12544 18629 13568
rect 18309 12480 18317 12544
rect 18381 12480 18397 12544
rect 18461 12480 18477 12544
rect 18541 12480 18557 12544
rect 18621 12480 18629 12544
rect 18309 11456 18629 12480
rect 18309 11392 18317 11456
rect 18381 11392 18397 11456
rect 18461 11392 18477 11456
rect 18541 11392 18557 11456
rect 18621 11392 18629 11456
rect 18309 10368 18629 11392
rect 18309 10304 18317 10368
rect 18381 10304 18397 10368
rect 18461 10304 18477 10368
rect 18541 10304 18557 10368
rect 18621 10304 18629 10368
rect 18309 9280 18629 10304
rect 18309 9216 18317 9280
rect 18381 9216 18397 9280
rect 18461 9216 18477 9280
rect 18541 9216 18557 9280
rect 18621 9216 18629 9280
rect 18309 8192 18629 9216
rect 18309 8128 18317 8192
rect 18381 8128 18397 8192
rect 18461 8128 18477 8192
rect 18541 8128 18557 8192
rect 18621 8128 18629 8192
rect 18309 7104 18629 8128
rect 18309 7040 18317 7104
rect 18381 7040 18397 7104
rect 18461 7040 18477 7104
rect 18541 7040 18557 7104
rect 18621 7040 18629 7104
rect 18309 6016 18629 7040
rect 18309 5952 18317 6016
rect 18381 5952 18397 6016
rect 18461 5952 18477 6016
rect 18541 5952 18557 6016
rect 18621 5952 18629 6016
rect 18309 4928 18629 5952
rect 18309 4864 18317 4928
rect 18381 4864 18397 4928
rect 18461 4864 18477 4928
rect 18541 4864 18557 4928
rect 18621 4864 18629 4928
rect 18309 3840 18629 4864
rect 18309 3776 18317 3840
rect 18381 3776 18397 3840
rect 18461 3776 18477 3840
rect 18541 3776 18557 3840
rect 18621 3776 18629 3840
rect 18309 2752 18629 3776
rect 18309 2688 18317 2752
rect 18381 2688 18397 2752
rect 18461 2688 18477 2752
rect 18541 2688 18557 2752
rect 18621 2688 18629 2752
rect 18309 2128 18629 2688
rect 21782 27232 22102 27792
rect 21782 27168 21790 27232
rect 21854 27168 21870 27232
rect 21934 27168 21950 27232
rect 22014 27168 22030 27232
rect 22094 27168 22102 27232
rect 21782 26144 22102 27168
rect 21782 26080 21790 26144
rect 21854 26080 21870 26144
rect 21934 26080 21950 26144
rect 22014 26080 22030 26144
rect 22094 26080 22102 26144
rect 21782 25056 22102 26080
rect 21782 24992 21790 25056
rect 21854 24992 21870 25056
rect 21934 24992 21950 25056
rect 22014 24992 22030 25056
rect 22094 24992 22102 25056
rect 21782 23968 22102 24992
rect 21782 23904 21790 23968
rect 21854 23904 21870 23968
rect 21934 23904 21950 23968
rect 22014 23904 22030 23968
rect 22094 23904 22102 23968
rect 21782 22880 22102 23904
rect 21782 22816 21790 22880
rect 21854 22816 21870 22880
rect 21934 22816 21950 22880
rect 22014 22816 22030 22880
rect 22094 22816 22102 22880
rect 21782 21792 22102 22816
rect 21782 21728 21790 21792
rect 21854 21728 21870 21792
rect 21934 21728 21950 21792
rect 22014 21728 22030 21792
rect 22094 21728 22102 21792
rect 21782 20704 22102 21728
rect 21782 20640 21790 20704
rect 21854 20640 21870 20704
rect 21934 20640 21950 20704
rect 22014 20640 22030 20704
rect 22094 20640 22102 20704
rect 21782 19616 22102 20640
rect 21782 19552 21790 19616
rect 21854 19552 21870 19616
rect 21934 19552 21950 19616
rect 22014 19552 22030 19616
rect 22094 19552 22102 19616
rect 21782 18528 22102 19552
rect 21782 18464 21790 18528
rect 21854 18464 21870 18528
rect 21934 18464 21950 18528
rect 22014 18464 22030 18528
rect 22094 18464 22102 18528
rect 21782 17440 22102 18464
rect 21782 17376 21790 17440
rect 21854 17376 21870 17440
rect 21934 17376 21950 17440
rect 22014 17376 22030 17440
rect 22094 17376 22102 17440
rect 21782 16352 22102 17376
rect 21782 16288 21790 16352
rect 21854 16288 21870 16352
rect 21934 16288 21950 16352
rect 22014 16288 22030 16352
rect 22094 16288 22102 16352
rect 21782 15264 22102 16288
rect 21782 15200 21790 15264
rect 21854 15200 21870 15264
rect 21934 15200 21950 15264
rect 22014 15200 22030 15264
rect 22094 15200 22102 15264
rect 21782 14176 22102 15200
rect 21782 14112 21790 14176
rect 21854 14112 21870 14176
rect 21934 14112 21950 14176
rect 22014 14112 22030 14176
rect 22094 14112 22102 14176
rect 21782 13088 22102 14112
rect 21782 13024 21790 13088
rect 21854 13024 21870 13088
rect 21934 13024 21950 13088
rect 22014 13024 22030 13088
rect 22094 13024 22102 13088
rect 21782 12000 22102 13024
rect 21782 11936 21790 12000
rect 21854 11936 21870 12000
rect 21934 11936 21950 12000
rect 22014 11936 22030 12000
rect 22094 11936 22102 12000
rect 21782 10912 22102 11936
rect 21782 10848 21790 10912
rect 21854 10848 21870 10912
rect 21934 10848 21950 10912
rect 22014 10848 22030 10912
rect 22094 10848 22102 10912
rect 21782 9824 22102 10848
rect 21782 9760 21790 9824
rect 21854 9760 21870 9824
rect 21934 9760 21950 9824
rect 22014 9760 22030 9824
rect 22094 9760 22102 9824
rect 21782 8736 22102 9760
rect 21782 8672 21790 8736
rect 21854 8672 21870 8736
rect 21934 8672 21950 8736
rect 22014 8672 22030 8736
rect 22094 8672 22102 8736
rect 21782 7648 22102 8672
rect 21782 7584 21790 7648
rect 21854 7584 21870 7648
rect 21934 7584 21950 7648
rect 22014 7584 22030 7648
rect 22094 7584 22102 7648
rect 21782 6560 22102 7584
rect 21782 6496 21790 6560
rect 21854 6496 21870 6560
rect 21934 6496 21950 6560
rect 22014 6496 22030 6560
rect 22094 6496 22102 6560
rect 21782 5472 22102 6496
rect 21782 5408 21790 5472
rect 21854 5408 21870 5472
rect 21934 5408 21950 5472
rect 22014 5408 22030 5472
rect 22094 5408 22102 5472
rect 21782 4384 22102 5408
rect 21782 4320 21790 4384
rect 21854 4320 21870 4384
rect 21934 4320 21950 4384
rect 22014 4320 22030 4384
rect 22094 4320 22102 4384
rect 21782 3296 22102 4320
rect 21782 3232 21790 3296
rect 21854 3232 21870 3296
rect 21934 3232 21950 3296
rect 22014 3232 22030 3296
rect 22094 3232 22102 3296
rect 21782 2208 22102 3232
rect 21782 2144 21790 2208
rect 21854 2144 21870 2208
rect 21934 2144 21950 2208
rect 22014 2144 22030 2208
rect 22094 2144 22102 2208
rect 21782 2128 22102 2144
rect 25255 27776 25575 27792
rect 25255 27712 25263 27776
rect 25327 27712 25343 27776
rect 25407 27712 25423 27776
rect 25487 27712 25503 27776
rect 25567 27712 25575 27776
rect 25255 26688 25575 27712
rect 25255 26624 25263 26688
rect 25327 26624 25343 26688
rect 25407 26624 25423 26688
rect 25487 26624 25503 26688
rect 25567 26624 25575 26688
rect 25255 25600 25575 26624
rect 25255 25536 25263 25600
rect 25327 25536 25343 25600
rect 25407 25536 25423 25600
rect 25487 25536 25503 25600
rect 25567 25536 25575 25600
rect 25255 24512 25575 25536
rect 25255 24448 25263 24512
rect 25327 24448 25343 24512
rect 25407 24448 25423 24512
rect 25487 24448 25503 24512
rect 25567 24448 25575 24512
rect 25255 23424 25575 24448
rect 25255 23360 25263 23424
rect 25327 23360 25343 23424
rect 25407 23360 25423 23424
rect 25487 23360 25503 23424
rect 25567 23360 25575 23424
rect 25255 22336 25575 23360
rect 25255 22272 25263 22336
rect 25327 22272 25343 22336
rect 25407 22272 25423 22336
rect 25487 22272 25503 22336
rect 25567 22272 25575 22336
rect 25255 21248 25575 22272
rect 25255 21184 25263 21248
rect 25327 21184 25343 21248
rect 25407 21184 25423 21248
rect 25487 21184 25503 21248
rect 25567 21184 25575 21248
rect 25255 20160 25575 21184
rect 25255 20096 25263 20160
rect 25327 20096 25343 20160
rect 25407 20096 25423 20160
rect 25487 20096 25503 20160
rect 25567 20096 25575 20160
rect 25255 19072 25575 20096
rect 25255 19008 25263 19072
rect 25327 19008 25343 19072
rect 25407 19008 25423 19072
rect 25487 19008 25503 19072
rect 25567 19008 25575 19072
rect 25255 17984 25575 19008
rect 25255 17920 25263 17984
rect 25327 17920 25343 17984
rect 25407 17920 25423 17984
rect 25487 17920 25503 17984
rect 25567 17920 25575 17984
rect 25255 16896 25575 17920
rect 25255 16832 25263 16896
rect 25327 16832 25343 16896
rect 25407 16832 25423 16896
rect 25487 16832 25503 16896
rect 25567 16832 25575 16896
rect 25255 15808 25575 16832
rect 25255 15744 25263 15808
rect 25327 15744 25343 15808
rect 25407 15744 25423 15808
rect 25487 15744 25503 15808
rect 25567 15744 25575 15808
rect 25255 14720 25575 15744
rect 25255 14656 25263 14720
rect 25327 14656 25343 14720
rect 25407 14656 25423 14720
rect 25487 14656 25503 14720
rect 25567 14656 25575 14720
rect 25255 13632 25575 14656
rect 25255 13568 25263 13632
rect 25327 13568 25343 13632
rect 25407 13568 25423 13632
rect 25487 13568 25503 13632
rect 25567 13568 25575 13632
rect 25255 12544 25575 13568
rect 25255 12480 25263 12544
rect 25327 12480 25343 12544
rect 25407 12480 25423 12544
rect 25487 12480 25503 12544
rect 25567 12480 25575 12544
rect 25255 11456 25575 12480
rect 25255 11392 25263 11456
rect 25327 11392 25343 11456
rect 25407 11392 25423 11456
rect 25487 11392 25503 11456
rect 25567 11392 25575 11456
rect 25255 10368 25575 11392
rect 25255 10304 25263 10368
rect 25327 10304 25343 10368
rect 25407 10304 25423 10368
rect 25487 10304 25503 10368
rect 25567 10304 25575 10368
rect 25255 9280 25575 10304
rect 25255 9216 25263 9280
rect 25327 9216 25343 9280
rect 25407 9216 25423 9280
rect 25487 9216 25503 9280
rect 25567 9216 25575 9280
rect 25255 8192 25575 9216
rect 25255 8128 25263 8192
rect 25327 8128 25343 8192
rect 25407 8128 25423 8192
rect 25487 8128 25503 8192
rect 25567 8128 25575 8192
rect 25255 7104 25575 8128
rect 25255 7040 25263 7104
rect 25327 7040 25343 7104
rect 25407 7040 25423 7104
rect 25487 7040 25503 7104
rect 25567 7040 25575 7104
rect 25255 6016 25575 7040
rect 25255 5952 25263 6016
rect 25327 5952 25343 6016
rect 25407 5952 25423 6016
rect 25487 5952 25503 6016
rect 25567 5952 25575 6016
rect 25255 4928 25575 5952
rect 25255 4864 25263 4928
rect 25327 4864 25343 4928
rect 25407 4864 25423 4928
rect 25487 4864 25503 4928
rect 25567 4864 25575 4928
rect 25255 3840 25575 4864
rect 25255 3776 25263 3840
rect 25327 3776 25343 3840
rect 25407 3776 25423 3840
rect 25487 3776 25503 3840
rect 25567 3776 25575 3840
rect 25255 2752 25575 3776
rect 25255 2688 25263 2752
rect 25327 2688 25343 2752
rect 25407 2688 25423 2752
rect 25487 2688 25503 2752
rect 25567 2688 25575 2752
rect 25255 2128 25575 2688
rect 28728 27232 29048 27792
rect 28728 27168 28736 27232
rect 28800 27168 28816 27232
rect 28880 27168 28896 27232
rect 28960 27168 28976 27232
rect 29040 27168 29048 27232
rect 28728 26144 29048 27168
rect 28728 26080 28736 26144
rect 28800 26080 28816 26144
rect 28880 26080 28896 26144
rect 28960 26080 28976 26144
rect 29040 26080 29048 26144
rect 28728 25056 29048 26080
rect 28728 24992 28736 25056
rect 28800 24992 28816 25056
rect 28880 24992 28896 25056
rect 28960 24992 28976 25056
rect 29040 24992 29048 25056
rect 28728 23968 29048 24992
rect 28728 23904 28736 23968
rect 28800 23904 28816 23968
rect 28880 23904 28896 23968
rect 28960 23904 28976 23968
rect 29040 23904 29048 23968
rect 28728 22880 29048 23904
rect 28728 22816 28736 22880
rect 28800 22816 28816 22880
rect 28880 22816 28896 22880
rect 28960 22816 28976 22880
rect 29040 22816 29048 22880
rect 28728 21792 29048 22816
rect 28728 21728 28736 21792
rect 28800 21728 28816 21792
rect 28880 21728 28896 21792
rect 28960 21728 28976 21792
rect 29040 21728 29048 21792
rect 28728 20704 29048 21728
rect 28728 20640 28736 20704
rect 28800 20640 28816 20704
rect 28880 20640 28896 20704
rect 28960 20640 28976 20704
rect 29040 20640 29048 20704
rect 28728 19616 29048 20640
rect 28728 19552 28736 19616
rect 28800 19552 28816 19616
rect 28880 19552 28896 19616
rect 28960 19552 28976 19616
rect 29040 19552 29048 19616
rect 28728 18528 29048 19552
rect 28728 18464 28736 18528
rect 28800 18464 28816 18528
rect 28880 18464 28896 18528
rect 28960 18464 28976 18528
rect 29040 18464 29048 18528
rect 28728 17440 29048 18464
rect 28728 17376 28736 17440
rect 28800 17376 28816 17440
rect 28880 17376 28896 17440
rect 28960 17376 28976 17440
rect 29040 17376 29048 17440
rect 28728 16352 29048 17376
rect 28728 16288 28736 16352
rect 28800 16288 28816 16352
rect 28880 16288 28896 16352
rect 28960 16288 28976 16352
rect 29040 16288 29048 16352
rect 28728 15264 29048 16288
rect 28728 15200 28736 15264
rect 28800 15200 28816 15264
rect 28880 15200 28896 15264
rect 28960 15200 28976 15264
rect 29040 15200 29048 15264
rect 28728 14176 29048 15200
rect 28728 14112 28736 14176
rect 28800 14112 28816 14176
rect 28880 14112 28896 14176
rect 28960 14112 28976 14176
rect 29040 14112 29048 14176
rect 28728 13088 29048 14112
rect 28728 13024 28736 13088
rect 28800 13024 28816 13088
rect 28880 13024 28896 13088
rect 28960 13024 28976 13088
rect 29040 13024 29048 13088
rect 28728 12000 29048 13024
rect 28728 11936 28736 12000
rect 28800 11936 28816 12000
rect 28880 11936 28896 12000
rect 28960 11936 28976 12000
rect 29040 11936 29048 12000
rect 28728 10912 29048 11936
rect 28728 10848 28736 10912
rect 28800 10848 28816 10912
rect 28880 10848 28896 10912
rect 28960 10848 28976 10912
rect 29040 10848 29048 10912
rect 28728 9824 29048 10848
rect 28728 9760 28736 9824
rect 28800 9760 28816 9824
rect 28880 9760 28896 9824
rect 28960 9760 28976 9824
rect 29040 9760 29048 9824
rect 28728 8736 29048 9760
rect 28728 8672 28736 8736
rect 28800 8672 28816 8736
rect 28880 8672 28896 8736
rect 28960 8672 28976 8736
rect 29040 8672 29048 8736
rect 28728 7648 29048 8672
rect 28728 7584 28736 7648
rect 28800 7584 28816 7648
rect 28880 7584 28896 7648
rect 28960 7584 28976 7648
rect 29040 7584 29048 7648
rect 28728 6560 29048 7584
rect 28728 6496 28736 6560
rect 28800 6496 28816 6560
rect 28880 6496 28896 6560
rect 28960 6496 28976 6560
rect 29040 6496 29048 6560
rect 28728 5472 29048 6496
rect 28728 5408 28736 5472
rect 28800 5408 28816 5472
rect 28880 5408 28896 5472
rect 28960 5408 28976 5472
rect 29040 5408 29048 5472
rect 28728 4384 29048 5408
rect 28728 4320 28736 4384
rect 28800 4320 28816 4384
rect 28880 4320 28896 4384
rect 28960 4320 28976 4384
rect 29040 4320 29048 4384
rect 28728 3296 29048 4320
rect 28728 3232 28736 3296
rect 28800 3232 28816 3296
rect 28880 3232 28896 3296
rect 28960 3232 28976 3296
rect 29040 3232 29048 3296
rect 28728 2208 29048 3232
rect 28728 2144 28736 2208
rect 28800 2144 28816 2208
rect 28880 2144 28896 2208
rect 28960 2144 28976 2208
rect 29040 2144 29048 2208
rect 28728 2128 29048 2144
use sky130_fd_sc_hd__inv_2  _095_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 2944 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _096_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 2024 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _097_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 11040 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _098_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 12972 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _099_
timestamp 1688980957
transform 1 0 10580 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _100_
timestamp 1688980957
transform -1 0 13800 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _101_
timestamp 1688980957
transform 1 0 10764 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _102_
timestamp 1688980957
transform -1 0 13064 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _103_
timestamp 1688980957
transform 1 0 10212 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _104_
timestamp 1688980957
transform -1 0 12696 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _105_
timestamp 1688980957
transform -1 0 10856 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _106_
timestamp 1688980957
transform 1 0 9936 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _107_
timestamp 1688980957
transform 1 0 9660 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _108_
timestamp 1688980957
transform -1 0 10580 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _109_
timestamp 1688980957
transform 1 0 9200 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _110_
timestamp 1688980957
transform -1 0 11408 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _111_
timestamp 1688980957
transform 1 0 8372 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _112_
timestamp 1688980957
transform -1 0 11960 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _113_
timestamp 1688980957
transform 1 0 7820 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _114_
timestamp 1688980957
transform -1 0 9752 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _115_
timestamp 1688980957
transform 1 0 8096 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _116_
timestamp 1688980957
transform -1 0 9384 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _117_
timestamp 1688980957
transform 1 0 8924 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _118_
timestamp 1688980957
transform 1 0 8648 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _119_
timestamp 1688980957
transform -1 0 7820 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _120_
timestamp 1688980957
transform 1 0 6808 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _121_
timestamp 1688980957
transform 1 0 8188 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _122_
timestamp 1688980957
transform 1 0 11408 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _123_
timestamp 1688980957
transform 1 0 8924 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _124_
timestamp 1688980957
transform -1 0 13064 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _125_
timestamp 1688980957
transform -1 0 7544 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _126_
timestamp 1688980957
transform 1 0 6532 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _127_
timestamp 1688980957
transform 1 0 6440 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _128_
timestamp 1688980957
transform -1 0 8096 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _129_
timestamp 1688980957
transform 1 0 5244 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _130_
timestamp 1688980957
transform 1 0 6348 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _131_
timestamp 1688980957
transform 1 0 5612 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _132_
timestamp 1688980957
transform -1 0 8004 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _133_
timestamp 1688980957
transform 1 0 4876 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _134_
timestamp 1688980957
transform -1 0 11500 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _135_
timestamp 1688980957
transform 1 0 4968 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _136_
timestamp 1688980957
transform 1 0 5428 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _137_
timestamp 1688980957
transform 1 0 5244 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _138_
timestamp 1688980957
transform 1 0 10304 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _139_
timestamp 1688980957
transform 1 0 4784 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _140_
timestamp 1688980957
transform 1 0 6348 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _141_
timestamp 1688980957
transform 1 0 4876 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _142_
timestamp 1688980957
transform -1 0 9476 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _143_
timestamp 1688980957
transform 1 0 4600 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _144_
timestamp 1688980957
transform 1 0 5428 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _145_
timestamp 1688980957
transform 1 0 4140 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _146_
timestamp 1688980957
transform -1 0 5428 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _147_
timestamp 1688980957
transform 1 0 3864 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _148_
timestamp 1688980957
transform 1 0 8004 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _149_
timestamp 1688980957
transform 1 0 1380 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _150_
timestamp 1688980957
transform 1 0 4416 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _151_
timestamp 1688980957
transform 1 0 4784 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _152_
timestamp 1688980957
transform 1 0 7360 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _153_
timestamp 1688980957
transform 1 0 3220 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _154_
timestamp 1688980957
transform -1 0 6256 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _155_
timestamp 1688980957
transform 1 0 3772 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _156_
timestamp 1688980957
transform 1 0 4508 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _157_
timestamp 1688980957
transform 1 0 1472 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _158_
timestamp 1688980957
transform 1 0 2208 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__and3b_1  _159_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 4416 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _160_
timestamp 1688980957
transform 1 0 9292 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _161_
timestamp 1688980957
transform 1 0 6348 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _162_
timestamp 1688980957
transform 1 0 7360 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _163_
timestamp 1688980957
transform 1 0 8924 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__and2_2  _164_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 7084 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _165_
timestamp 1688980957
transform 1 0 9660 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__and2_2  _166_
timestamp 1688980957
transform 1 0 8924 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _167_
timestamp 1688980957
transform 1 0 9660 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _168_
timestamp 1688980957
transform 1 0 10212 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_2  _169_
timestamp 1688980957
transform 1 0 7360 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _170_
timestamp 1688980957
transform 1 0 12052 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_2  _171_
timestamp 1688980957
transform 1 0 4968 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _172_
timestamp 1688980957
transform 1 0 13984 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__and2_2  _173_
timestamp 1688980957
transform 1 0 10856 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__and2_2  _174_
timestamp 1688980957
transform 1 0 9016 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _175_
timestamp 1688980957
transform 1 0 15732 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__and2_2  _176_
timestamp 1688980957
transform 1 0 9660 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _177_
timestamp 1688980957
transform 1 0 13616 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _178_
timestamp 1688980957
transform 1 0 14076 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__and2_2  _179_
timestamp 1688980957
transform 1 0 9016 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _180_
timestamp 1688980957
transform 1 0 16928 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__and2_2  _181_
timestamp 1688980957
transform 1 0 9752 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _182_
timestamp 1688980957
transform 1 0 16468 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _183_
timestamp 1688980957
transform 1 0 15364 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _184_
timestamp 1688980957
transform 1 0 15088 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _185_
timestamp 1688980957
transform 1 0 16008 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _186_
timestamp 1688980957
transform 1 0 15916 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _187_
timestamp 1688980957
transform 1 0 15732 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _188_
timestamp 1688980957
transform 1 0 15456 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _189_
timestamp 1688980957
transform 1 0 15180 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _190_
timestamp 1688980957
transform 1 0 15548 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _191_
timestamp 1688980957
transform -1 0 1656 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _192_
timestamp 1688980957
transform -1 0 9568 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _193_
timestamp 1688980957
transform -1 0 10028 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _194_
timestamp 1688980957
transform 1 0 4324 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _195_
timestamp 1688980957
transform -1 0 9200 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _196_
timestamp 1688980957
transform -1 0 6624 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _197_
timestamp 1688980957
transform -1 0 8188 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _198_
timestamp 1688980957
transform 1 0 9660 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _199_
timestamp 1688980957
transform -1 0 10212 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _200_
timestamp 1688980957
transform -1 0 11408 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _201_
timestamp 1688980957
transform -1 0 4968 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _202_
timestamp 1688980957
transform -1 0 12880 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _203_
timestamp 1688980957
transform -1 0 7728 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _204_
timestamp 1688980957
transform -1 0 8280 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _205_
timestamp 1688980957
transform -1 0 10580 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _206_
timestamp 1688980957
transform -1 0 7820 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _207_
timestamp 1688980957
transform 1 0 14076 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _208_
timestamp 1688980957
transform 1 0 11684 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _209_
timestamp 1688980957
transform 1 0 6532 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _210_
timestamp 1688980957
transform -1 0 9752 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _211_
timestamp 1688980957
transform 1 0 9752 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _212_
timestamp 1688980957
transform -1 0 11408 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _213_
timestamp 1688980957
transform 1 0 11408 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _214_
timestamp 1688980957
transform -1 0 13892 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _215_
timestamp 1688980957
transform -1 0 13708 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _216_
timestamp 1688980957
transform -1 0 11132 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _217_
timestamp 1688980957
transform -1 0 14812 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _218_
timestamp 1688980957
transform -1 0 14076 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _219_
timestamp 1688980957
transform -1 0 15088 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _220_
timestamp 1688980957
transform -1 0 14352 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_2  _221_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 2392 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _222_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 4140 0 -1 3264
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _223_
timestamp 1688980957
transform 1 0 5244 0 1 3264
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _224_
timestamp 1688980957
transform 1 0 6716 0 1 4352
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _225_
timestamp 1688980957
transform 1 0 3956 0 1 5440
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _226_
timestamp 1688980957
transform 1 0 7728 0 -1 6528
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _227_
timestamp 1688980957
transform 1 0 5060 0 1 6528
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _228_
timestamp 1688980957
transform 1 0 5152 0 1 7616
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _229_
timestamp 1688980957
transform 1 0 8924 0 1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _230_
timestamp 1688980957
transform 1 0 5796 0 1 8704
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _231_
timestamp 1688980957
transform 1 0 9936 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _232_
timestamp 1688980957
transform 1 0 4968 0 1 9792
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _233_
timestamp 1688980957
transform 1 0 11500 0 -1 10880
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _234_
timestamp 1688980957
transform 1 0 6072 0 1 10880
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _235_
timestamp 1688980957
transform 1 0 5704 0 1 13056
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _236_
timestamp 1688980957
transform -1 0 9016 0 -1 11968
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _237_
timestamp 1688980957
transform 1 0 5888 0 1 14144
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _238_
timestamp 1688980957
transform 1 0 11960 0 -1 11968
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _239_
timestamp 1688980957
transform 1 0 11500 0 1 10880
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _240_
timestamp 1688980957
transform 1 0 6072 0 1 16320
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _241_
timestamp 1688980957
transform 1 0 8280 0 -1 13056
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _242_
timestamp 1688980957
transform 1 0 8924 0 1 16320
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _243_
timestamp 1688980957
transform 1 0 8280 0 -1 16320
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _244_
timestamp 1688980957
transform 1 0 11500 0 -1 16320
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _245_
timestamp 1688980957
transform 1 0 11684 0 1 16320
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _246_
timestamp 1688980957
transform 1 0 11408 0 1 17408
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _247_
timestamp 1688980957
transform 1 0 9384 0 1 13056
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _248_
timestamp 1688980957
transform 1 0 11684 0 -1 17408
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _249_
timestamp 1688980957
transform 1 0 11868 0 1 13056
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _250_
timestamp 1688980957
transform 1 0 12052 0 -1 14144
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _251_
timestamp 1688980957
transform 1 0 11868 0 1 14144
box -38 -48 2154 592
use sky130_fd_sc_hd__dfxtp_2  _252_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 3496 0 1 3264
box -38 -48 1602 592
use sky130_fd_sc_hd__diode_2  ANTENNA__095__A dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3128 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__096__D
timestamp 1688980957
transform -1 0 2852 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__098__A0
timestamp 1688980957
transform -1 0 12144 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__100__A0
timestamp 1688980957
transform 1 0 14260 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__102__A0
timestamp 1688980957
transform -1 0 12236 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__104__A0
timestamp 1688980957
transform 1 0 12696 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__106__A0
timestamp 1688980957
transform 1 0 11684 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__108__A0
timestamp 1688980957
transform -1 0 9752 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__110__A0
timestamp 1688980957
transform 1 0 11224 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__112__A0
timestamp 1688980957
transform -1 0 11132 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__114__A0
timestamp 1688980957
transform 1 0 10212 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__114__S
timestamp 1688980957
transform 1 0 8648 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__116__A0
timestamp 1688980957
transform 1 0 9108 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__116__S
timestamp 1688980957
transform -1 0 8556 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__118__A0
timestamp 1688980957
transform 1 0 9476 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__118__S
timestamp 1688980957
transform 1 0 8464 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__120__A0
timestamp 1688980957
transform 1 0 7636 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__122__S
timestamp 1688980957
transform 1 0 11224 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__126__A0
timestamp 1688980957
transform 1 0 7544 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__128__A0
timestamp 1688980957
transform -1 0 5244 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__130__A0
timestamp 1688980957
transform -1 0 5520 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__132__A0
timestamp 1688980957
transform -1 0 8188 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__136__A0
timestamp 1688980957
transform 1 0 4784 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__138__S
timestamp 1688980957
transform 1 0 12052 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__140__A0
timestamp 1688980957
transform -1 0 4876 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__140__S
timestamp 1688980957
transform 1 0 4324 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__142__S
timestamp 1688980957
transform 1 0 11132 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__144__A0
timestamp 1688980957
transform -1 0 4784 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__144__S
timestamp 1688980957
transform 1 0 4232 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__146__A0
timestamp 1688980957
transform -1 0 4140 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__146__S
timestamp 1688980957
transform 1 0 3496 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__148__S
timestamp 1688980957
transform 1 0 10672 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__150__A0
timestamp 1688980957
transform 1 0 10120 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__150__S
timestamp 1688980957
transform 1 0 10856 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__152__S
timestamp 1688980957
transform 1 0 10120 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__154__A0
timestamp 1688980957
transform 1 0 10488 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__154__S
timestamp 1688980957
transform 1 0 10856 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__156__A0
timestamp 1688980957
transform 1 0 11132 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__156__S
timestamp 1688980957
transform 1 0 11684 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__158__S
timestamp 1688980957
transform -1 0 12328 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__161__A
timestamp 1688980957
transform 1 0 11776 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__162__A
timestamp 1688980957
transform 1 0 10764 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__164__A
timestamp 1688980957
transform -1 0 10580 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__166__A
timestamp 1688980957
transform -1 0 9568 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__167__A
timestamp 1688980957
transform -1 0 10580 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__169__A
timestamp 1688980957
transform -1 0 8832 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__171__A
timestamp 1688980957
transform -1 0 4692 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__173__A
timestamp 1688980957
transform -1 0 11776 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__174__A
timestamp 1688980957
transform 1 0 8648 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__175__A
timestamp 1688980957
transform -1 0 15732 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__176__A
timestamp 1688980957
transform 1 0 9752 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__179__A
timestamp 1688980957
transform 1 0 10672 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__180__A
timestamp 1688980957
transform -1 0 17756 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__181__A
timestamp 1688980957
transform -1 0 10488 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__182__A
timestamp 1688980957
transform 1 0 16284 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__183__A
timestamp 1688980957
transform 1 0 15180 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__184__A
timestamp 1688980957
transform -1 0 15088 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__185__A
timestamp 1688980957
transform 1 0 16652 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__186__A
timestamp 1688980957
transform -1 0 15916 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__187__A
timestamp 1688980957
transform -1 0 16560 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__188__A
timestamp 1688980957
transform 1 0 15272 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__189__A
timestamp 1688980957
transform -1 0 15180 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__190__A
timestamp 1688980957
transform 1 0 15364 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__191__A
timestamp 1688980957
transform 1 0 2116 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__192__A
timestamp 1688980957
transform 1 0 9752 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__193__A
timestamp 1688980957
transform 1 0 10120 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__194__A
timestamp 1688980957
transform 1 0 4140 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__195__A
timestamp 1688980957
transform 1 0 9752 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__196__A
timestamp 1688980957
transform 1 0 10488 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__197__A
timestamp 1688980957
transform 1 0 10028 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__198__A
timestamp 1688980957
transform 1 0 10304 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__199__A
timestamp 1688980957
transform 1 0 10764 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__200__A
timestamp 1688980957
transform 1 0 11684 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__217__A
timestamp 1688980957
transform -1 0 15180 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__218__A
timestamp 1688980957
transform 1 0 14260 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__219__A
timestamp 1688980957
transform 1 0 14628 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__220__A
timestamp 1688980957
transform 1 0 14536 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout161_A
timestamp 1688980957
transform 1 0 4784 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout163_A
timestamp 1688980957
transform 1 0 4416 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold94_A
timestamp 1688980957
transform -1 0 3220 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output100_A
timestamp 1688980957
transform 1 0 26680 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output102_A
timestamp 1688980957
transform 1 0 26956 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output103_A
timestamp 1688980957
transform 1 0 26680 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output104_A
timestamp 1688980957
transform 1 0 26680 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output105_A
timestamp 1688980957
transform -1 0 27140 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output108_A
timestamp 1688980957
transform 1 0 26680 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output109_A
timestamp 1688980957
transform 1 0 23736 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output110_A
timestamp 1688980957
transform -1 0 27140 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output111_A
timestamp 1688980957
transform -1 0 27140 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output112_A
timestamp 1688980957
transform 1 0 26680 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output113_A
timestamp 1688980957
transform 1 0 26680 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output114_A
timestamp 1688980957
transform -1 0 27140 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output115_A
timestamp 1688980957
transform -1 0 27140 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output116_A
timestamp 1688980957
transform 1 0 26680 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output117_A
timestamp 1688980957
transform 1 0 26680 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output118_A
timestamp 1688980957
transform -1 0 27140 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output119_A
timestamp 1688980957
transform -1 0 27140 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output120_A
timestamp 1688980957
transform -1 0 25668 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output121_A
timestamp 1688980957
transform 1 0 26680 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output123_A
timestamp 1688980957
transform -1 0 26864 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output125_A
timestamp 1688980957
transform 1 0 26956 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output126_A
timestamp 1688980957
transform 1 0 26680 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output128_A
timestamp 1688980957
transform -1 0 27140 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output129_A
timestamp 1688980957
transform 1 0 20056 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output132_A
timestamp 1688980957
transform -1 0 24288 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output137_A
timestamp 1688980957
transform -1 0 27692 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output160_A
timestamp 1688980957
transform 1 0 26680 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_wb_clk_i dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 7084 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_0__f_wb_clk_i
timestamp 1688980957
transform -1 0 4416 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_1__f_wb_clk_i
timestamp 1688980957
transform 1 0 6072 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_2__f_wb_clk_i
timestamp 1688980957
transform -1 0 7084 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_3__f_wb_clk_i
timestamp 1688980957
transform 1 0 7820 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_8  fanout161 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 8188 0 1 9792
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  fanout162
timestamp 1688980957
transform 1 0 3772 0 1 3264
box -38 -48 1050 592
use sky130_fd_sc_hd__buf_8  fanout163 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  fanout164
timestamp 1688980957
transform 1 0 3036 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_3 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1380 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_133 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 13340 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_139
timestamp 1688980957
transform 1 0 13892 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_141 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_153
timestamp 1688980957
transform 1 0 15180 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_165 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_169 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 16652 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_177
timestamp 1688980957
transform 1 0 17388 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_197
timestamp 1688980957
transform 1 0 19228 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_205
timestamp 1688980957
transform 1 0 19964 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_241
timestamp 1688980957
transform 1 0 23276 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_249
timestamp 1688980957
transform 1 0 24012 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_269
timestamp 1688980957
transform 1 0 25852 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_277
timestamp 1688980957
transform 1 0 26588 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_297 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 28428 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_3
timestamp 1688980957
transform 1 0 1380 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_62
timestamp 1688980957
transform 1 0 6808 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_111
timestamp 1688980957
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_125
timestamp 1688980957
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_137
timestamp 1688980957
transform 1 0 13708 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_149
timestamp 1688980957
transform 1 0 14812 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_161
timestamp 1688980957
transform 1 0 15916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_167
timestamp 1688980957
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_169
timestamp 1688980957
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_181
timestamp 1688980957
transform 1 0 17756 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_189
timestamp 1688980957
transform 1 0 18492 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_273
timestamp 1688980957
transform 1 0 26220 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_279
timestamp 1688980957
transform 1 0 26772 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_297
timestamp 1688980957
transform 1 0 28428 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_3
timestamp 1688980957
transform 1 0 1380 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_7
timestamp 1688980957
transform 1 0 1748 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_26
timestamp 1688980957
transform 1 0 3496 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_73
timestamp 1688980957
transform 1 0 7820 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_82
timestamp 1688980957
transform 1 0 8648 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_93
timestamp 1688980957
transform 1 0 9660 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_114
timestamp 1688980957
transform 1 0 11592 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_118
timestamp 1688980957
transform 1 0 11960 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_122
timestamp 1688980957
transform 1 0 12328 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_134
timestamp 1688980957
transform 1 0 13432 0 1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_141
timestamp 1688980957
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_153
timestamp 1688980957
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_165
timestamp 1688980957
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_177
timestamp 1688980957
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_189
timestamp 1688980957
transform 1 0 18492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_195
timestamp 1688980957
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_197
timestamp 1688980957
transform 1 0 19228 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_205
timestamp 1688980957
transform 1 0 19964 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_238
timestamp 1688980957
transform 1 0 23000 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_285
timestamp 1688980957
transform 1 0 27324 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_289
timestamp 1688980957
transform 1 0 27692 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_295
timestamp 1688980957
transform 1 0 28244 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_35
timestamp 1688980957
transform 1 0 4324 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_46
timestamp 1688980957
transform 1 0 5336 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_103
timestamp 1688980957
transform 1 0 10580 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_107
timestamp 1688980957
transform 1 0 10948 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_111
timestamp 1688980957
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_113
timestamp 1688980957
transform 1 0 11500 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_117
timestamp 1688980957
transform 1 0 11868 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_129
timestamp 1688980957
transform 1 0 12972 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_141
timestamp 1688980957
transform 1 0 14076 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_153
timestamp 1688980957
transform 1 0 15180 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_165
timestamp 1688980957
transform 1 0 16284 0 -1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_169
timestamp 1688980957
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_181
timestamp 1688980957
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_193
timestamp 1688980957
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_205
timestamp 1688980957
transform 1 0 19964 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_225
timestamp 1688980957
transform 1 0 21804 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_279
timestamp 1688980957
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_297
timestamp 1688980957
transform 1 0 28428 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_3
timestamp 1688980957
transform 1 0 1380 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_60
timestamp 1688980957
transform 1 0 6624 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_96
timestamp 1688980957
transform 1 0 9936 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_100
timestamp 1688980957
transform 1 0 10304 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_104
timestamp 1688980957
transform 1 0 10672 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_108
timestamp 1688980957
transform 1 0 11040 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_120
timestamp 1688980957
transform 1 0 12144 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_132
timestamp 1688980957
transform 1 0 13248 0 1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_141
timestamp 1688980957
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_153
timestamp 1688980957
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_165
timestamp 1688980957
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_177
timestamp 1688980957
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_189
timestamp 1688980957
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_195
timestamp 1688980957
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_197
timestamp 1688980957
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_209
timestamp 1688980957
transform 1 0 20332 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_217
timestamp 1688980957
transform 1 0 21068 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_285
timestamp 1688980957
transform 1 0 27324 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_297
timestamp 1688980957
transform 1 0 28428 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_45
timestamp 1688980957
transform 1 0 5244 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_55
timestamp 1688980957
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_92
timestamp 1688980957
transform 1 0 9568 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_96
timestamp 1688980957
transform 1 0 9936 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_100
timestamp 1688980957
transform 1 0 10304 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_104
timestamp 1688980957
transform 1 0 10672 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_108 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 11040 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_113
timestamp 1688980957
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_125
timestamp 1688980957
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_137
timestamp 1688980957
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_149
timestamp 1688980957
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_161
timestamp 1688980957
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_167
timestamp 1688980957
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_169
timestamp 1688980957
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_181
timestamp 1688980957
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_193
timestamp 1688980957
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_205
timestamp 1688980957
transform 1 0 19964 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_217
timestamp 1688980957
transform 1 0 21068 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_223
timestamp 1688980957
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_225
timestamp 1688980957
transform 1 0 21804 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_274
timestamp 1688980957
transform 1 0 26312 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_297
timestamp 1688980957
transform 1 0 28428 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_27
timestamp 1688980957
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_29
timestamp 1688980957
transform 1 0 3772 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_80
timestamp 1688980957
transform 1 0 8464 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_88
timestamp 1688980957
transform 1 0 9200 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_92
timestamp 1688980957
transform 1 0 9568 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_96
timestamp 1688980957
transform 1 0 9936 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_100
timestamp 1688980957
transform 1 0 10304 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_112
timestamp 1688980957
transform 1 0 11408 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_124
timestamp 1688980957
transform 1 0 12512 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_136
timestamp 1688980957
transform 1 0 13616 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_141
timestamp 1688980957
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_153
timestamp 1688980957
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_165
timestamp 1688980957
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_177
timestamp 1688980957
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_189
timestamp 1688980957
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_195
timestamp 1688980957
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_197
timestamp 1688980957
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_209
timestamp 1688980957
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_221
timestamp 1688980957
transform 1 0 21436 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_233
timestamp 1688980957
transform 1 0 22540 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_253
timestamp 1688980957
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_265
timestamp 1688980957
transform 1 0 25484 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_19
timestamp 1688980957
transform 1 0 2852 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_28
timestamp 1688980957
transform 1 0 3680 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_54
timestamp 1688980957
transform 1 0 6072 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_71
timestamp 1688980957
transform 1 0 7636 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_95
timestamp 1688980957
transform 1 0 9844 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_99
timestamp 1688980957
transform 1 0 10212 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_103
timestamp 1688980957
transform 1 0 10580 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_111
timestamp 1688980957
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_113
timestamp 1688980957
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_125
timestamp 1688980957
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_137
timestamp 1688980957
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_149
timestamp 1688980957
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_161
timestamp 1688980957
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_167
timestamp 1688980957
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_169
timestamp 1688980957
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_181
timestamp 1688980957
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_193
timestamp 1688980957
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_205
timestamp 1688980957
transform 1 0 19964 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_217
timestamp 1688980957
transform 1 0 21068 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_223
timestamp 1688980957
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_225
timestamp 1688980957
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_237
timestamp 1688980957
transform 1 0 22908 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_245
timestamp 1688980957
transform 1 0 23644 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_281
timestamp 1688980957
transform 1 0 26956 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_3
timestamp 1688980957
transform 1 0 1380 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_29
timestamp 1688980957
transform 1 0 3772 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_66
timestamp 1688980957
transform 1 0 7176 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_98
timestamp 1688980957
transform 1 0 10120 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_102
timestamp 1688980957
transform 1 0 10488 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_106
timestamp 1688980957
transform 1 0 10856 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_118
timestamp 1688980957
transform 1 0 11960 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_130
timestamp 1688980957
transform 1 0 13064 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_138
timestamp 1688980957
transform 1 0 13800 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_141
timestamp 1688980957
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_153
timestamp 1688980957
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_165
timestamp 1688980957
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_177
timestamp 1688980957
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_189
timestamp 1688980957
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_195
timestamp 1688980957
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_197
timestamp 1688980957
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_209
timestamp 1688980957
transform 1 0 20332 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_221
timestamp 1688980957
transform 1 0 21436 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_233
timestamp 1688980957
transform 1 0 22540 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_245
timestamp 1688980957
transform 1 0 23644 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_251
timestamp 1688980957
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_253
timestamp 1688980957
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_3
timestamp 1688980957
transform 1 0 1380 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_32
timestamp 1688980957
transform 1 0 4048 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_73
timestamp 1688980957
transform 1 0 7820 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_91
timestamp 1688980957
transform 1 0 9476 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_99
timestamp 1688980957
transform 1 0 10212 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_103
timestamp 1688980957
transform 1 0 10580 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_107
timestamp 1688980957
transform 1 0 10948 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_111
timestamp 1688980957
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_113
timestamp 1688980957
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_125
timestamp 1688980957
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_137
timestamp 1688980957
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_149
timestamp 1688980957
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_161
timestamp 1688980957
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_167
timestamp 1688980957
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_169
timestamp 1688980957
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_181
timestamp 1688980957
transform 1 0 17756 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_193
timestamp 1688980957
transform 1 0 18860 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_205
timestamp 1688980957
transform 1 0 19964 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_217
timestamp 1688980957
transform 1 0 21068 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_223
timestamp 1688980957
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_225
timestamp 1688980957
transform 1 0 21804 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_237
timestamp 1688980957
transform 1 0 22908 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_249
timestamp 1688980957
transform 1 0 24012 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_261
timestamp 1688980957
transform 1 0 25116 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_281
timestamp 1688980957
transform 1 0 26956 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_10
timestamp 1688980957
transform 1 0 2024 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_18
timestamp 1688980957
transform 1 0 2760 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_34
timestamp 1688980957
transform 1 0 4232 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_43
timestamp 1688980957
transform 1 0 5060 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_67
timestamp 1688980957
transform 1 0 7268 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_82
timestamp 1688980957
transform 1 0 8648 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_98
timestamp 1688980957
transform 1 0 10120 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_116
timestamp 1688980957
transform 1 0 11776 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_128
timestamp 1688980957
transform 1 0 12880 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_141
timestamp 1688980957
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_153
timestamp 1688980957
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_165
timestamp 1688980957
transform 1 0 16284 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_177
timestamp 1688980957
transform 1 0 17388 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_189
timestamp 1688980957
transform 1 0 18492 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_195
timestamp 1688980957
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_197
timestamp 1688980957
transform 1 0 19228 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_209
timestamp 1688980957
transform 1 0 20332 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_221
timestamp 1688980957
transform 1 0 21436 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_233
timestamp 1688980957
transform 1 0 22540 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_245
timestamp 1688980957
transform 1 0 23644 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_251
timestamp 1688980957
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_253
timestamp 1688980957
transform 1 0 24380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_265
timestamp 1688980957
transform 1 0 25484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_277
timestamp 1688980957
transform 1 0 26588 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_27
timestamp 1688980957
transform 1 0 3588 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_33
timestamp 1688980957
transform 1 0 4140 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_37
timestamp 1688980957
transform 1 0 4508 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_46
timestamp 1688980957
transform 1 0 5336 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_55
timestamp 1688980957
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_121
timestamp 1688980957
transform 1 0 12236 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_133
timestamp 1688980957
transform 1 0 13340 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_145
timestamp 1688980957
transform 1 0 14444 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_157
timestamp 1688980957
transform 1 0 15548 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_165
timestamp 1688980957
transform 1 0 16284 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_169
timestamp 1688980957
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_181
timestamp 1688980957
transform 1 0 17756 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_193
timestamp 1688980957
transform 1 0 18860 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_205
timestamp 1688980957
transform 1 0 19964 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_217
timestamp 1688980957
transform 1 0 21068 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_223
timestamp 1688980957
transform 1 0 21620 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_225
timestamp 1688980957
transform 1 0 21804 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_237
timestamp 1688980957
transform 1 0 22908 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_249
timestamp 1688980957
transform 1 0 24012 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_261
timestamp 1688980957
transform 1 0 25116 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_273
timestamp 1688980957
transform 1 0 26220 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_277
timestamp 1688980957
transform 1 0 26588 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_281
timestamp 1688980957
transform 1 0 26956 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_18
timestamp 1688980957
transform 1 0 2760 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_24
timestamp 1688980957
transform 1 0 3312 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_29
timestamp 1688980957
transform 1 0 3772 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_33
timestamp 1688980957
transform 1 0 4140 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_36
timestamp 1688980957
transform 1 0 4416 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_50
timestamp 1688980957
transform 1 0 5704 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_74
timestamp 1688980957
transform 1 0 7912 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_112
timestamp 1688980957
transform 1 0 11408 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_116
timestamp 1688980957
transform 1 0 11776 0 1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_124
timestamp 1688980957
transform 1 0 12512 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_136
timestamp 1688980957
transform 1 0 13616 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_141
timestamp 1688980957
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_153
timestamp 1688980957
transform 1 0 15180 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_165
timestamp 1688980957
transform 1 0 16284 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_177
timestamp 1688980957
transform 1 0 17388 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_189
timestamp 1688980957
transform 1 0 18492 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_195
timestamp 1688980957
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_197
timestamp 1688980957
transform 1 0 19228 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_209
timestamp 1688980957
transform 1 0 20332 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_221
timestamp 1688980957
transform 1 0 21436 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_233
timestamp 1688980957
transform 1 0 22540 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_245
timestamp 1688980957
transform 1 0 23644 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_251
timestamp 1688980957
transform 1 0 24196 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_253
timestamp 1688980957
transform 1 0 24380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_265
timestamp 1688980957
transform 1 0 25484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_277
timestamp 1688980957
transform 1 0 26588 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_15
timestamp 1688980957
transform 1 0 2484 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_19
timestamp 1688980957
transform 1 0 2852 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_23
timestamp 1688980957
transform 1 0 3220 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_31
timestamp 1688980957
transform 1 0 3956 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_35
timestamp 1688980957
transform 1 0 4324 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_85
timestamp 1688980957
transform 1 0 8924 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_113
timestamp 1688980957
transform 1 0 11500 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_117
timestamp 1688980957
transform 1 0 11868 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_121
timestamp 1688980957
transform 1 0 12236 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_133
timestamp 1688980957
transform 1 0 13340 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_139
timestamp 1688980957
transform 1 0 13892 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_145
timestamp 1688980957
transform 1 0 14444 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_157
timestamp 1688980957
transform 1 0 15548 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_165
timestamp 1688980957
transform 1 0 16284 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_169
timestamp 1688980957
transform 1 0 16652 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_181
timestamp 1688980957
transform 1 0 17756 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_193
timestamp 1688980957
transform 1 0 18860 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_205
timestamp 1688980957
transform 1 0 19964 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_217
timestamp 1688980957
transform 1 0 21068 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_223
timestamp 1688980957
transform 1 0 21620 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_225
timestamp 1688980957
transform 1 0 21804 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_237
timestamp 1688980957
transform 1 0 22908 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_249
timestamp 1688980957
transform 1 0 24012 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_261
timestamp 1688980957
transform 1 0 25116 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_273
timestamp 1688980957
transform 1 0 26220 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_279
timestamp 1688980957
transform 1 0 26772 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_281
timestamp 1688980957
transform 1 0 26956 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_293
timestamp 1688980957
transform 1 0 28060 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_9
timestamp 1688980957
transform 1 0 1932 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_13
timestamp 1688980957
transform 1 0 2300 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_25
timestamp 1688980957
transform 1 0 3404 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_29
timestamp 1688980957
transform 1 0 3772 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_37
timestamp 1688980957
transform 1 0 4508 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_65
timestamp 1688980957
transform 1 0 7084 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_77
timestamp 1688980957
transform 1 0 8188 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_81
timestamp 1688980957
transform 1 0 8556 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_85
timestamp 1688980957
transform 1 0 8924 0 1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_128
timestamp 1688980957
transform 1 0 12880 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_141
timestamp 1688980957
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_153
timestamp 1688980957
transform 1 0 15180 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_165
timestamp 1688980957
transform 1 0 16284 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_177
timestamp 1688980957
transform 1 0 17388 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_189
timestamp 1688980957
transform 1 0 18492 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_195
timestamp 1688980957
transform 1 0 19044 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_197
timestamp 1688980957
transform 1 0 19228 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_209
timestamp 1688980957
transform 1 0 20332 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_221
timestamp 1688980957
transform 1 0 21436 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_233
timestamp 1688980957
transform 1 0 22540 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_245
timestamp 1688980957
transform 1 0 23644 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_251
timestamp 1688980957
transform 1 0 24196 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_253
timestamp 1688980957
transform 1 0 24380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_265
timestamp 1688980957
transform 1 0 25484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_277
timestamp 1688980957
transform 1 0 26588 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_9
timestamp 1688980957
transform 1 0 1932 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_21
timestamp 1688980957
transform 1 0 3036 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_33
timestamp 1688980957
transform 1 0 4140 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_38
timestamp 1688980957
transform 1 0 4600 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_72
timestamp 1688980957
transform 1 0 7728 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_93
timestamp 1688980957
transform 1 0 9660 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_110
timestamp 1688980957
transform 1 0 11224 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_141
timestamp 1688980957
transform 1 0 14076 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_153
timestamp 1688980957
transform 1 0 15180 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_164
timestamp 1688980957
transform 1 0 16192 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_169
timestamp 1688980957
transform 1 0 16652 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_181
timestamp 1688980957
transform 1 0 17756 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_193
timestamp 1688980957
transform 1 0 18860 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_205
timestamp 1688980957
transform 1 0 19964 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_217
timestamp 1688980957
transform 1 0 21068 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_223
timestamp 1688980957
transform 1 0 21620 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_225
timestamp 1688980957
transform 1 0 21804 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_237
timestamp 1688980957
transform 1 0 22908 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_249
timestamp 1688980957
transform 1 0 24012 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_261
timestamp 1688980957
transform 1 0 25116 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_273
timestamp 1688980957
transform 1 0 26220 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_279
timestamp 1688980957
transform 1 0 26772 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_281
timestamp 1688980957
transform 1 0 26956 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_9
timestamp 1688980957
transform 1 0 1932 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_21
timestamp 1688980957
transform 1 0 3036 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_27
timestamp 1688980957
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_29
timestamp 1688980957
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_82
timestamp 1688980957
transform 1 0 8648 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_90
timestamp 1688980957
transform 1 0 9384 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_99
timestamp 1688980957
transform 1 0 10212 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_103
timestamp 1688980957
transform 1 0 10580 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_136
timestamp 1688980957
transform 1 0 13616 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_146
timestamp 1688980957
transform 1 0 14536 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_158
timestamp 1688980957
transform 1 0 15640 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_170
timestamp 1688980957
transform 1 0 16744 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_182
timestamp 1688980957
transform 1 0 17848 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_194
timestamp 1688980957
transform 1 0 18952 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_197
timestamp 1688980957
transform 1 0 19228 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_209
timestamp 1688980957
transform 1 0 20332 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_221
timestamp 1688980957
transform 1 0 21436 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_233
timestamp 1688980957
transform 1 0 22540 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_245
timestamp 1688980957
transform 1 0 23644 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_251
timestamp 1688980957
transform 1 0 24196 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_253
timestamp 1688980957
transform 1 0 24380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_265
timestamp 1688980957
transform 1 0 25484 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_277
timestamp 1688980957
transform 1 0 26588 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_289
timestamp 1688980957
transform 1 0 27692 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_297
timestamp 1688980957
transform 1 0 28428 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_9
timestamp 1688980957
transform 1 0 1932 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_21
timestamp 1688980957
transform 1 0 3036 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_33
timestamp 1688980957
transform 1 0 4140 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_45
timestamp 1688980957
transform 1 0 5244 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_54
timestamp 1688980957
transform 1 0 6072 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_57
timestamp 1688980957
transform 1 0 6348 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_92
timestamp 1688980957
transform 1 0 9568 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_96
timestamp 1688980957
transform 1 0 9936 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_102
timestamp 1688980957
transform 1 0 10488 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_106
timestamp 1688980957
transform 1 0 10856 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_113
timestamp 1688980957
transform 1 0 11500 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_141
timestamp 1688980957
transform 1 0 14076 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_153
timestamp 1688980957
transform 1 0 15180 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_165
timestamp 1688980957
transform 1 0 16284 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_169
timestamp 1688980957
transform 1 0 16652 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_177
timestamp 1688980957
transform 1 0 17388 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_181
timestamp 1688980957
transform 1 0 17756 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_193
timestamp 1688980957
transform 1 0 18860 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_205
timestamp 1688980957
transform 1 0 19964 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_217
timestamp 1688980957
transform 1 0 21068 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_223
timestamp 1688980957
transform 1 0 21620 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_225
timestamp 1688980957
transform 1 0 21804 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_237
timestamp 1688980957
transform 1 0 22908 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_249
timestamp 1688980957
transform 1 0 24012 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_261
timestamp 1688980957
transform 1 0 25116 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_273
timestamp 1688980957
transform 1 0 26220 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_277
timestamp 1688980957
transform 1 0 26588 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_281
timestamp 1688980957
transform 1 0 26956 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_9
timestamp 1688980957
transform 1 0 1932 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_21
timestamp 1688980957
transform 1 0 3036 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_27
timestamp 1688980957
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_29
timestamp 1688980957
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_41
timestamp 1688980957
transform 1 0 4876 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_65
timestamp 1688980957
transform 1 0 7084 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_93
timestamp 1688980957
transform 1 0 9660 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_103
timestamp 1688980957
transform 1 0 10580 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_138
timestamp 1688980957
transform 1 0 13800 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_144
timestamp 1688980957
transform 1 0 14352 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_152
timestamp 1688980957
transform 1 0 15088 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_160
timestamp 1688980957
transform 1 0 15824 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_164
timestamp 1688980957
transform 1 0 16192 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_172
timestamp 1688980957
transform 1 0 16928 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_184
timestamp 1688980957
transform 1 0 18032 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_197
timestamp 1688980957
transform 1 0 19228 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_209
timestamp 1688980957
transform 1 0 20332 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_221
timestamp 1688980957
transform 1 0 21436 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_233
timestamp 1688980957
transform 1 0 22540 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_245
timestamp 1688980957
transform 1 0 23644 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_251
timestamp 1688980957
transform 1 0 24196 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_253
timestamp 1688980957
transform 1 0 24380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_265
timestamp 1688980957
transform 1 0 25484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_277
timestamp 1688980957
transform 1 0 26588 0 1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_9
timestamp 1688980957
transform 1 0 1932 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_21
timestamp 1688980957
transform 1 0 3036 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_33
timestamp 1688980957
transform 1 0 4140 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_45
timestamp 1688980957
transform 1 0 5244 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_109
timestamp 1688980957
transform 1 0 11132 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_113
timestamp 1688980957
transform 1 0 11500 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_141
timestamp 1688980957
transform 1 0 14076 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_145
timestamp 1688980957
transform 1 0 14444 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_149
timestamp 1688980957
transform 1 0 14812 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_157
timestamp 1688980957
transform 1 0 15548 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_166
timestamp 1688980957
transform 1 0 16376 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_169
timestamp 1688980957
transform 1 0 16652 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_181
timestamp 1688980957
transform 1 0 17756 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_193
timestamp 1688980957
transform 1 0 18860 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_205
timestamp 1688980957
transform 1 0 19964 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_217
timestamp 1688980957
transform 1 0 21068 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_223
timestamp 1688980957
transform 1 0 21620 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_225
timestamp 1688980957
transform 1 0 21804 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_237
timestamp 1688980957
transform 1 0 22908 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_249
timestamp 1688980957
transform 1 0 24012 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_261
timestamp 1688980957
transform 1 0 25116 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_273
timestamp 1688980957
transform 1 0 26220 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_279
timestamp 1688980957
transform 1 0 26772 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_281
timestamp 1688980957
transform 1 0 26956 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_293
timestamp 1688980957
transform 1 0 28060 0 -1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_9
timestamp 1688980957
transform 1 0 1932 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_21
timestamp 1688980957
transform 1 0 3036 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_27
timestamp 1688980957
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_29
timestamp 1688980957
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_41
timestamp 1688980957
transform 1 0 4876 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_73
timestamp 1688980957
transform 1 0 7820 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_113
timestamp 1688980957
transform 1 0 11500 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_141
timestamp 1688980957
transform 1 0 14076 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_153
timestamp 1688980957
transform 1 0 15180 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_161
timestamp 1688980957
transform 1 0 15916 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_167
timestamp 1688980957
transform 1 0 16468 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_171
timestamp 1688980957
transform 1 0 16836 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_183
timestamp 1688980957
transform 1 0 17940 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_195
timestamp 1688980957
transform 1 0 19044 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_197
timestamp 1688980957
transform 1 0 19228 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_209
timestamp 1688980957
transform 1 0 20332 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_221
timestamp 1688980957
transform 1 0 21436 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_233
timestamp 1688980957
transform 1 0 22540 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_245
timestamp 1688980957
transform 1 0 23644 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_251
timestamp 1688980957
transform 1 0 24196 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_253
timestamp 1688980957
transform 1 0 24380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_265
timestamp 1688980957
transform 1 0 25484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_277
timestamp 1688980957
transform 1 0 26588 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_9
timestamp 1688980957
transform 1 0 1932 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_21
timestamp 1688980957
transform 1 0 3036 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_33
timestamp 1688980957
transform 1 0 4140 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_45
timestamp 1688980957
transform 1 0 5244 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_53
timestamp 1688980957
transform 1 0 5980 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_57
timestamp 1688980957
transform 1 0 6348 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_68
timestamp 1688980957
transform 1 0 7360 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_72
timestamp 1688980957
transform 1 0 7728 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_77
timestamp 1688980957
transform 1 0 8188 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_94
timestamp 1688980957
transform 1 0 9752 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_110
timestamp 1688980957
transform 1 0 11224 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_113
timestamp 1688980957
transform 1 0 11500 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_117
timestamp 1688980957
transform 1 0 11868 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_142
timestamp 1688980957
transform 1 0 14168 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_146
timestamp 1688980957
transform 1 0 14536 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_149
timestamp 1688980957
transform 1 0 14812 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_158
timestamp 1688980957
transform 1 0 15640 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_164
timestamp 1688980957
transform 1 0 16192 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_169
timestamp 1688980957
transform 1 0 16652 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_181
timestamp 1688980957
transform 1 0 17756 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_193
timestamp 1688980957
transform 1 0 18860 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_205
timestamp 1688980957
transform 1 0 19964 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_217
timestamp 1688980957
transform 1 0 21068 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_223
timestamp 1688980957
transform 1 0 21620 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_225
timestamp 1688980957
transform 1 0 21804 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_237
timestamp 1688980957
transform 1 0 22908 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_249
timestamp 1688980957
transform 1 0 24012 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_261
timestamp 1688980957
transform 1 0 25116 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_273
timestamp 1688980957
transform 1 0 26220 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_277
timestamp 1688980957
transform 1 0 26588 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_281
timestamp 1688980957
transform 1 0 26956 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_9
timestamp 1688980957
transform 1 0 1932 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_21
timestamp 1688980957
transform 1 0 3036 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_27
timestamp 1688980957
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_29
timestamp 1688980957
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_41
timestamp 1688980957
transform 1 0 4876 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_49
timestamp 1688980957
transform 1 0 5612 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_75
timestamp 1688980957
transform 1 0 8004 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_83
timestamp 1688980957
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_85
timestamp 1688980957
transform 1 0 8924 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_93
timestamp 1688980957
transform 1 0 9660 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_113
timestamp 1688980957
transform 1 0 11500 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_152
timestamp 1688980957
transform 1 0 15088 0 1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_162
timestamp 1688980957
transform 1 0 16008 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_174
timestamp 1688980957
transform 1 0 17112 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_186
timestamp 1688980957
transform 1 0 18216 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_194
timestamp 1688980957
transform 1 0 18952 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_197
timestamp 1688980957
transform 1 0 19228 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_209
timestamp 1688980957
transform 1 0 20332 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_221
timestamp 1688980957
transform 1 0 21436 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_233
timestamp 1688980957
transform 1 0 22540 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_245
timestamp 1688980957
transform 1 0 23644 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_251
timestamp 1688980957
transform 1 0 24196 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_253
timestamp 1688980957
transform 1 0 24380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_265
timestamp 1688980957
transform 1 0 25484 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_277
timestamp 1688980957
transform 1 0 26588 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_289
timestamp 1688980957
transform 1 0 27692 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_297
timestamp 1688980957
transform 1 0 28428 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_6
timestamp 1688980957
transform 1 0 1656 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_18
timestamp 1688980957
transform 1 0 2760 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_30
timestamp 1688980957
transform 1 0 3864 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_42
timestamp 1688980957
transform 1 0 4968 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_54
timestamp 1688980957
transform 1 0 6072 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_73
timestamp 1688980957
transform 1 0 7820 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_85
timestamp 1688980957
transform 1 0 8924 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_97
timestamp 1688980957
transform 1 0 10028 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_109
timestamp 1688980957
transform 1 0 11132 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_113
timestamp 1688980957
transform 1 0 11500 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_117
timestamp 1688980957
transform 1 0 11868 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_138
timestamp 1688980957
transform 1 0 13800 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_144
timestamp 1688980957
transform 1 0 14352 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_148
timestamp 1688980957
transform 1 0 14720 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_160
timestamp 1688980957
transform 1 0 15824 0 -1 15232
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_169
timestamp 1688980957
transform 1 0 16652 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_181
timestamp 1688980957
transform 1 0 17756 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_193
timestamp 1688980957
transform 1 0 18860 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_205
timestamp 1688980957
transform 1 0 19964 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_217
timestamp 1688980957
transform 1 0 21068 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_223
timestamp 1688980957
transform 1 0 21620 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_225
timestamp 1688980957
transform 1 0 21804 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_237
timestamp 1688980957
transform 1 0 22908 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_249
timestamp 1688980957
transform 1 0 24012 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_261
timestamp 1688980957
transform 1 0 25116 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_273
timestamp 1688980957
transform 1 0 26220 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_277
timestamp 1688980957
transform 1 0 26588 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_281
timestamp 1688980957
transform 1 0 26956 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_9
timestamp 1688980957
transform 1 0 1932 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_21
timestamp 1688980957
transform 1 0 3036 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_27
timestamp 1688980957
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_29
timestamp 1688980957
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_41
timestamp 1688980957
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_53
timestamp 1688980957
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_65
timestamp 1688980957
transform 1 0 7084 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_73
timestamp 1688980957
transform 1 0 7820 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_81
timestamp 1688980957
transform 1 0 8556 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_97
timestamp 1688980957
transform 1 0 10028 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_101
timestamp 1688980957
transform 1 0 10396 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_137
timestamp 1688980957
transform 1 0 13708 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_141
timestamp 1688980957
transform 1 0 14076 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_145
timestamp 1688980957
transform 1 0 14444 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_157
timestamp 1688980957
transform 1 0 15548 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_169
timestamp 1688980957
transform 1 0 16652 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_181
timestamp 1688980957
transform 1 0 17756 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_193
timestamp 1688980957
transform 1 0 18860 0 1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_197
timestamp 1688980957
transform 1 0 19228 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_209
timestamp 1688980957
transform 1 0 20332 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_221
timestamp 1688980957
transform 1 0 21436 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_233
timestamp 1688980957
transform 1 0 22540 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_245
timestamp 1688980957
transform 1 0 23644 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_251
timestamp 1688980957
transform 1 0 24196 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_253
timestamp 1688980957
transform 1 0 24380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_265
timestamp 1688980957
transform 1 0 25484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_277
timestamp 1688980957
transform 1 0 26588 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_9
timestamp 1688980957
transform 1 0 1932 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_21
timestamp 1688980957
transform 1 0 3036 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_33
timestamp 1688980957
transform 1 0 4140 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_45
timestamp 1688980957
transform 1 0 5244 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_53
timestamp 1688980957
transform 1 0 5980 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_57
timestamp 1688980957
transform 1 0 6348 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_71
timestamp 1688980957
transform 1 0 7636 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_139
timestamp 1688980957
transform 1 0 13892 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_151
timestamp 1688980957
transform 1 0 14996 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_163
timestamp 1688980957
transform 1 0 16100 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_167
timestamp 1688980957
transform 1 0 16468 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_169
timestamp 1688980957
transform 1 0 16652 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_181
timestamp 1688980957
transform 1 0 17756 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_193
timestamp 1688980957
transform 1 0 18860 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_205
timestamp 1688980957
transform 1 0 19964 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_217
timestamp 1688980957
transform 1 0 21068 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_223
timestamp 1688980957
transform 1 0 21620 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_225
timestamp 1688980957
transform 1 0 21804 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_237
timestamp 1688980957
transform 1 0 22908 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_249
timestamp 1688980957
transform 1 0 24012 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_261
timestamp 1688980957
transform 1 0 25116 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_273
timestamp 1688980957
transform 1 0 26220 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_279
timestamp 1688980957
transform 1 0 26772 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_281
timestamp 1688980957
transform 1 0 26956 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_293
timestamp 1688980957
transform 1 0 28060 0 -1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_9
timestamp 1688980957
transform 1 0 1932 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_21
timestamp 1688980957
transform 1 0 3036 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_27
timestamp 1688980957
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_29
timestamp 1688980957
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_41
timestamp 1688980957
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_53
timestamp 1688980957
transform 1 0 5980 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_77
timestamp 1688980957
transform 1 0 8188 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_108
timestamp 1688980957
transform 1 0 11040 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_138
timestamp 1688980957
transform 1 0 13800 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_141
timestamp 1688980957
transform 1 0 14076 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_153
timestamp 1688980957
transform 1 0 15180 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_165
timestamp 1688980957
transform 1 0 16284 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_177
timestamp 1688980957
transform 1 0 17388 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_189
timestamp 1688980957
transform 1 0 18492 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_195
timestamp 1688980957
transform 1 0 19044 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_197
timestamp 1688980957
transform 1 0 19228 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_209
timestamp 1688980957
transform 1 0 20332 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_221
timestamp 1688980957
transform 1 0 21436 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_233
timestamp 1688980957
transform 1 0 22540 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_245
timestamp 1688980957
transform 1 0 23644 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_251
timestamp 1688980957
transform 1 0 24196 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_253
timestamp 1688980957
transform 1 0 24380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_265
timestamp 1688980957
transform 1 0 25484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_277
timestamp 1688980957
transform 1 0 26588 0 1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_9
timestamp 1688980957
transform 1 0 1932 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_21
timestamp 1688980957
transform 1 0 3036 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_33
timestamp 1688980957
transform 1 0 4140 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_45
timestamp 1688980957
transform 1 0 5244 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_53
timestamp 1688980957
transform 1 0 5980 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_57
timestamp 1688980957
transform 1 0 6348 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_73
timestamp 1688980957
transform 1 0 7820 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_90
timestamp 1688980957
transform 1 0 9384 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_113
timestamp 1688980957
transform 1 0 11500 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_149
timestamp 1688980957
transform 1 0 14812 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_153
timestamp 1688980957
transform 1 0 15180 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_165
timestamp 1688980957
transform 1 0 16284 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_169
timestamp 1688980957
transform 1 0 16652 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_181
timestamp 1688980957
transform 1 0 17756 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_193
timestamp 1688980957
transform 1 0 18860 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_205
timestamp 1688980957
transform 1 0 19964 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_217
timestamp 1688980957
transform 1 0 21068 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_223
timestamp 1688980957
transform 1 0 21620 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_225
timestamp 1688980957
transform 1 0 21804 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_237
timestamp 1688980957
transform 1 0 22908 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_249
timestamp 1688980957
transform 1 0 24012 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_261
timestamp 1688980957
transform 1 0 25116 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_273
timestamp 1688980957
transform 1 0 26220 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_279
timestamp 1688980957
transform 1 0 26772 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_281
timestamp 1688980957
transform 1 0 26956 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_9
timestamp 1688980957
transform 1 0 1932 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_21
timestamp 1688980957
transform 1 0 3036 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_27
timestamp 1688980957
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_29
timestamp 1688980957
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_41
timestamp 1688980957
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_53
timestamp 1688980957
transform 1 0 5980 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_65
timestamp 1688980957
transform 1 0 7084 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_77
timestamp 1688980957
transform 1 0 8188 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_81
timestamp 1688980957
transform 1 0 8556 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_85
timestamp 1688980957
transform 1 0 8924 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_97
timestamp 1688980957
transform 1 0 10028 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_135
timestamp 1688980957
transform 1 0 13524 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_139
timestamp 1688980957
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_141
timestamp 1688980957
transform 1 0 14076 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_153
timestamp 1688980957
transform 1 0 15180 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_165
timestamp 1688980957
transform 1 0 16284 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_177
timestamp 1688980957
transform 1 0 17388 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_189
timestamp 1688980957
transform 1 0 18492 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_195
timestamp 1688980957
transform 1 0 19044 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_197
timestamp 1688980957
transform 1 0 19228 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_209
timestamp 1688980957
transform 1 0 20332 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_221
timestamp 1688980957
transform 1 0 21436 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_233
timestamp 1688980957
transform 1 0 22540 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_245
timestamp 1688980957
transform 1 0 23644 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_251
timestamp 1688980957
transform 1 0 24196 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_253
timestamp 1688980957
transform 1 0 24380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_265
timestamp 1688980957
transform 1 0 25484 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_277
timestamp 1688980957
transform 1 0 26588 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_289
timestamp 1688980957
transform 1 0 27692 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_297
timestamp 1688980957
transform 1 0 28428 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_9
timestamp 1688980957
transform 1 0 1932 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_21
timestamp 1688980957
transform 1 0 3036 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_33
timestamp 1688980957
transform 1 0 4140 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_45
timestamp 1688980957
transform 1 0 5244 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_53
timestamp 1688980957
transform 1 0 5980 0 -1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_57
timestamp 1688980957
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_69
timestamp 1688980957
transform 1 0 7452 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_81
timestamp 1688980957
transform 1 0 8556 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_87
timestamp 1688980957
transform 1 0 9108 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_98
timestamp 1688980957
transform 1 0 10120 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_110
timestamp 1688980957
transform 1 0 11224 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_113
timestamp 1688980957
transform 1 0 11500 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_134
timestamp 1688980957
transform 1 0 13432 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_146
timestamp 1688980957
transform 1 0 14536 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_158
timestamp 1688980957
transform 1 0 15640 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_166
timestamp 1688980957
transform 1 0 16376 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_169
timestamp 1688980957
transform 1 0 16652 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_181
timestamp 1688980957
transform 1 0 17756 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_193
timestamp 1688980957
transform 1 0 18860 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_205
timestamp 1688980957
transform 1 0 19964 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_217
timestamp 1688980957
transform 1 0 21068 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_223
timestamp 1688980957
transform 1 0 21620 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_225
timestamp 1688980957
transform 1 0 21804 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_237
timestamp 1688980957
transform 1 0 22908 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_249
timestamp 1688980957
transform 1 0 24012 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_261
timestamp 1688980957
transform 1 0 25116 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_273
timestamp 1688980957
transform 1 0 26220 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_277
timestamp 1688980957
transform 1 0 26588 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_281
timestamp 1688980957
transform 1 0 26956 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_9
timestamp 1688980957
transform 1 0 1932 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_21
timestamp 1688980957
transform 1 0 3036 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_27
timestamp 1688980957
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_29
timestamp 1688980957
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_41
timestamp 1688980957
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_53
timestamp 1688980957
transform 1 0 5980 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_65
timestamp 1688980957
transform 1 0 7084 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_77
timestamp 1688980957
transform 1 0 8188 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_83
timestamp 1688980957
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_85
timestamp 1688980957
transform 1 0 8924 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_97
timestamp 1688980957
transform 1 0 10028 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_109
timestamp 1688980957
transform 1 0 11132 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_121
timestamp 1688980957
transform 1 0 12236 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_125
timestamp 1688980957
transform 1 0 12604 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_128
timestamp 1688980957
transform 1 0 12880 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_141
timestamp 1688980957
transform 1 0 14076 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_153
timestamp 1688980957
transform 1 0 15180 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_165
timestamp 1688980957
transform 1 0 16284 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_177
timestamp 1688980957
transform 1 0 17388 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_189
timestamp 1688980957
transform 1 0 18492 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_195
timestamp 1688980957
transform 1 0 19044 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_197
timestamp 1688980957
transform 1 0 19228 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_209
timestamp 1688980957
transform 1 0 20332 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_221
timestamp 1688980957
transform 1 0 21436 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_233
timestamp 1688980957
transform 1 0 22540 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_245
timestamp 1688980957
transform 1 0 23644 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_251
timestamp 1688980957
transform 1 0 24196 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_253
timestamp 1688980957
transform 1 0 24380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_265
timestamp 1688980957
transform 1 0 25484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_277
timestamp 1688980957
transform 1 0 26588 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_9
timestamp 1688980957
transform 1 0 1932 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_21
timestamp 1688980957
transform 1 0 3036 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_33
timestamp 1688980957
transform 1 0 4140 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_45
timestamp 1688980957
transform 1 0 5244 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_53
timestamp 1688980957
transform 1 0 5980 0 -1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_57
timestamp 1688980957
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_69
timestamp 1688980957
transform 1 0 7452 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_81
timestamp 1688980957
transform 1 0 8556 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_93
timestamp 1688980957
transform 1 0 9660 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_105
timestamp 1688980957
transform 1 0 10764 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_111
timestamp 1688980957
transform 1 0 11316 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_113
timestamp 1688980957
transform 1 0 11500 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_125
timestamp 1688980957
transform 1 0 12604 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_137
timestamp 1688980957
transform 1 0 13708 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_149
timestamp 1688980957
transform 1 0 14812 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_161
timestamp 1688980957
transform 1 0 15916 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_167
timestamp 1688980957
transform 1 0 16468 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_169
timestamp 1688980957
transform 1 0 16652 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_181
timestamp 1688980957
transform 1 0 17756 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_193
timestamp 1688980957
transform 1 0 18860 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_205
timestamp 1688980957
transform 1 0 19964 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_217
timestamp 1688980957
transform 1 0 21068 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_223
timestamp 1688980957
transform 1 0 21620 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_225
timestamp 1688980957
transform 1 0 21804 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_237
timestamp 1688980957
transform 1 0 22908 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_249
timestamp 1688980957
transform 1 0 24012 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_261
timestamp 1688980957
transform 1 0 25116 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_273
timestamp 1688980957
transform 1 0 26220 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_279
timestamp 1688980957
transform 1 0 26772 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_281
timestamp 1688980957
transform 1 0 26956 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_293
timestamp 1688980957
transform 1 0 28060 0 -1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_9
timestamp 1688980957
transform 1 0 1932 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_21
timestamp 1688980957
transform 1 0 3036 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_27
timestamp 1688980957
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_29
timestamp 1688980957
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_41
timestamp 1688980957
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_53
timestamp 1688980957
transform 1 0 5980 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_65
timestamp 1688980957
transform 1 0 7084 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_77
timestamp 1688980957
transform 1 0 8188 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_83
timestamp 1688980957
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_85
timestamp 1688980957
transform 1 0 8924 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_97
timestamp 1688980957
transform 1 0 10028 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_109
timestamp 1688980957
transform 1 0 11132 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_121
timestamp 1688980957
transform 1 0 12236 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_133
timestamp 1688980957
transform 1 0 13340 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_139
timestamp 1688980957
transform 1 0 13892 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_141
timestamp 1688980957
transform 1 0 14076 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_153
timestamp 1688980957
transform 1 0 15180 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_165
timestamp 1688980957
transform 1 0 16284 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_177
timestamp 1688980957
transform 1 0 17388 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_189
timestamp 1688980957
transform 1 0 18492 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_195
timestamp 1688980957
transform 1 0 19044 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_197
timestamp 1688980957
transform 1 0 19228 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_209
timestamp 1688980957
transform 1 0 20332 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_221
timestamp 1688980957
transform 1 0 21436 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_233
timestamp 1688980957
transform 1 0 22540 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_245
timestamp 1688980957
transform 1 0 23644 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_251
timestamp 1688980957
transform 1 0 24196 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_253
timestamp 1688980957
transform 1 0 24380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_265
timestamp 1688980957
transform 1 0 25484 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_277
timestamp 1688980957
transform 1 0 26588 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_9
timestamp 1688980957
transform 1 0 1932 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_21
timestamp 1688980957
transform 1 0 3036 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_33
timestamp 1688980957
transform 1 0 4140 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_45
timestamp 1688980957
transform 1 0 5244 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_53
timestamp 1688980957
transform 1 0 5980 0 -1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_57
timestamp 1688980957
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_69
timestamp 1688980957
transform 1 0 7452 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_81
timestamp 1688980957
transform 1 0 8556 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_93
timestamp 1688980957
transform 1 0 9660 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_105
timestamp 1688980957
transform 1 0 10764 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_111
timestamp 1688980957
transform 1 0 11316 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_113
timestamp 1688980957
transform 1 0 11500 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_125
timestamp 1688980957
transform 1 0 12604 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_137
timestamp 1688980957
transform 1 0 13708 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_149
timestamp 1688980957
transform 1 0 14812 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_161
timestamp 1688980957
transform 1 0 15916 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_167
timestamp 1688980957
transform 1 0 16468 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_169
timestamp 1688980957
transform 1 0 16652 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_181
timestamp 1688980957
transform 1 0 17756 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_193
timestamp 1688980957
transform 1 0 18860 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_205
timestamp 1688980957
transform 1 0 19964 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_217
timestamp 1688980957
transform 1 0 21068 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_223
timestamp 1688980957
transform 1 0 21620 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_225
timestamp 1688980957
transform 1 0 21804 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_237
timestamp 1688980957
transform 1 0 22908 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_249
timestamp 1688980957
transform 1 0 24012 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_261
timestamp 1688980957
transform 1 0 25116 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_273
timestamp 1688980957
transform 1 0 26220 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_277
timestamp 1688980957
transform 1 0 26588 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_281
timestamp 1688980957
transform 1 0 26956 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_9
timestamp 1688980957
transform 1 0 1932 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_21
timestamp 1688980957
transform 1 0 3036 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_27
timestamp 1688980957
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_29
timestamp 1688980957
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_41
timestamp 1688980957
transform 1 0 4876 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_53
timestamp 1688980957
transform 1 0 5980 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_65
timestamp 1688980957
transform 1 0 7084 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_77
timestamp 1688980957
transform 1 0 8188 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_83
timestamp 1688980957
transform 1 0 8740 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_85
timestamp 1688980957
transform 1 0 8924 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_97
timestamp 1688980957
transform 1 0 10028 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_109
timestamp 1688980957
transform 1 0 11132 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_121
timestamp 1688980957
transform 1 0 12236 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_133
timestamp 1688980957
transform 1 0 13340 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_139
timestamp 1688980957
transform 1 0 13892 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_141
timestamp 1688980957
transform 1 0 14076 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_153
timestamp 1688980957
transform 1 0 15180 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_165
timestamp 1688980957
transform 1 0 16284 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_177
timestamp 1688980957
transform 1 0 17388 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_189
timestamp 1688980957
transform 1 0 18492 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_195
timestamp 1688980957
transform 1 0 19044 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_197
timestamp 1688980957
transform 1 0 19228 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_209
timestamp 1688980957
transform 1 0 20332 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_221
timestamp 1688980957
transform 1 0 21436 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_233
timestamp 1688980957
transform 1 0 22540 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_245
timestamp 1688980957
transform 1 0 23644 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_251
timestamp 1688980957
transform 1 0 24196 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_253
timestamp 1688980957
transform 1 0 24380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_265
timestamp 1688980957
transform 1 0 25484 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_277
timestamp 1688980957
transform 1 0 26588 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_289
timestamp 1688980957
transform 1 0 27692 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_297
timestamp 1688980957
transform 1 0 28428 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_9
timestamp 1688980957
transform 1 0 1932 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_21
timestamp 1688980957
transform 1 0 3036 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_33
timestamp 1688980957
transform 1 0 4140 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_45
timestamp 1688980957
transform 1 0 5244 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_53
timestamp 1688980957
transform 1 0 5980 0 -1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_57
timestamp 1688980957
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_69
timestamp 1688980957
transform 1 0 7452 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_81
timestamp 1688980957
transform 1 0 8556 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_93
timestamp 1688980957
transform 1 0 9660 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_105
timestamp 1688980957
transform 1 0 10764 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_111
timestamp 1688980957
transform 1 0 11316 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_113
timestamp 1688980957
transform 1 0 11500 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_125
timestamp 1688980957
transform 1 0 12604 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_137
timestamp 1688980957
transform 1 0 13708 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_149
timestamp 1688980957
transform 1 0 14812 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_161
timestamp 1688980957
transform 1 0 15916 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_167
timestamp 1688980957
transform 1 0 16468 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_169
timestamp 1688980957
transform 1 0 16652 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_181
timestamp 1688980957
transform 1 0 17756 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_193
timestamp 1688980957
transform 1 0 18860 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_205
timestamp 1688980957
transform 1 0 19964 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_217
timestamp 1688980957
transform 1 0 21068 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_223
timestamp 1688980957
transform 1 0 21620 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_225
timestamp 1688980957
transform 1 0 21804 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_237
timestamp 1688980957
transform 1 0 22908 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_249
timestamp 1688980957
transform 1 0 24012 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_261
timestamp 1688980957
transform 1 0 25116 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_273
timestamp 1688980957
transform 1 0 26220 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_277
timestamp 1688980957
transform 1 0 26588 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_281
timestamp 1688980957
transform 1 0 26956 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_9
timestamp 1688980957
transform 1 0 1932 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_21
timestamp 1688980957
transform 1 0 3036 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_27
timestamp 1688980957
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_29
timestamp 1688980957
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_41
timestamp 1688980957
transform 1 0 4876 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_53
timestamp 1688980957
transform 1 0 5980 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_65
timestamp 1688980957
transform 1 0 7084 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_77
timestamp 1688980957
transform 1 0 8188 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_83
timestamp 1688980957
transform 1 0 8740 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_85
timestamp 1688980957
transform 1 0 8924 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_97
timestamp 1688980957
transform 1 0 10028 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_109
timestamp 1688980957
transform 1 0 11132 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_121
timestamp 1688980957
transform 1 0 12236 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_133
timestamp 1688980957
transform 1 0 13340 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_139
timestamp 1688980957
transform 1 0 13892 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_141
timestamp 1688980957
transform 1 0 14076 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_153
timestamp 1688980957
transform 1 0 15180 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_165
timestamp 1688980957
transform 1 0 16284 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_177
timestamp 1688980957
transform 1 0 17388 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_189
timestamp 1688980957
transform 1 0 18492 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_195
timestamp 1688980957
transform 1 0 19044 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_197
timestamp 1688980957
transform 1 0 19228 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_209
timestamp 1688980957
transform 1 0 20332 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_221
timestamp 1688980957
transform 1 0 21436 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_233
timestamp 1688980957
transform 1 0 22540 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_245
timestamp 1688980957
transform 1 0 23644 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_251
timestamp 1688980957
transform 1 0 24196 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_253
timestamp 1688980957
transform 1 0 24380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_265
timestamp 1688980957
transform 1 0 25484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_277
timestamp 1688980957
transform 1 0 26588 0 1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_9
timestamp 1688980957
transform 1 0 1932 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_21
timestamp 1688980957
transform 1 0 3036 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_33
timestamp 1688980957
transform 1 0 4140 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_45
timestamp 1688980957
transform 1 0 5244 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_53
timestamp 1688980957
transform 1 0 5980 0 -1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_57
timestamp 1688980957
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_69
timestamp 1688980957
transform 1 0 7452 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_81
timestamp 1688980957
transform 1 0 8556 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_93
timestamp 1688980957
transform 1 0 9660 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_105
timestamp 1688980957
transform 1 0 10764 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_111
timestamp 1688980957
transform 1 0 11316 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_113
timestamp 1688980957
transform 1 0 11500 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_125
timestamp 1688980957
transform 1 0 12604 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_137
timestamp 1688980957
transform 1 0 13708 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_149
timestamp 1688980957
transform 1 0 14812 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_161
timestamp 1688980957
transform 1 0 15916 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_167
timestamp 1688980957
transform 1 0 16468 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_169
timestamp 1688980957
transform 1 0 16652 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_181
timestamp 1688980957
transform 1 0 17756 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_193
timestamp 1688980957
transform 1 0 18860 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_205
timestamp 1688980957
transform 1 0 19964 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_217
timestamp 1688980957
transform 1 0 21068 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_223
timestamp 1688980957
transform 1 0 21620 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_225
timestamp 1688980957
transform 1 0 21804 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_237
timestamp 1688980957
transform 1 0 22908 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_249
timestamp 1688980957
transform 1 0 24012 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_261
timestamp 1688980957
transform 1 0 25116 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_273
timestamp 1688980957
transform 1 0 26220 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_279
timestamp 1688980957
transform 1 0 26772 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_281
timestamp 1688980957
transform 1 0 26956 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_293
timestamp 1688980957
transform 1 0 28060 0 -1 22848
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_9
timestamp 1688980957
transform 1 0 1932 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_21
timestamp 1688980957
transform 1 0 3036 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_27
timestamp 1688980957
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_29
timestamp 1688980957
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_41
timestamp 1688980957
transform 1 0 4876 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_53
timestamp 1688980957
transform 1 0 5980 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_65
timestamp 1688980957
transform 1 0 7084 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_77
timestamp 1688980957
transform 1 0 8188 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_83
timestamp 1688980957
transform 1 0 8740 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_85
timestamp 1688980957
transform 1 0 8924 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_97
timestamp 1688980957
transform 1 0 10028 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_109
timestamp 1688980957
transform 1 0 11132 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_121
timestamp 1688980957
transform 1 0 12236 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_133
timestamp 1688980957
transform 1 0 13340 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_139
timestamp 1688980957
transform 1 0 13892 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_141
timestamp 1688980957
transform 1 0 14076 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_153
timestamp 1688980957
transform 1 0 15180 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_165
timestamp 1688980957
transform 1 0 16284 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_177
timestamp 1688980957
transform 1 0 17388 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_189
timestamp 1688980957
transform 1 0 18492 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_195
timestamp 1688980957
transform 1 0 19044 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_197
timestamp 1688980957
transform 1 0 19228 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_209
timestamp 1688980957
transform 1 0 20332 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_221
timestamp 1688980957
transform 1 0 21436 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_233
timestamp 1688980957
transform 1 0 22540 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_245
timestamp 1688980957
transform 1 0 23644 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_251
timestamp 1688980957
transform 1 0 24196 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_253
timestamp 1688980957
transform 1 0 24380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_265
timestamp 1688980957
transform 1 0 25484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_277
timestamp 1688980957
transform 1 0 26588 0 1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_6
timestamp 1688980957
transform 1 0 1656 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_18
timestamp 1688980957
transform 1 0 2760 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_30
timestamp 1688980957
transform 1 0 3864 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_42
timestamp 1688980957
transform 1 0 4968 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_54
timestamp 1688980957
transform 1 0 6072 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_57
timestamp 1688980957
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_69
timestamp 1688980957
transform 1 0 7452 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_81
timestamp 1688980957
transform 1 0 8556 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_93
timestamp 1688980957
transform 1 0 9660 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_105
timestamp 1688980957
transform 1 0 10764 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_111
timestamp 1688980957
transform 1 0 11316 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_113
timestamp 1688980957
transform 1 0 11500 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_125
timestamp 1688980957
transform 1 0 12604 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_137
timestamp 1688980957
transform 1 0 13708 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_149
timestamp 1688980957
transform 1 0 14812 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_161
timestamp 1688980957
transform 1 0 15916 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_167
timestamp 1688980957
transform 1 0 16468 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_169
timestamp 1688980957
transform 1 0 16652 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_181
timestamp 1688980957
transform 1 0 17756 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_193
timestamp 1688980957
transform 1 0 18860 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_205
timestamp 1688980957
transform 1 0 19964 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_217
timestamp 1688980957
transform 1 0 21068 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_223
timestamp 1688980957
transform 1 0 21620 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_225
timestamp 1688980957
transform 1 0 21804 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_237
timestamp 1688980957
transform 1 0 22908 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_249
timestamp 1688980957
transform 1 0 24012 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_261
timestamp 1688980957
transform 1 0 25116 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_273
timestamp 1688980957
transform 1 0 26220 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_277
timestamp 1688980957
transform 1 0 26588 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_281
timestamp 1688980957
transform 1 0 26956 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_3
timestamp 1688980957
transform 1 0 1380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_15
timestamp 1688980957
transform 1 0 2484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_27
timestamp 1688980957
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_29
timestamp 1688980957
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_41
timestamp 1688980957
transform 1 0 4876 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_53
timestamp 1688980957
transform 1 0 5980 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_65
timestamp 1688980957
transform 1 0 7084 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_77
timestamp 1688980957
transform 1 0 8188 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_83
timestamp 1688980957
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_85
timestamp 1688980957
transform 1 0 8924 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_97
timestamp 1688980957
transform 1 0 10028 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_109
timestamp 1688980957
transform 1 0 11132 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_121
timestamp 1688980957
transform 1 0 12236 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_133
timestamp 1688980957
transform 1 0 13340 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_139
timestamp 1688980957
transform 1 0 13892 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_141
timestamp 1688980957
transform 1 0 14076 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_153
timestamp 1688980957
transform 1 0 15180 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_165
timestamp 1688980957
transform 1 0 16284 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_177
timestamp 1688980957
transform 1 0 17388 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_189
timestamp 1688980957
transform 1 0 18492 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_195
timestamp 1688980957
transform 1 0 19044 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_197
timestamp 1688980957
transform 1 0 19228 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_209
timestamp 1688980957
transform 1 0 20332 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_221
timestamp 1688980957
transform 1 0 21436 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_233
timestamp 1688980957
transform 1 0 22540 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_245
timestamp 1688980957
transform 1 0 23644 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_251
timestamp 1688980957
transform 1 0 24196 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_253
timestamp 1688980957
transform 1 0 24380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_265
timestamp 1688980957
transform 1 0 25484 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_277
timestamp 1688980957
transform 1 0 26588 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_289
timestamp 1688980957
transform 1 0 27692 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_297
timestamp 1688980957
transform 1 0 28428 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_3
timestamp 1688980957
transform 1 0 1380 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_15
timestamp 1688980957
transform 1 0 2484 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_27
timestamp 1688980957
transform 1 0 3588 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_39
timestamp 1688980957
transform 1 0 4692 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_51
timestamp 1688980957
transform 1 0 5796 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_55
timestamp 1688980957
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_57
timestamp 1688980957
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_69
timestamp 1688980957
transform 1 0 7452 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_81
timestamp 1688980957
transform 1 0 8556 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_93
timestamp 1688980957
transform 1 0 9660 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_105
timestamp 1688980957
transform 1 0 10764 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_111
timestamp 1688980957
transform 1 0 11316 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_113
timestamp 1688980957
transform 1 0 11500 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_125
timestamp 1688980957
transform 1 0 12604 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_137
timestamp 1688980957
transform 1 0 13708 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_149
timestamp 1688980957
transform 1 0 14812 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_161
timestamp 1688980957
transform 1 0 15916 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_167
timestamp 1688980957
transform 1 0 16468 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_169
timestamp 1688980957
transform 1 0 16652 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_181
timestamp 1688980957
transform 1 0 17756 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_193
timestamp 1688980957
transform 1 0 18860 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_205
timestamp 1688980957
transform 1 0 19964 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_217
timestamp 1688980957
transform 1 0 21068 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_223
timestamp 1688980957
transform 1 0 21620 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_225
timestamp 1688980957
transform 1 0 21804 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_237
timestamp 1688980957
transform 1 0 22908 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_249
timestamp 1688980957
transform 1 0 24012 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_261
timestamp 1688980957
transform 1 0 25116 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_273
timestamp 1688980957
transform 1 0 26220 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_277
timestamp 1688980957
transform 1 0 26588 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_281
timestamp 1688980957
transform 1 0 26956 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_3
timestamp 1688980957
transform 1 0 1380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_15
timestamp 1688980957
transform 1 0 2484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_27
timestamp 1688980957
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_29
timestamp 1688980957
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_41
timestamp 1688980957
transform 1 0 4876 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_53
timestamp 1688980957
transform 1 0 5980 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_65
timestamp 1688980957
transform 1 0 7084 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_77
timestamp 1688980957
transform 1 0 8188 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_83
timestamp 1688980957
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_85
timestamp 1688980957
transform 1 0 8924 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_97
timestamp 1688980957
transform 1 0 10028 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_109
timestamp 1688980957
transform 1 0 11132 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_121
timestamp 1688980957
transform 1 0 12236 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_133
timestamp 1688980957
transform 1 0 13340 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_139
timestamp 1688980957
transform 1 0 13892 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_141
timestamp 1688980957
transform 1 0 14076 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_153
timestamp 1688980957
transform 1 0 15180 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_165
timestamp 1688980957
transform 1 0 16284 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_177
timestamp 1688980957
transform 1 0 17388 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_189
timestamp 1688980957
transform 1 0 18492 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_195
timestamp 1688980957
transform 1 0 19044 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_197
timestamp 1688980957
transform 1 0 19228 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_209
timestamp 1688980957
transform 1 0 20332 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_221
timestamp 1688980957
transform 1 0 21436 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_233
timestamp 1688980957
transform 1 0 22540 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_245
timestamp 1688980957
transform 1 0 23644 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_251
timestamp 1688980957
transform 1 0 24196 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_253
timestamp 1688980957
transform 1 0 24380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_265
timestamp 1688980957
transform 1 0 25484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_277
timestamp 1688980957
transform 1 0 26588 0 1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_3
timestamp 1688980957
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_15
timestamp 1688980957
transform 1 0 2484 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_27
timestamp 1688980957
transform 1 0 3588 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_39
timestamp 1688980957
transform 1 0 4692 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_51
timestamp 1688980957
transform 1 0 5796 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_55
timestamp 1688980957
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_57
timestamp 1688980957
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_69
timestamp 1688980957
transform 1 0 7452 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_81
timestamp 1688980957
transform 1 0 8556 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_93
timestamp 1688980957
transform 1 0 9660 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_105
timestamp 1688980957
transform 1 0 10764 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_111
timestamp 1688980957
transform 1 0 11316 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_113
timestamp 1688980957
transform 1 0 11500 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_125
timestamp 1688980957
transform 1 0 12604 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_137
timestamp 1688980957
transform 1 0 13708 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_149
timestamp 1688980957
transform 1 0 14812 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_161
timestamp 1688980957
transform 1 0 15916 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_167
timestamp 1688980957
transform 1 0 16468 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_169
timestamp 1688980957
transform 1 0 16652 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_181
timestamp 1688980957
transform 1 0 17756 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_193
timestamp 1688980957
transform 1 0 18860 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_205
timestamp 1688980957
transform 1 0 19964 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_217
timestamp 1688980957
transform 1 0 21068 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_223
timestamp 1688980957
transform 1 0 21620 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_225
timestamp 1688980957
transform 1 0 21804 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_237
timestamp 1688980957
transform 1 0 22908 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_249
timestamp 1688980957
transform 1 0 24012 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_261
timestamp 1688980957
transform 1 0 25116 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_273
timestamp 1688980957
transform 1 0 26220 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_279
timestamp 1688980957
transform 1 0 26772 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_281
timestamp 1688980957
transform 1 0 26956 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_293
timestamp 1688980957
transform 1 0 28060 0 -1 26112
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_3
timestamp 1688980957
transform 1 0 1380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_15
timestamp 1688980957
transform 1 0 2484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_27
timestamp 1688980957
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_29
timestamp 1688980957
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_41
timestamp 1688980957
transform 1 0 4876 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_53
timestamp 1688980957
transform 1 0 5980 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_65
timestamp 1688980957
transform 1 0 7084 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_77
timestamp 1688980957
transform 1 0 8188 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_83
timestamp 1688980957
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_85
timestamp 1688980957
transform 1 0 8924 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_97
timestamp 1688980957
transform 1 0 10028 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_109
timestamp 1688980957
transform 1 0 11132 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_121
timestamp 1688980957
transform 1 0 12236 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_133
timestamp 1688980957
transform 1 0 13340 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_139
timestamp 1688980957
transform 1 0 13892 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_141
timestamp 1688980957
transform 1 0 14076 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_153
timestamp 1688980957
transform 1 0 15180 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_165
timestamp 1688980957
transform 1 0 16284 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_177
timestamp 1688980957
transform 1 0 17388 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_189
timestamp 1688980957
transform 1 0 18492 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_195
timestamp 1688980957
transform 1 0 19044 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_197
timestamp 1688980957
transform 1 0 19228 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_209
timestamp 1688980957
transform 1 0 20332 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_221
timestamp 1688980957
transform 1 0 21436 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_233
timestamp 1688980957
transform 1 0 22540 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_245
timestamp 1688980957
transform 1 0 23644 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_251
timestamp 1688980957
transform 1 0 24196 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_253
timestamp 1688980957
transform 1 0 24380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_265
timestamp 1688980957
transform 1 0 25484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_44_277
timestamp 1688980957
transform 1 0 26588 0 1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_3
timestamp 1688980957
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_15
timestamp 1688980957
transform 1 0 2484 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_27
timestamp 1688980957
transform 1 0 3588 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_39
timestamp 1688980957
transform 1 0 4692 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_51
timestamp 1688980957
transform 1 0 5796 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_55
timestamp 1688980957
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_57
timestamp 1688980957
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_69
timestamp 1688980957
transform 1 0 7452 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_81
timestamp 1688980957
transform 1 0 8556 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_93
timestamp 1688980957
transform 1 0 9660 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_105
timestamp 1688980957
transform 1 0 10764 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_111
timestamp 1688980957
transform 1 0 11316 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_113
timestamp 1688980957
transform 1 0 11500 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_125
timestamp 1688980957
transform 1 0 12604 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_137
timestamp 1688980957
transform 1 0 13708 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_149
timestamp 1688980957
transform 1 0 14812 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_161
timestamp 1688980957
transform 1 0 15916 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_167
timestamp 1688980957
transform 1 0 16468 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_169
timestamp 1688980957
transform 1 0 16652 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_181
timestamp 1688980957
transform 1 0 17756 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_193
timestamp 1688980957
transform 1 0 18860 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_205
timestamp 1688980957
transform 1 0 19964 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_217
timestamp 1688980957
transform 1 0 21068 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_223
timestamp 1688980957
transform 1 0 21620 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_225
timestamp 1688980957
transform 1 0 21804 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_237
timestamp 1688980957
transform 1 0 22908 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_249
timestamp 1688980957
transform 1 0 24012 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_261
timestamp 1688980957
transform 1 0 25116 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_273
timestamp 1688980957
transform 1 0 26220 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_277
timestamp 1688980957
transform 1 0 26588 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_281
timestamp 1688980957
transform 1 0 26956 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_3
timestamp 1688980957
transform 1 0 1380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_15
timestamp 1688980957
transform 1 0 2484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_27
timestamp 1688980957
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_29
timestamp 1688980957
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_41
timestamp 1688980957
transform 1 0 4876 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_53
timestamp 1688980957
transform 1 0 5980 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_57
timestamp 1688980957
transform 1 0 6348 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_69
timestamp 1688980957
transform 1 0 7452 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_81
timestamp 1688980957
transform 1 0 8556 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_85
timestamp 1688980957
transform 1 0 8924 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_97
timestamp 1688980957
transform 1 0 10028 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_109
timestamp 1688980957
transform 1 0 11132 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_113
timestamp 1688980957
transform 1 0 11500 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_125
timestamp 1688980957
transform 1 0 12604 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_137
timestamp 1688980957
transform 1 0 13708 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_141
timestamp 1688980957
transform 1 0 14076 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_153
timestamp 1688980957
transform 1 0 15180 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_165
timestamp 1688980957
transform 1 0 16284 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_169
timestamp 1688980957
transform 1 0 16652 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_181
timestamp 1688980957
transform 1 0 17756 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_193
timestamp 1688980957
transform 1 0 18860 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_197
timestamp 1688980957
transform 1 0 19228 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_209
timestamp 1688980957
transform 1 0 20332 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_221
timestamp 1688980957
transform 1 0 21436 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_225
timestamp 1688980957
transform 1 0 21804 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_237
timestamp 1688980957
transform 1 0 22908 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_249
timestamp 1688980957
transform 1 0 24012 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_253
timestamp 1688980957
transform 1 0 24380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_265
timestamp 1688980957
transform 1 0 25484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_277
timestamp 1688980957
transform 1 0 26588 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_281
timestamp 1688980957
transform 1 0 26956 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_293
timestamp 1688980957
transform 1 0 28060 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1840 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp 1688980957
transform -1 0 2668 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp 1688980957
transform 1 0 1840 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp 1688980957
transform -1 0 4048 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold5
timestamp 1688980957
transform 1 0 2576 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold6
timestamp 1688980957
transform 1 0 1472 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold7
timestamp 1688980957
transform -1 0 3680 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold8
timestamp 1688980957
transform -1 0 2392 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold9
timestamp 1688980957
transform -1 0 4600 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold10
timestamp 1688980957
transform 1 0 1380 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold11
timestamp 1688980957
transform 1 0 2852 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold12
timestamp 1688980957
transform -1 0 7084 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold13
timestamp 1688980957
transform 1 0 8556 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold14
timestamp 1688980957
transform 1 0 2944 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold15
timestamp 1688980957
transform -1 0 6072 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold16
timestamp 1688980957
transform 1 0 1472 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold17
timestamp 1688980957
transform -1 0 5888 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold18
timestamp 1688980957
transform -1 0 6256 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold19
timestamp 1688980957
transform 1 0 8924 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold20
timestamp 1688980957
transform -1 0 6624 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold21
timestamp 1688980957
transform -1 0 6164 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold22
timestamp 1688980957
transform 1 0 2944 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold23
timestamp 1688980957
transform -1 0 5336 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold24
timestamp 1688980957
transform -1 0 6072 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold25
timestamp 1688980957
transform 1 0 1380 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold26
timestamp 1688980957
transform 1 0 1472 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold27
timestamp 1688980957
transform -1 0 7360 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold28
timestamp 1688980957
transform 1 0 5520 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold29
timestamp 1688980957
transform -1 0 7820 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold30
timestamp 1688980957
transform 1 0 8096 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold31
timestamp 1688980957
transform 1 0 2116 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold32
timestamp 1688980957
transform 1 0 2208 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold33
timestamp 1688980957
transform 1 0 7268 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold34
timestamp 1688980957
transform 1 0 2208 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold35
timestamp 1688980957
transform -1 0 6164 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold36
timestamp 1688980957
transform -1 0 10488 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold37
timestamp 1688980957
transform 1 0 7820 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold38
timestamp 1688980957
transform 1 0 4416 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold39
timestamp 1688980957
transform -1 0 10212 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold40
timestamp 1688980957
transform -1 0 10580 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold41
timestamp 1688980957
transform 1 0 10304 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold42
timestamp 1688980957
transform -1 0 10580 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold43
timestamp 1688980957
transform 1 0 11500 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold44
timestamp 1688980957
transform -1 0 12236 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold45
timestamp 1688980957
transform -1 0 13432 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold46
timestamp 1688980957
transform 1 0 7360 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold47
timestamp 1688980957
transform -1 0 9660 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold48
timestamp 1688980957
transform -1 0 8832 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold49
timestamp 1688980957
transform 1 0 7912 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold50
timestamp 1688980957
transform -1 0 8924 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold51
timestamp 1688980957
transform 1 0 10672 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold52
timestamp 1688980957
transform 1 0 9936 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold53
timestamp 1688980957
transform -1 0 11776 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold54
timestamp 1688980957
transform -1 0 13800 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold55
timestamp 1688980957
transform -1 0 7360 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold56
timestamp 1688980957
transform 1 0 8924 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold57
timestamp 1688980957
transform -1 0 13800 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold58
timestamp 1688980957
transform -1 0 4784 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold59
timestamp 1688980957
transform 1 0 4324 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold60
timestamp 1688980957
transform -1 0 12604 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold61
timestamp 1688980957
transform 1 0 4784 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold62
timestamp 1688980957
transform -1 0 7084 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold63
timestamp 1688980957
transform -1 0 9660 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold64
timestamp 1688980957
transform 1 0 7084 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold65
timestamp 1688980957
transform -1 0 7084 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold66
timestamp 1688980957
transform -1 0 6256 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold67
timestamp 1688980957
transform 1 0 6900 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold68
timestamp 1688980957
transform -1 0 7912 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold69
timestamp 1688980957
transform -1 0 7084 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold70
timestamp 1688980957
transform 1 0 10672 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold71
timestamp 1688980957
transform -1 0 11408 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold72
timestamp 1688980957
transform -1 0 14812 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold73
timestamp 1688980957
transform 1 0 8372 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold74
timestamp 1688980957
transform -1 0 8832 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold75
timestamp 1688980957
transform -1 0 10028 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold76
timestamp 1688980957
transform 1 0 9200 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold77
timestamp 1688980957
transform 1 0 9200 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold78
timestamp 1688980957
transform 1 0 10672 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold79
timestamp 1688980957
transform 1 0 9752 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold80
timestamp 1688980957
transform -1 0 10304 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold81
timestamp 1688980957
transform -1 0 14536 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold82
timestamp 1688980957
transform -1 0 8832 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold83
timestamp 1688980957
transform 1 0 7912 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold84
timestamp 1688980957
transform -1 0 11132 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold85
timestamp 1688980957
transform -1 0 11316 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold86
timestamp 1688980957
transform -1 0 11224 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold87
timestamp 1688980957
transform -1 0 13432 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold88
timestamp 1688980957
transform 1 0 7636 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold89
timestamp 1688980957
transform 1 0 6348 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold90
timestamp 1688980957
transform -1 0 7360 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold91
timestamp 1688980957
transform 1 0 9108 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold92
timestamp 1688980957
transform 1 0 7912 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold93
timestamp 1688980957
transform -1 0 12696 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold94
timestamp 1688980957
transform 1 0 2944 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold95
timestamp 1688980957
transform 1 0 2116 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input1 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 2944 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1688980957
transform -1 0 1932 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1688980957
transform -1 0 1656 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input4 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1656 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input5
timestamp 1688980957
transform 1 0 1380 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1688980957
transform -1 0 1932 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input7
timestamp 1688980957
transform 1 0 1380 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1688980957
transform -1 0 1932 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input9
timestamp 1688980957
transform 1 0 1380 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input10
timestamp 1688980957
transform 1 0 1656 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1688980957
transform -1 0 1656 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1688980957
transform -1 0 2484 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input13
timestamp 1688980957
transform 1 0 1656 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 1688980957
transform -1 0 1656 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input15
timestamp 1688980957
transform 1 0 1656 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input16
timestamp 1688980957
transform 1 0 1380 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input17
timestamp 1688980957
transform 1 0 1656 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input18
timestamp 1688980957
transform 1 0 1380 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input19
timestamp 1688980957
transform 1 0 1656 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input20
timestamp 1688980957
transform 1 0 1380 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input21
timestamp 1688980957
transform 1 0 1656 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input22
timestamp 1688980957
transform 1 0 1380 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input23
timestamp 1688980957
transform -1 0 2484 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input24
timestamp 1688980957
transform 1 0 1380 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input25
timestamp 1688980957
transform -1 0 1840 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input26
timestamp 1688980957
transform -1 0 3588 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input27
timestamp 1688980957
transform -1 0 2208 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input28
timestamp 1688980957
transform -1 0 1932 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input29
timestamp 1688980957
transform -1 0 1656 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input30
timestamp 1688980957
transform -1 0 1932 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input31
timestamp 1688980957
transform -1 0 1656 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input32
timestamp 1688980957
transform -1 0 1932 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input33
timestamp 1688980957
transform 1 0 1380 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input34
timestamp 1688980957
transform -1 0 1932 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input35
timestamp 1688980957
transform -1 0 1656 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input36
timestamp 1688980957
transform -1 0 1932 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input37
timestamp 1688980957
transform -1 0 1656 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input38
timestamp 1688980957
transform 1 0 1656 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input39
timestamp 1688980957
transform -1 0 1656 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input40
timestamp 1688980957
transform 1 0 1656 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input41
timestamp 1688980957
transform 1 0 1380 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input42
timestamp 1688980957
transform -1 0 1932 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input43
timestamp 1688980957
transform -1 0 1656 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input44
timestamp 1688980957
transform 1 0 1380 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input45
timestamp 1688980957
transform -1 0 1932 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input46
timestamp 1688980957
transform -1 0 1656 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input47
timestamp 1688980957
transform -1 0 1932 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input48
timestamp 1688980957
transform -1 0 1656 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input49
timestamp 1688980957
transform 1 0 1656 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input50
timestamp 1688980957
transform 1 0 1380 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input51
timestamp 1688980957
transform 1 0 1656 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input52
timestamp 1688980957
transform 1 0 1380 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input53
timestamp 1688980957
transform 1 0 1656 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input54
timestamp 1688980957
transform -1 0 1932 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input55
timestamp 1688980957
transform 1 0 1380 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input56
timestamp 1688980957
transform 1 0 1380 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input57
timestamp 1688980957
transform -1 0 1932 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input58
timestamp 1688980957
transform 1 0 1380 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input59
timestamp 1688980957
transform 1 0 1656 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input60
timestamp 1688980957
transform 1 0 1380 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input61
timestamp 1688980957
transform -1 0 1656 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input62
timestamp 1688980957
transform -1 0 1932 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input63
timestamp 1688980957
transform 1 0 2484 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input64
timestamp 1688980957
transform -1 0 2484 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input65
timestamp 1688980957
transform -1 0 13340 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input66
timestamp 1688980957
transform 1 0 11316 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input67
timestamp 1688980957
transform -1 0 13064 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input68
timestamp 1688980957
transform -1 0 1748 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input69
timestamp 1688980957
transform 1 0 8740 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input70
timestamp 1688980957
transform 1 0 12052 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input71
timestamp 1688980957
transform 1 0 10304 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input72
timestamp 1688980957
transform 1 0 7912 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input73
timestamp 1688980957
transform -1 0 4048 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input74
timestamp 1688980957
transform -1 0 8740 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input75
timestamp 1688980957
transform 1 0 8188 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input76
timestamp 1688980957
transform 1 0 2484 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input77
timestamp 1688980957
transform 1 0 11776 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input78
timestamp 1688980957
transform 1 0 9384 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input79
timestamp 1688980957
transform -1 0 6624 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input80
timestamp 1688980957
transform 1 0 11040 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input81
timestamp 1688980957
transform 1 0 10028 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input82
timestamp 1688980957
transform 1 0 10764 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input83
timestamp 1688980957
transform -1 0 9200 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input84
timestamp 1688980957
transform -1 0 10764 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input85
timestamp 1688980957
transform 1 0 12512 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input86
timestamp 1688980957
transform 1 0 11500 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input87
timestamp 1688980957
transform -1 0 2484 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input88
timestamp 1688980957
transform 1 0 12236 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input89
timestamp 1688980957
transform 1 0 3036 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input90
timestamp 1688980957
transform 1 0 2484 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input91
timestamp 1688980957
transform -1 0 3036 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input92
timestamp 1688980957
transform 1 0 9016 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input93
timestamp 1688980957
transform 1 0 12328 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input94
timestamp 1688980957
transform 1 0 9660 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input95
timestamp 1688980957
transform 1 0 8188 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input96
timestamp 1688980957
transform -1 0 2208 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input97
timestamp 1688980957
transform 1 0 1932 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_12  output98 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 20240 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output99
timestamp 1688980957
transform 1 0 27140 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output100
timestamp 1688980957
transform 1 0 27140 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output101
timestamp 1688980957
transform 1 0 27140 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output102
timestamp 1688980957
transform 1 0 27140 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output103
timestamp 1688980957
transform 1 0 27140 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output104
timestamp 1688980957
transform 1 0 27140 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output105
timestamp 1688980957
transform 1 0 27140 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output106
timestamp 1688980957
transform 1 0 27140 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output107
timestamp 1688980957
transform 1 0 27140 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output108
timestamp 1688980957
transform 1 0 27140 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output109
timestamp 1688980957
transform 1 0 23920 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output110
timestamp 1688980957
transform 1 0 27140 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output111
timestamp 1688980957
transform 1 0 27140 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output112
timestamp 1688980957
transform 1 0 27140 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output113
timestamp 1688980957
transform 1 0 27140 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output114
timestamp 1688980957
transform 1 0 27140 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output115
timestamp 1688980957
transform 1 0 27140 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output116
timestamp 1688980957
transform 1 0 27140 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output117
timestamp 1688980957
transform 1 0 27140 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output118
timestamp 1688980957
transform 1 0 27140 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output119
timestamp 1688980957
transform 1 0 27140 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output120
timestamp 1688980957
transform 1 0 25668 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output121
timestamp 1688980957
transform 1 0 27140 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output122
timestamp 1688980957
transform 1 0 27140 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output123
timestamp 1688980957
transform 1 0 27140 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output124
timestamp 1688980957
transform 1 0 27140 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output125
timestamp 1688980957
transform 1 0 27140 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output126
timestamp 1688980957
transform 1 0 27140 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output127
timestamp 1688980957
transform 1 0 27140 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output128
timestamp 1688980957
transform 1 0 27140 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output129
timestamp 1688980957
transform 1 0 20240 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output130
timestamp 1688980957
transform 1 0 21804 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output131
timestamp 1688980957
transform 1 0 24380 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output132
timestamp 1688980957
transform 1 0 25300 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output133
timestamp 1688980957
transform 1 0 25852 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output134
timestamp 1688980957
transform 1 0 26956 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output135
timestamp 1688980957
transform 1 0 24840 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output136
timestamp 1688980957
transform 1 0 25852 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output137
timestamp 1688980957
transform 1 0 26956 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output138
timestamp 1688980957
transform 1 0 25668 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output139
timestamp 1688980957
transform 1 0 26956 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output140
timestamp 1688980957
transform 1 0 25392 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output141
timestamp 1688980957
transform 1 0 21804 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output142
timestamp 1688980957
transform 1 0 22816 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output143
timestamp 1688980957
transform 1 0 23368 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output144
timestamp 1688980957
transform 1 0 20240 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output145
timestamp 1688980957
transform 1 0 20056 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output146
timestamp 1688980957
transform 1 0 27140 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output147
timestamp 1688980957
transform 1 0 22816 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output148
timestamp 1688980957
transform 1 0 21896 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output149
timestamp 1688980957
transform 1 0 21344 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output150
timestamp 1688980957
transform 1 0 18768 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output151
timestamp 1688980957
transform 1 0 17664 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output152
timestamp 1688980957
transform 1 0 21528 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output153
timestamp 1688980957
transform 1 0 25392 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output154
timestamp 1688980957
transform 1 0 23276 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output155
timestamp 1688980957
transform 1 0 24380 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output156
timestamp 1688980957
transform 1 0 22356 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output157
timestamp 1688980957
transform 1 0 24748 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output158
timestamp 1688980957
transform 1 0 24380 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output159
timestamp 1688980957
transform 1 0 23828 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output160
timestamp 1688980957
transform 1 0 26956 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1688980957
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1688980957
transform -1 0 28888 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1688980957
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1688980957
transform -1 0 28888 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1688980957
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1688980957
transform -1 0 28888 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1688980957
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1688980957
transform -1 0 28888 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1688980957
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1688980957
transform -1 0 28888 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1688980957
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1688980957
transform -1 0 28888 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1688980957
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1688980957
transform -1 0 28888 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1688980957
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1688980957
transform -1 0 28888 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1688980957
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1688980957
transform -1 0 28888 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1688980957
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1688980957
transform -1 0 28888 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1688980957
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1688980957
transform -1 0 28888 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1688980957
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1688980957
transform -1 0 28888 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1688980957
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1688980957
transform -1 0 28888 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1688980957
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1688980957
transform -1 0 28888 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1688980957
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1688980957
transform -1 0 28888 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1688980957
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1688980957
transform -1 0 28888 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1688980957
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1688980957
transform -1 0 28888 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1688980957
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1688980957
transform -1 0 28888 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1688980957
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1688980957
transform -1 0 28888 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1688980957
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1688980957
transform -1 0 28888 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1688980957
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1688980957
transform -1 0 28888 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1688980957
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1688980957
transform -1 0 28888 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1688980957
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1688980957
transform -1 0 28888 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1688980957
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1688980957
transform -1 0 28888 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1688980957
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1688980957
transform -1 0 28888 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1688980957
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1688980957
transform -1 0 28888 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1688980957
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1688980957
transform -1 0 28888 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1688980957
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1688980957
transform -1 0 28888 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1688980957
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1688980957
transform -1 0 28888 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1688980957
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1688980957
transform -1 0 28888 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1688980957
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1688980957
transform -1 0 28888 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1688980957
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1688980957
transform -1 0 28888 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1688980957
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1688980957
transform -1 0 28888 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1688980957
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1688980957
transform -1 0 28888 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1688980957
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1688980957
transform -1 0 28888 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1688980957
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1688980957
transform -1 0 28888 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1688980957
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1688980957
transform -1 0 28888 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1688980957
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1688980957
transform -1 0 28888 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1688980957
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1688980957
transform -1 0 28888 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1688980957
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1688980957
transform -1 0 28888 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1688980957
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1688980957
transform -1 0 28888 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1688980957
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1688980957
transform -1 0 28888 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1688980957
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1688980957
transform -1 0 28888 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1688980957
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1688980957
transform -1 0 28888 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1688980957
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1688980957
transform -1 0 28888 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1688980957
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1688980957
transform -1 0 28888 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1688980957
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1688980957
transform -1 0 28888 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1688980957
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1688980957
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1688980957
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1688980957
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1688980957
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1688980957
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1688980957
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1688980957
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1688980957
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1688980957
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1688980957
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1688980957
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1688980957
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1688980957
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1688980957
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1688980957
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1688980957
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1688980957
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1688980957
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1688980957
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1688980957
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1688980957
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1688980957
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1688980957
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1688980957
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1688980957
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1688980957
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1688980957
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1688980957
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1688980957
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1688980957
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1688980957
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1688980957
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1688980957
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1688980957
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1688980957
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1688980957
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1688980957
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1688980957
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1688980957
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1688980957
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1688980957
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1688980957
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1688980957
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1688980957
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1688980957
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1688980957
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1688980957
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1688980957
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1688980957
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1688980957
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1688980957
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1688980957
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1688980957
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1688980957
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1688980957
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1688980957
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1688980957
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1688980957
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1688980957
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1688980957
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1688980957
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1688980957
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1688980957
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1688980957
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1688980957
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1688980957
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1688980957
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1688980957
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1688980957
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1688980957
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1688980957
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1688980957
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1688980957
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1688980957
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1688980957
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1688980957
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1688980957
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1688980957
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1688980957
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1688980957
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1688980957
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1688980957
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1688980957
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1688980957
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1688980957
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1688980957
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1688980957
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1688980957
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1688980957
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1688980957
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1688980957
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1688980957
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1688980957
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1688980957
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1688980957
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1688980957
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1688980957
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1688980957
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1688980957
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1688980957
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1688980957
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1688980957
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1688980957
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1688980957
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1688980957
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1688980957
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1688980957
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1688980957
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1688980957
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1688980957
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1688980957
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1688980957
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1688980957
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1688980957
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1688980957
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1688980957
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1688980957
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1688980957
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1688980957
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1688980957
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1688980957
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1688980957
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1688980957
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1688980957
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1688980957
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1688980957
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1688980957
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1688980957
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1688980957
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1688980957
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1688980957
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1688980957
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1688980957
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1688980957
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1688980957
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1688980957
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1688980957
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1688980957
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1688980957
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1688980957
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1688980957
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1688980957
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1688980957
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1688980957
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1688980957
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1688980957
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1688980957
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1688980957
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1688980957
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1688980957
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1688980957
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1688980957
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1688980957
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1688980957
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1688980957
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1688980957
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1688980957
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1688980957
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1688980957
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1688980957
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1688980957
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1688980957
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1688980957
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1688980957
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1688980957
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1688980957
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1688980957
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1688980957
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1688980957
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1688980957
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1688980957
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1688980957
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1688980957
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1688980957
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1688980957
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1688980957
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1688980957
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1688980957
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1688980957
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1688980957
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1688980957
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1688980957
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1688980957
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1688980957
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1688980957
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1688980957
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1688980957
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1688980957
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1688980957
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1688980957
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1688980957
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1688980957
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1688980957
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1688980957
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1688980957
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1688980957
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1688980957
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1688980957
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1688980957
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1688980957
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1688980957
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1688980957
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1688980957
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1688980957
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1688980957
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1688980957
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1688980957
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1688980957
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1688980957
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1688980957
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1688980957
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1688980957
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1688980957
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1688980957
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1688980957
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1688980957
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1688980957
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1688980957
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1688980957
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1688980957
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1688980957
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1688980957
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1688980957
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1688980957
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1688980957
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1688980957
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1688980957
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1688980957
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1688980957
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1688980957
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1688980957
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1688980957
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1688980957
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1688980957
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1688980957
transform 1 0 6256 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1688980957
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1688980957
transform 1 0 11408 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1688980957
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1688980957
transform 1 0 16560 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1688980957
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1688980957
transform 1 0 21712 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1688980957
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1688980957
transform 1 0 26864 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  wishbone_register_m_165 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 28336 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  wishbone_register_m_166
timestamp 1688980957
transform 1 0 28336 0 1 3264
box -38 -48 314 592
<< labels >>
flabel metal3 s 0 6264 800 6384 0 FreeSans 480 0 0 0 access_read_mask_i[0]
port 0 nsew signal input
flabel metal3 s 0 8984 800 9104 0 FreeSans 480 0 0 0 access_read_mask_i[10]
port 1 nsew signal input
flabel metal3 s 0 9256 800 9376 0 FreeSans 480 0 0 0 access_read_mask_i[11]
port 2 nsew signal input
flabel metal3 s 0 9528 800 9648 0 FreeSans 480 0 0 0 access_read_mask_i[12]
port 3 nsew signal input
flabel metal3 s 0 9800 800 9920 0 FreeSans 480 0 0 0 access_read_mask_i[13]
port 4 nsew signal input
flabel metal3 s 0 10072 800 10192 0 FreeSans 480 0 0 0 access_read_mask_i[14]
port 5 nsew signal input
flabel metal3 s 0 10344 800 10464 0 FreeSans 480 0 0 0 access_read_mask_i[15]
port 6 nsew signal input
flabel metal3 s 0 10616 800 10736 0 FreeSans 480 0 0 0 access_read_mask_i[16]
port 7 nsew signal input
flabel metal3 s 0 10888 800 11008 0 FreeSans 480 0 0 0 access_read_mask_i[17]
port 8 nsew signal input
flabel metal3 s 0 11160 800 11280 0 FreeSans 480 0 0 0 access_read_mask_i[18]
port 9 nsew signal input
flabel metal3 s 0 11432 800 11552 0 FreeSans 480 0 0 0 access_read_mask_i[19]
port 10 nsew signal input
flabel metal3 s 0 6536 800 6656 0 FreeSans 480 0 0 0 access_read_mask_i[1]
port 11 nsew signal input
flabel metal3 s 0 11704 800 11824 0 FreeSans 480 0 0 0 access_read_mask_i[20]
port 12 nsew signal input
flabel metal3 s 0 11976 800 12096 0 FreeSans 480 0 0 0 access_read_mask_i[21]
port 13 nsew signal input
flabel metal3 s 0 12248 800 12368 0 FreeSans 480 0 0 0 access_read_mask_i[22]
port 14 nsew signal input
flabel metal3 s 0 12520 800 12640 0 FreeSans 480 0 0 0 access_read_mask_i[23]
port 15 nsew signal input
flabel metal3 s 0 12792 800 12912 0 FreeSans 480 0 0 0 access_read_mask_i[24]
port 16 nsew signal input
flabel metal3 s 0 13064 800 13184 0 FreeSans 480 0 0 0 access_read_mask_i[25]
port 17 nsew signal input
flabel metal3 s 0 13336 800 13456 0 FreeSans 480 0 0 0 access_read_mask_i[26]
port 18 nsew signal input
flabel metal3 s 0 13608 800 13728 0 FreeSans 480 0 0 0 access_read_mask_i[27]
port 19 nsew signal input
flabel metal3 s 0 13880 800 14000 0 FreeSans 480 0 0 0 access_read_mask_i[28]
port 20 nsew signal input
flabel metal3 s 0 14152 800 14272 0 FreeSans 480 0 0 0 access_read_mask_i[29]
port 21 nsew signal input
flabel metal3 s 0 6808 800 6928 0 FreeSans 480 0 0 0 access_read_mask_i[2]
port 22 nsew signal input
flabel metal3 s 0 14424 800 14544 0 FreeSans 480 0 0 0 access_read_mask_i[30]
port 23 nsew signal input
flabel metal3 s 0 14696 800 14816 0 FreeSans 480 0 0 0 access_read_mask_i[31]
port 24 nsew signal input
flabel metal3 s 0 7080 800 7200 0 FreeSans 480 0 0 0 access_read_mask_i[3]
port 25 nsew signal input
flabel metal3 s 0 7352 800 7472 0 FreeSans 480 0 0 0 access_read_mask_i[4]
port 26 nsew signal input
flabel metal3 s 0 7624 800 7744 0 FreeSans 480 0 0 0 access_read_mask_i[5]
port 27 nsew signal input
flabel metal3 s 0 7896 800 8016 0 FreeSans 480 0 0 0 access_read_mask_i[6]
port 28 nsew signal input
flabel metal3 s 0 8168 800 8288 0 FreeSans 480 0 0 0 access_read_mask_i[7]
port 29 nsew signal input
flabel metal3 s 0 8440 800 8560 0 FreeSans 480 0 0 0 access_read_mask_i[8]
port 30 nsew signal input
flabel metal3 s 0 8712 800 8832 0 FreeSans 480 0 0 0 access_read_mask_i[9]
port 31 nsew signal input
flabel metal3 s 0 14968 800 15088 0 FreeSans 480 0 0 0 access_write_mask_i[0]
port 32 nsew signal input
flabel metal3 s 0 17688 800 17808 0 FreeSans 480 0 0 0 access_write_mask_i[10]
port 33 nsew signal input
flabel metal3 s 0 17960 800 18080 0 FreeSans 480 0 0 0 access_write_mask_i[11]
port 34 nsew signal input
flabel metal3 s 0 18232 800 18352 0 FreeSans 480 0 0 0 access_write_mask_i[12]
port 35 nsew signal input
flabel metal3 s 0 18504 800 18624 0 FreeSans 480 0 0 0 access_write_mask_i[13]
port 36 nsew signal input
flabel metal3 s 0 18776 800 18896 0 FreeSans 480 0 0 0 access_write_mask_i[14]
port 37 nsew signal input
flabel metal3 s 0 19048 800 19168 0 FreeSans 480 0 0 0 access_write_mask_i[15]
port 38 nsew signal input
flabel metal3 s 0 19320 800 19440 0 FreeSans 480 0 0 0 access_write_mask_i[16]
port 39 nsew signal input
flabel metal3 s 0 19592 800 19712 0 FreeSans 480 0 0 0 access_write_mask_i[17]
port 40 nsew signal input
flabel metal3 s 0 19864 800 19984 0 FreeSans 480 0 0 0 access_write_mask_i[18]
port 41 nsew signal input
flabel metal3 s 0 20136 800 20256 0 FreeSans 480 0 0 0 access_write_mask_i[19]
port 42 nsew signal input
flabel metal3 s 0 15240 800 15360 0 FreeSans 480 0 0 0 access_write_mask_i[1]
port 43 nsew signal input
flabel metal3 s 0 20408 800 20528 0 FreeSans 480 0 0 0 access_write_mask_i[20]
port 44 nsew signal input
flabel metal3 s 0 20680 800 20800 0 FreeSans 480 0 0 0 access_write_mask_i[21]
port 45 nsew signal input
flabel metal3 s 0 20952 800 21072 0 FreeSans 480 0 0 0 access_write_mask_i[22]
port 46 nsew signal input
flabel metal3 s 0 21224 800 21344 0 FreeSans 480 0 0 0 access_write_mask_i[23]
port 47 nsew signal input
flabel metal3 s 0 21496 800 21616 0 FreeSans 480 0 0 0 access_write_mask_i[24]
port 48 nsew signal input
flabel metal3 s 0 21768 800 21888 0 FreeSans 480 0 0 0 access_write_mask_i[25]
port 49 nsew signal input
flabel metal3 s 0 22040 800 22160 0 FreeSans 480 0 0 0 access_write_mask_i[26]
port 50 nsew signal input
flabel metal3 s 0 22312 800 22432 0 FreeSans 480 0 0 0 access_write_mask_i[27]
port 51 nsew signal input
flabel metal3 s 0 22584 800 22704 0 FreeSans 480 0 0 0 access_write_mask_i[28]
port 52 nsew signal input
flabel metal3 s 0 22856 800 22976 0 FreeSans 480 0 0 0 access_write_mask_i[29]
port 53 nsew signal input
flabel metal3 s 0 15512 800 15632 0 FreeSans 480 0 0 0 access_write_mask_i[2]
port 54 nsew signal input
flabel metal3 s 0 23128 800 23248 0 FreeSans 480 0 0 0 access_write_mask_i[30]
port 55 nsew signal input
flabel metal3 s 0 23400 800 23520 0 FreeSans 480 0 0 0 access_write_mask_i[31]
port 56 nsew signal input
flabel metal3 s 0 15784 800 15904 0 FreeSans 480 0 0 0 access_write_mask_i[3]
port 57 nsew signal input
flabel metal3 s 0 16056 800 16176 0 FreeSans 480 0 0 0 access_write_mask_i[4]
port 58 nsew signal input
flabel metal3 s 0 16328 800 16448 0 FreeSans 480 0 0 0 access_write_mask_i[5]
port 59 nsew signal input
flabel metal3 s 0 16600 800 16720 0 FreeSans 480 0 0 0 access_write_mask_i[6]
port 60 nsew signal input
flabel metal3 s 0 16872 800 16992 0 FreeSans 480 0 0 0 access_write_mask_i[7]
port 61 nsew signal input
flabel metal3 s 0 17144 800 17264 0 FreeSans 480 0 0 0 access_write_mask_i[8]
port 62 nsew signal input
flabel metal3 s 0 17416 800 17536 0 FreeSans 480 0 0 0 access_write_mask_i[9]
port 63 nsew signal input
flabel metal3 s 29200 2184 30000 2304 0 FreeSans 480 0 0 0 reg_o[0]
port 64 nsew signal tristate
flabel metal3 s 29200 10344 30000 10464 0 FreeSans 480 0 0 0 reg_o[10]
port 65 nsew signal tristate
flabel metal3 s 29200 11160 30000 11280 0 FreeSans 480 0 0 0 reg_o[11]
port 66 nsew signal tristate
flabel metal3 s 29200 11976 30000 12096 0 FreeSans 480 0 0 0 reg_o[12]
port 67 nsew signal tristate
flabel metal3 s 29200 12792 30000 12912 0 FreeSans 480 0 0 0 reg_o[13]
port 68 nsew signal tristate
flabel metal3 s 29200 13608 30000 13728 0 FreeSans 480 0 0 0 reg_o[14]
port 69 nsew signal tristate
flabel metal3 s 29200 14424 30000 14544 0 FreeSans 480 0 0 0 reg_o[15]
port 70 nsew signal tristate
flabel metal3 s 29200 15240 30000 15360 0 FreeSans 480 0 0 0 reg_o[16]
port 71 nsew signal tristate
flabel metal3 s 29200 16056 30000 16176 0 FreeSans 480 0 0 0 reg_o[17]
port 72 nsew signal tristate
flabel metal3 s 29200 16872 30000 16992 0 FreeSans 480 0 0 0 reg_o[18]
port 73 nsew signal tristate
flabel metal3 s 29200 17688 30000 17808 0 FreeSans 480 0 0 0 reg_o[19]
port 74 nsew signal tristate
flabel metal3 s 29200 3000 30000 3120 0 FreeSans 480 0 0 0 reg_o[1]
port 75 nsew signal tristate
flabel metal3 s 29200 18504 30000 18624 0 FreeSans 480 0 0 0 reg_o[20]
port 76 nsew signal tristate
flabel metal3 s 29200 19320 30000 19440 0 FreeSans 480 0 0 0 reg_o[21]
port 77 nsew signal tristate
flabel metal3 s 29200 20136 30000 20256 0 FreeSans 480 0 0 0 reg_o[22]
port 78 nsew signal tristate
flabel metal3 s 29200 20952 30000 21072 0 FreeSans 480 0 0 0 reg_o[23]
port 79 nsew signal tristate
flabel metal3 s 29200 21768 30000 21888 0 FreeSans 480 0 0 0 reg_o[24]
port 80 nsew signal tristate
flabel metal3 s 29200 22584 30000 22704 0 FreeSans 480 0 0 0 reg_o[25]
port 81 nsew signal tristate
flabel metal3 s 29200 23400 30000 23520 0 FreeSans 480 0 0 0 reg_o[26]
port 82 nsew signal tristate
flabel metal3 s 29200 24216 30000 24336 0 FreeSans 480 0 0 0 reg_o[27]
port 83 nsew signal tristate
flabel metal3 s 29200 25032 30000 25152 0 FreeSans 480 0 0 0 reg_o[28]
port 84 nsew signal tristate
flabel metal3 s 29200 25848 30000 25968 0 FreeSans 480 0 0 0 reg_o[29]
port 85 nsew signal tristate
flabel metal3 s 29200 3816 30000 3936 0 FreeSans 480 0 0 0 reg_o[2]
port 86 nsew signal tristate
flabel metal3 s 29200 26664 30000 26784 0 FreeSans 480 0 0 0 reg_o[30]
port 87 nsew signal tristate
flabel metal3 s 29200 27480 30000 27600 0 FreeSans 480 0 0 0 reg_o[31]
port 88 nsew signal tristate
flabel metal3 s 29200 4632 30000 4752 0 FreeSans 480 0 0 0 reg_o[3]
port 89 nsew signal tristate
flabel metal3 s 29200 5448 30000 5568 0 FreeSans 480 0 0 0 reg_o[4]
port 90 nsew signal tristate
flabel metal3 s 29200 6264 30000 6384 0 FreeSans 480 0 0 0 reg_o[5]
port 91 nsew signal tristate
flabel metal3 s 29200 7080 30000 7200 0 FreeSans 480 0 0 0 reg_o[6]
port 92 nsew signal tristate
flabel metal3 s 29200 7896 30000 8016 0 FreeSans 480 0 0 0 reg_o[7]
port 93 nsew signal tristate
flabel metal3 s 29200 8712 30000 8832 0 FreeSans 480 0 0 0 reg_o[8]
port 94 nsew signal tristate
flabel metal3 s 29200 9528 30000 9648 0 FreeSans 480 0 0 0 reg_o[9]
port 95 nsew signal tristate
flabel metal4 s 4417 2128 4737 27792 0 FreeSans 1920 90 0 0 vccd1
port 96 nsew power bidirectional
flabel metal4 s 11363 2128 11683 27792 0 FreeSans 1920 90 0 0 vccd1
port 96 nsew power bidirectional
flabel metal4 s 18309 2128 18629 27792 0 FreeSans 1920 90 0 0 vccd1
port 96 nsew power bidirectional
flabel metal4 s 25255 2128 25575 27792 0 FreeSans 1920 90 0 0 vccd1
port 96 nsew power bidirectional
flabel metal4 s 7890 2128 8210 27792 0 FreeSans 1920 90 0 0 vssd1
port 97 nsew ground bidirectional
flabel metal4 s 14836 2128 15156 27792 0 FreeSans 1920 90 0 0 vssd1
port 97 nsew ground bidirectional
flabel metal4 s 21782 2128 22102 27792 0 FreeSans 1920 90 0 0 vssd1
port 97 nsew ground bidirectional
flabel metal4 s 28728 2128 29048 27792 0 FreeSans 1920 90 0 0 vssd1
port 97 nsew ground bidirectional
flabel metal2 s 478 0 534 800 0 FreeSans 224 90 0 0 wb_clk_i
port 98 nsew signal input
flabel metal2 s 754 0 810 800 0 FreeSans 224 90 0 0 wb_rst_i
port 99 nsew signal input
flabel metal2 s 20626 0 20682 800 0 FreeSans 224 90 0 0 wbs_ack_o
port 100 nsew signal tristate
flabel metal2 s 11794 0 11850 800 0 FreeSans 224 90 0 0 wbs_adr_i[0]
port 101 nsew signal input
flabel metal2 s 14554 0 14610 800 0 FreeSans 224 90 0 0 wbs_adr_i[10]
port 102 nsew signal input
flabel metal2 s 14830 0 14886 800 0 FreeSans 224 90 0 0 wbs_adr_i[11]
port 103 nsew signal input
flabel metal2 s 15106 0 15162 800 0 FreeSans 224 90 0 0 wbs_adr_i[12]
port 104 nsew signal input
flabel metal2 s 15382 0 15438 800 0 FreeSans 224 90 0 0 wbs_adr_i[13]
port 105 nsew signal input
flabel metal2 s 15658 0 15714 800 0 FreeSans 224 90 0 0 wbs_adr_i[14]
port 106 nsew signal input
flabel metal2 s 15934 0 15990 800 0 FreeSans 224 90 0 0 wbs_adr_i[15]
port 107 nsew signal input
flabel metal2 s 16210 0 16266 800 0 FreeSans 224 90 0 0 wbs_adr_i[16]
port 108 nsew signal input
flabel metal2 s 16486 0 16542 800 0 FreeSans 224 90 0 0 wbs_adr_i[17]
port 109 nsew signal input
flabel metal2 s 16762 0 16818 800 0 FreeSans 224 90 0 0 wbs_adr_i[18]
port 110 nsew signal input
flabel metal2 s 17038 0 17094 800 0 FreeSans 224 90 0 0 wbs_adr_i[19]
port 111 nsew signal input
flabel metal2 s 12070 0 12126 800 0 FreeSans 224 90 0 0 wbs_adr_i[1]
port 112 nsew signal input
flabel metal2 s 17314 0 17370 800 0 FreeSans 224 90 0 0 wbs_adr_i[20]
port 113 nsew signal input
flabel metal2 s 17590 0 17646 800 0 FreeSans 224 90 0 0 wbs_adr_i[21]
port 114 nsew signal input
flabel metal2 s 17866 0 17922 800 0 FreeSans 224 90 0 0 wbs_adr_i[22]
port 115 nsew signal input
flabel metal2 s 18142 0 18198 800 0 FreeSans 224 90 0 0 wbs_adr_i[23]
port 116 nsew signal input
flabel metal2 s 18418 0 18474 800 0 FreeSans 224 90 0 0 wbs_adr_i[24]
port 117 nsew signal input
flabel metal2 s 18694 0 18750 800 0 FreeSans 224 90 0 0 wbs_adr_i[25]
port 118 nsew signal input
flabel metal2 s 18970 0 19026 800 0 FreeSans 224 90 0 0 wbs_adr_i[26]
port 119 nsew signal input
flabel metal2 s 19246 0 19302 800 0 FreeSans 224 90 0 0 wbs_adr_i[27]
port 120 nsew signal input
flabel metal2 s 19522 0 19578 800 0 FreeSans 224 90 0 0 wbs_adr_i[28]
port 121 nsew signal input
flabel metal2 s 19798 0 19854 800 0 FreeSans 224 90 0 0 wbs_adr_i[29]
port 122 nsew signal input
flabel metal2 s 12346 0 12402 800 0 FreeSans 224 90 0 0 wbs_adr_i[2]
port 123 nsew signal input
flabel metal2 s 20074 0 20130 800 0 FreeSans 224 90 0 0 wbs_adr_i[30]
port 124 nsew signal input
flabel metal2 s 20350 0 20406 800 0 FreeSans 224 90 0 0 wbs_adr_i[31]
port 125 nsew signal input
flabel metal2 s 12622 0 12678 800 0 FreeSans 224 90 0 0 wbs_adr_i[3]
port 126 nsew signal input
flabel metal2 s 12898 0 12954 800 0 FreeSans 224 90 0 0 wbs_adr_i[4]
port 127 nsew signal input
flabel metal2 s 13174 0 13230 800 0 FreeSans 224 90 0 0 wbs_adr_i[5]
port 128 nsew signal input
flabel metal2 s 13450 0 13506 800 0 FreeSans 224 90 0 0 wbs_adr_i[6]
port 129 nsew signal input
flabel metal2 s 13726 0 13782 800 0 FreeSans 224 90 0 0 wbs_adr_i[7]
port 130 nsew signal input
flabel metal2 s 14002 0 14058 800 0 FreeSans 224 90 0 0 wbs_adr_i[8]
port 131 nsew signal input
flabel metal2 s 14278 0 14334 800 0 FreeSans 224 90 0 0 wbs_adr_i[9]
port 132 nsew signal input
flabel metal2 s 1306 0 1362 800 0 FreeSans 224 90 0 0 wbs_cyc_i
port 133 nsew signal input
flabel metal2 s 2962 0 3018 800 0 FreeSans 224 90 0 0 wbs_dat_i[0]
port 134 nsew signal input
flabel metal2 s 5722 0 5778 800 0 FreeSans 224 90 0 0 wbs_dat_i[10]
port 135 nsew signal input
flabel metal2 s 5998 0 6054 800 0 FreeSans 224 90 0 0 wbs_dat_i[11]
port 136 nsew signal input
flabel metal2 s 6274 0 6330 800 0 FreeSans 224 90 0 0 wbs_dat_i[12]
port 137 nsew signal input
flabel metal2 s 6550 0 6606 800 0 FreeSans 224 90 0 0 wbs_dat_i[13]
port 138 nsew signal input
flabel metal2 s 6826 0 6882 800 0 FreeSans 224 90 0 0 wbs_dat_i[14]
port 139 nsew signal input
flabel metal2 s 7102 0 7158 800 0 FreeSans 224 90 0 0 wbs_dat_i[15]
port 140 nsew signal input
flabel metal2 s 7378 0 7434 800 0 FreeSans 224 90 0 0 wbs_dat_i[16]
port 141 nsew signal input
flabel metal2 s 7654 0 7710 800 0 FreeSans 224 90 0 0 wbs_dat_i[17]
port 142 nsew signal input
flabel metal2 s 7930 0 7986 800 0 FreeSans 224 90 0 0 wbs_dat_i[18]
port 143 nsew signal input
flabel metal2 s 8206 0 8262 800 0 FreeSans 224 90 0 0 wbs_dat_i[19]
port 144 nsew signal input
flabel metal2 s 3238 0 3294 800 0 FreeSans 224 90 0 0 wbs_dat_i[1]
port 145 nsew signal input
flabel metal2 s 8482 0 8538 800 0 FreeSans 224 90 0 0 wbs_dat_i[20]
port 146 nsew signal input
flabel metal2 s 8758 0 8814 800 0 FreeSans 224 90 0 0 wbs_dat_i[21]
port 147 nsew signal input
flabel metal2 s 9034 0 9090 800 0 FreeSans 224 90 0 0 wbs_dat_i[22]
port 148 nsew signal input
flabel metal2 s 9310 0 9366 800 0 FreeSans 224 90 0 0 wbs_dat_i[23]
port 149 nsew signal input
flabel metal2 s 9586 0 9642 800 0 FreeSans 224 90 0 0 wbs_dat_i[24]
port 150 nsew signal input
flabel metal2 s 9862 0 9918 800 0 FreeSans 224 90 0 0 wbs_dat_i[25]
port 151 nsew signal input
flabel metal2 s 10138 0 10194 800 0 FreeSans 224 90 0 0 wbs_dat_i[26]
port 152 nsew signal input
flabel metal2 s 10414 0 10470 800 0 FreeSans 224 90 0 0 wbs_dat_i[27]
port 153 nsew signal input
flabel metal2 s 10690 0 10746 800 0 FreeSans 224 90 0 0 wbs_dat_i[28]
port 154 nsew signal input
flabel metal2 s 10966 0 11022 800 0 FreeSans 224 90 0 0 wbs_dat_i[29]
port 155 nsew signal input
flabel metal2 s 3514 0 3570 800 0 FreeSans 224 90 0 0 wbs_dat_i[2]
port 156 nsew signal input
flabel metal2 s 11242 0 11298 800 0 FreeSans 224 90 0 0 wbs_dat_i[30]
port 157 nsew signal input
flabel metal2 s 11518 0 11574 800 0 FreeSans 224 90 0 0 wbs_dat_i[31]
port 158 nsew signal input
flabel metal2 s 3790 0 3846 800 0 FreeSans 224 90 0 0 wbs_dat_i[3]
port 159 nsew signal input
flabel metal2 s 4066 0 4122 800 0 FreeSans 224 90 0 0 wbs_dat_i[4]
port 160 nsew signal input
flabel metal2 s 4342 0 4398 800 0 FreeSans 224 90 0 0 wbs_dat_i[5]
port 161 nsew signal input
flabel metal2 s 4618 0 4674 800 0 FreeSans 224 90 0 0 wbs_dat_i[6]
port 162 nsew signal input
flabel metal2 s 4894 0 4950 800 0 FreeSans 224 90 0 0 wbs_dat_i[7]
port 163 nsew signal input
flabel metal2 s 5170 0 5226 800 0 FreeSans 224 90 0 0 wbs_dat_i[8]
port 164 nsew signal input
flabel metal2 s 5446 0 5502 800 0 FreeSans 224 90 0 0 wbs_dat_i[9]
port 165 nsew signal input
flabel metal2 s 20902 0 20958 800 0 FreeSans 224 90 0 0 wbs_dat_o[0]
port 166 nsew signal tristate
flabel metal2 s 23662 0 23718 800 0 FreeSans 224 90 0 0 wbs_dat_o[10]
port 167 nsew signal tristate
flabel metal2 s 23938 0 23994 800 0 FreeSans 224 90 0 0 wbs_dat_o[11]
port 168 nsew signal tristate
flabel metal2 s 24214 0 24270 800 0 FreeSans 224 90 0 0 wbs_dat_o[12]
port 169 nsew signal tristate
flabel metal2 s 24490 0 24546 800 0 FreeSans 224 90 0 0 wbs_dat_o[13]
port 170 nsew signal tristate
flabel metal2 s 24766 0 24822 800 0 FreeSans 224 90 0 0 wbs_dat_o[14]
port 171 nsew signal tristate
flabel metal2 s 25042 0 25098 800 0 FreeSans 224 90 0 0 wbs_dat_o[15]
port 172 nsew signal tristate
flabel metal2 s 25318 0 25374 800 0 FreeSans 224 90 0 0 wbs_dat_o[16]
port 173 nsew signal tristate
flabel metal2 s 25594 0 25650 800 0 FreeSans 224 90 0 0 wbs_dat_o[17]
port 174 nsew signal tristate
flabel metal2 s 25870 0 25926 800 0 FreeSans 224 90 0 0 wbs_dat_o[18]
port 175 nsew signal tristate
flabel metal2 s 26146 0 26202 800 0 FreeSans 224 90 0 0 wbs_dat_o[19]
port 176 nsew signal tristate
flabel metal2 s 21178 0 21234 800 0 FreeSans 224 90 0 0 wbs_dat_o[1]
port 177 nsew signal tristate
flabel metal2 s 26422 0 26478 800 0 FreeSans 224 90 0 0 wbs_dat_o[20]
port 178 nsew signal tristate
flabel metal2 s 26698 0 26754 800 0 FreeSans 224 90 0 0 wbs_dat_o[21]
port 179 nsew signal tristate
flabel metal2 s 26974 0 27030 800 0 FreeSans 224 90 0 0 wbs_dat_o[22]
port 180 nsew signal tristate
flabel metal2 s 27250 0 27306 800 0 FreeSans 224 90 0 0 wbs_dat_o[23]
port 181 nsew signal tristate
flabel metal2 s 27526 0 27582 800 0 FreeSans 224 90 0 0 wbs_dat_o[24]
port 182 nsew signal tristate
flabel metal2 s 27802 0 27858 800 0 FreeSans 224 90 0 0 wbs_dat_o[25]
port 183 nsew signal tristate
flabel metal2 s 28078 0 28134 800 0 FreeSans 224 90 0 0 wbs_dat_o[26]
port 184 nsew signal tristate
flabel metal2 s 28354 0 28410 800 0 FreeSans 224 90 0 0 wbs_dat_o[27]
port 185 nsew signal tristate
flabel metal2 s 28630 0 28686 800 0 FreeSans 224 90 0 0 wbs_dat_o[28]
port 186 nsew signal tristate
flabel metal2 s 28906 0 28962 800 0 FreeSans 224 90 0 0 wbs_dat_o[29]
port 187 nsew signal tristate
flabel metal2 s 21454 0 21510 800 0 FreeSans 224 90 0 0 wbs_dat_o[2]
port 188 nsew signal tristate
flabel metal2 s 29182 0 29238 800 0 FreeSans 224 90 0 0 wbs_dat_o[30]
port 189 nsew signal tristate
flabel metal2 s 29458 0 29514 800 0 FreeSans 224 90 0 0 wbs_dat_o[31]
port 190 nsew signal tristate
flabel metal2 s 21730 0 21786 800 0 FreeSans 224 90 0 0 wbs_dat_o[3]
port 191 nsew signal tristate
flabel metal2 s 22006 0 22062 800 0 FreeSans 224 90 0 0 wbs_dat_o[4]
port 192 nsew signal tristate
flabel metal2 s 22282 0 22338 800 0 FreeSans 224 90 0 0 wbs_dat_o[5]
port 193 nsew signal tristate
flabel metal2 s 22558 0 22614 800 0 FreeSans 224 90 0 0 wbs_dat_o[6]
port 194 nsew signal tristate
flabel metal2 s 22834 0 22890 800 0 FreeSans 224 90 0 0 wbs_dat_o[7]
port 195 nsew signal tristate
flabel metal2 s 23110 0 23166 800 0 FreeSans 224 90 0 0 wbs_dat_o[8]
port 196 nsew signal tristate
flabel metal2 s 23386 0 23442 800 0 FreeSans 224 90 0 0 wbs_dat_o[9]
port 197 nsew signal tristate
flabel metal2 s 1858 0 1914 800 0 FreeSans 224 90 0 0 wbs_sel_i[0]
port 198 nsew signal input
flabel metal2 s 2134 0 2190 800 0 FreeSans 224 90 0 0 wbs_sel_i[1]
port 199 nsew signal input
flabel metal2 s 2410 0 2466 800 0 FreeSans 224 90 0 0 wbs_sel_i[2]
port 200 nsew signal input
flabel metal2 s 2686 0 2742 800 0 FreeSans 224 90 0 0 wbs_sel_i[3]
port 201 nsew signal input
flabel metal2 s 1030 0 1086 800 0 FreeSans 224 90 0 0 wbs_stb_i
port 202 nsew signal input
flabel metal2 s 1582 0 1638 800 0 FreeSans 224 90 0 0 wbs_we_i
port 203 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 30000 30000
<< end >>
