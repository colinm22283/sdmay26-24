// This is the unpowered netlist.
module spi_mem_m (clk_i,
    nrst_i,
    spi_clk_o,
    spi_cs_o,
    spi_dqsm_i,
    spi_dqsm_o,
    spi_miso_i,
    spi_mosi_o,
    sport_i,
    sport_o);
 input clk_i;
 input nrst_i;
 output spi_clk_o;
 output spi_cs_o;
 input spi_dqsm_i;
 output spi_dqsm_o;
 input [3:0] spi_miso_i;
 output [3:0] spi_mosi_o;
 input [56:0] sport_i;
 output [33:0] sport_o;

 wire net108;
 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire clknet_0_clk_i;
 wire clknet_3_0__leaf_clk_i;
 wire clknet_3_1__leaf_clk_i;
 wire clknet_3_2__leaf_clk_i;
 wire clknet_3_3__leaf_clk_i;
 wire clknet_3_4__leaf_clk_i;
 wire clknet_3_5__leaf_clk_i;
 wire clknet_3_6__leaf_clk_i;
 wire clknet_3_7__leaf_clk_i;
 wire clock_enable;
 wire current_dqsm;
 wire \current_nibble[0] ;
 wire \current_nibble[1] ;
 wire \current_nibble[2] ;
 wire \latency_count[0] ;
 wire \latency_count[1] ;
 wire \latency_count[2] ;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net15;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net16;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net17;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net18;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net19;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net2;
 wire net20;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net21;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net22;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net23;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net24;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net25;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net26;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net27;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net28;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net29;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net3;
 wire net30;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net31;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net32;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net33;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net34;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net35;
 wire net350;
 wire net351;
 wire net352;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net4;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net5;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net6;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net7;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net8;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire \pre_cycle[0] ;
 wire \pre_cycle[1] ;
 wire \read_buf[0] ;
 wire \read_buf[10] ;
 wire \read_buf[11] ;
 wire \read_buf[12] ;
 wire \read_buf[13] ;
 wire \read_buf[14] ;
 wire \read_buf[15] ;
 wire \read_buf[16] ;
 wire \read_buf[17] ;
 wire \read_buf[18] ;
 wire \read_buf[19] ;
 wire \read_buf[1] ;
 wire \read_buf[20] ;
 wire \read_buf[21] ;
 wire \read_buf[22] ;
 wire \read_buf[23] ;
 wire \read_buf[24] ;
 wire \read_buf[25] ;
 wire \read_buf[26] ;
 wire \read_buf[27] ;
 wire \read_buf[28] ;
 wire \read_buf[29] ;
 wire \read_buf[2] ;
 wire \read_buf[30] ;
 wire \read_buf[31] ;
 wire \read_buf[3] ;
 wire \read_buf[4] ;
 wire \read_buf[5] ;
 wire \read_buf[6] ;
 wire \read_buf[7] ;
 wire \read_buf[8] ;
 wire \read_buf[9] ;
 wire \read_byte[0] ;
 wire \read_byte[1] ;
 wire \read_byte[2] ;
 wire \read_word[0] ;
 wire \read_word[1] ;
 wire \read_word[2] ;
 wire \state[0] ;
 wire \state[10] ;
 wire \state[11] ;
 wire \state[1] ;
 wire \state[2] ;
 wire \state[3] ;
 wire \state[4] ;
 wire \state[5] ;
 wire \state[6] ;
 wire \state[7] ;
 wire \state[8] ;
 wire \state[9] ;
 wire word_ready;
 wire \write_buf[0] ;
 wire \write_buf[10] ;
 wire \write_buf[11] ;
 wire \write_buf[12] ;
 wire \write_buf[13] ;
 wire \write_buf[14] ;
 wire \write_buf[15] ;
 wire \write_buf[16] ;
 wire \write_buf[17] ;
 wire \write_buf[18] ;
 wire \write_buf[19] ;
 wire \write_buf[1] ;
 wire \write_buf[20] ;
 wire \write_buf[21] ;
 wire \write_buf[22] ;
 wire \write_buf[23] ;
 wire \write_buf[24] ;
 wire \write_buf[25] ;
 wire \write_buf[26] ;
 wire \write_buf[27] ;
 wire \write_buf[28] ;
 wire \write_buf[29] ;
 wire \write_buf[2] ;
 wire \write_buf[30] ;
 wire \write_buf[31] ;
 wire \write_buf[3] ;
 wire \write_buf[4] ;
 wire \write_buf[5] ;
 wire \write_buf[6] ;
 wire \write_buf[7] ;
 wire \write_buf[8] ;
 wire \write_buf[9] ;
 wire \write_byte[0] ;
 wire \write_byte[1] ;
 wire \write_byte[2] ;
 wire \write_word[0] ;
 wire \write_word[1] ;
 wire \write_word[2] ;

 sky130_fd_sc_hd__diode_2 ANTENNA__0783__B (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__0785__A (.DIODE(_0249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0789__A (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__0793__A (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__0797__A (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA__0801__A (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__0818__B (.DIODE(_0274_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0819__A (.DIODE(_0274_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0822__A (.DIODE(_0274_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0825__A (.DIODE(_0274_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0828__A (.DIODE(_0274_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0843__A (.DIODE(_0249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0848__C_N (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA__0855__A1 (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA__0857__A (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__0858__B (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__0863__B (.DIODE(_0310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0872__B (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__0872__C (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__0873__A (.DIODE(_0310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0875__A (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__0876__B (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__0878__A (.DIODE(_0325_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0884__A3 (.DIODE(_0326_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0887__A (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__0892__B (.DIODE(_0013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0895__A (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__0896__B (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__0898__B (.DIODE(_0341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0901__A (.DIODE(_0343_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0903__A (.DIODE(_0310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0913__B (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__0915__A2 (.DIODE(_0013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0917__A (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__0924__A (.DIODE(word_ready));
 sky130_fd_sc_hd__diode_2 ANTENNA__0925__A (.DIODE(_0325_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0926__A (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__0926__B (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__0926__C (.DIODE(_0274_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0927__A2 (.DIODE(_0364_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0936__A (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__0937__A (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__0938__A1 (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA__0945__A (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__0946__A (.DIODE(_0380_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0952__C (.DIODE(_0380_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0967__A (.DIODE(_0343_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0981__A (.DIODE(_0274_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0983__A (.DIODE(_0274_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0985__A (.DIODE(_0274_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0987__A (.DIODE(_0274_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1004__B1 (.DIODE(_0249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1005__B (.DIODE(_0249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1008__A (.DIODE(_0249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1014__1_A (.DIODE(clknet_3_1__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1015__A (.DIODE(_0341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1016__A (.DIODE(_0341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1017__A (.DIODE(_0341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1018__A (.DIODE(_0341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1019__A (.DIODE(_0341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1020__A (.DIODE(_0341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1021__A (.DIODE(_0341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1022__A (.DIODE(_0341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1023__A (.DIODE(_0341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1024__A (.DIODE(_0341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1025__A (.DIODE(_0341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1026__A (.DIODE(_0341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1027__A (.DIODE(_0341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1028__A (.DIODE(_0341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1029__A (.DIODE(_0341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1030__B (.DIODE(_0326_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1031__A2 (.DIODE(_0364_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1033__A (.DIODE(_0425_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1034__A (.DIODE(_0425_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1037__B (.DIODE(_0326_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1038__A2 (.DIODE(_0364_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1041__B (.DIODE(_0325_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1042__A2 (.DIODE(_0364_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1045__B (.DIODE(_0325_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1046__A2 (.DIODE(_0364_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1049__B (.DIODE(_0325_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1050__A2 (.DIODE(_0364_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1053__B (.DIODE(_0325_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1054__A2 (.DIODE(_0364_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1057__B (.DIODE(_0325_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1058__A2 (.DIODE(_0364_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1061__B (.DIODE(_0325_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1062__A2 (.DIODE(_0364_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1065__A (.DIODE(_0326_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1091__A (.DIODE(_0425_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1092__A (.DIODE(_0425_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1116__A (.DIODE(_0326_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1119__A (.DIODE(_0326_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1122__A (.DIODE(_0326_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1125__A (.DIODE(_0326_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1128__A (.DIODE(_0326_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1131__A (.DIODE(_0326_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1134__A (.DIODE(_0326_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1137__A (.DIODE(_0326_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1144__B1 (.DIODE(word_ready));
 sky130_fd_sc_hd__diode_2 ANTENNA__1154__A (.DIODE(_0310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1155__B (.DIODE(_0514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1165__B (.DIODE(_0514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1169__B (.DIODE(_0343_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1174__A (.DIODE(_0380_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1176__C (.DIODE(_0343_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1177__A (.DIODE(_0380_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1179__C (.DIODE(_0310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1187__B (.DIODE(_0514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1197__B (.DIODE(_0326_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1199__C1 (.DIODE(_0364_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1203__S (.DIODE(_0310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1204__C (.DIODE(_0310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1205__A (.DIODE(_0343_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1206__B (.DIODE(_0310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1212__B1 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__1222__B (.DIODE(_0514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1232__B (.DIODE(_0343_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1235__B (.DIODE(_0514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1244__B (.DIODE(_0514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1250__B (.DIODE(_0343_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1258__B (.DIODE(_0514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1264__B (.DIODE(_0343_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1270__B (.DIODE(_0326_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1272__C1 (.DIODE(_0364_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1275__S (.DIODE(_0310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1277__A (.DIODE(_0343_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1280__S (.DIODE(_0310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1283__A (.DIODE(_0514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1292__B (.DIODE(_0514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1296__B (.DIODE(_0343_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1302__B (.DIODE(_0514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1306__B (.DIODE(_0343_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1311__A (.DIODE(_0380_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1313__C (.DIODE(_0343_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1314__A (.DIODE(_0380_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1316__C (.DIODE(_0310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1323__B (.DIODE(_0514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1331__B (.DIODE(_0326_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1333__C1 (.DIODE(_0364_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1336__S (.DIODE(_0310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1338__A1 (.DIODE(_0343_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1349__B (.DIODE(_0514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1359__B (.DIODE(_0343_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1362__B (.DIODE(_0310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1371__B (.DIODE(_0514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1377__B (.DIODE(_0343_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1385__B (.DIODE(_0514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1389__C (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__1391__B (.DIODE(_0343_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1397__B (.DIODE(_0326_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1399__C1 (.DIODE(_0364_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1402__S (.DIODE(_0310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1404__S (.DIODE(_0310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1408__S (.DIODE(_0310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1411__A (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__1417__C (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__1496__B (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__1501__A1 (.DIODE(_0514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1502__A1 (.DIODE(_0514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1514__A (.DIODE(_0013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1517__A2 (.DIODE(_0013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1565__RESET_B (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__1566__CLK (.DIODE(clknet_3_3__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1568__CLK (.DIODE(clknet_3_1__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1568__RESET_B (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__1572__RESET_B (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__1573__RESET_B (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__1574__RESET_B (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__1582__CLK (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__1583__CLK (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__1584__CLK (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__1594__CLK (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__1595__CLK (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__1596__CLK (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__1597__RESET_B (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__1598__CLK (.DIODE(_0013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1617__CLK (.DIODE(clknet_3_1__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1618__CLK (.DIODE(clknet_3_1__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1621__CLK (.DIODE(clknet_3_1__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1631__CLK (.DIODE(clknet_3_3__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1641__CLK (.DIODE(clknet_3_3__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1642__CLK (.DIODE(clknet_3_3__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1645__CLK (.DIODE(clknet_3_3__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1646__CLK (.DIODE(clknet_3_3__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1683__RESET_B (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__1684__RESET_B (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__1685__CLK (.DIODE(clknet_3_3__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1685__RESET_B (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__1687__CLK (.DIODE(clknet_3_3__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1687__RESET_B (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__1688__CLK (.DIODE(clknet_3_1__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1688__RESET_B (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__1689__CLK (.DIODE(clknet_3_1__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1689__RESET_B (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__1690__CLK (.DIODE(clknet_3_1__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__1690__RESET_B (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__1693__RESET_B (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__1694__RESET_B (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__1695__RESET_B (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__1696__RESET_B (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_0__f_clk_i_A (.DIODE(clknet_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_1__f_clk_i_A (.DIODE(clknet_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_2__f_clk_i_A (.DIODE(clknet_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_3__f_clk_i_A (.DIODE(clknet_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_4__f_clk_i_A (.DIODE(clknet_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_5__f_clk_i_A (.DIODE(clknet_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_6__f_clk_i_A (.DIODE(clknet_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_7__f_clk_i_A (.DIODE(clknet_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout103_A (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout104_A (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout105_A (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout106_A (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout107_A (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold156_A (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold215_A (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold234_A (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold241_A (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold85_A (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold88_A (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_output63_A (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA_output64_A (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA_output65_A (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA_output66_A (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA_output68_A (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_output93_A (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA_output94_A (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA_output95_A (.DIODE(net95));
 sky130_fd_sc_hd__decap_8 FILLER_0_0_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_43 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_43 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_550 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_485 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_555 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_604 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_620 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_51 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_515 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_552 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_580 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_588 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_518 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_555 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_605 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_43 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_534 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_579 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_605 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_520 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_557 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_586 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_593 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_500 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_525 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_569 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_94 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_511 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_575 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_579 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_58 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_621 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_56 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_560 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_564 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_68 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_88 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_516 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_566 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_570 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_583 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_591 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_621 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_620 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_91 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_592 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_35 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_43 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_546 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_564 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_574 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_32 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_497 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_579 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_602 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_43 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_480 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_550 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_562 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_582 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_96 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_457 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_466 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_543 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_78 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_96 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_11 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_472 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_499 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_506 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_512 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_569 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_610 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_40 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_590 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_602 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_80 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_84 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_124 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_415 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_504 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_511 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_564 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_568 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_409 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_472 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_552 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_564 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_572 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_588 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_92 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_508 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_537 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_551 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_60 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_600 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_623 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_76 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_127 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_399 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_46 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_570 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_574 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_602 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_35 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_385 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_424 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_512 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_623 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_91 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_435 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_479 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_48 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_483 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_588 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_70 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_84 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_98 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_450 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_454 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_471 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_483 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_510 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_58 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_624 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_403 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_452 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_468 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_523 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_572 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_582 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_598 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_86 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_397 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_428 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_440 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_491 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_507 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_560 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_564 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_592 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_72 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_442 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_468 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_534 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_63 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_127 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_504 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_508 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_547 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_420 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_52 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_532 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_603 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_613 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_114 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_40 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_450 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_460 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_52 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_610 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_95 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_516 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_73 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_178 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_43 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_462 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_570 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_61 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_67 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_71 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_91 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_36 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_385 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_427 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_46 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_492 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_500 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_514 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_523 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_586 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_86 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_94 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_100 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_406 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_440 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_515 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_534 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_606 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_504 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_547 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_606 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_66 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_532 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_620 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_43 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_481 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_491 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_506 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_40 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_596 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_43 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_38 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_58 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_620 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_189 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_46 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_40 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_624 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_49 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_624 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_28 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_40 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_43 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_618 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_43 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_43 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_43 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_93 ();
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_148 ();
 sky130_fd_sc_hd__decap_3 PHY_149 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_150 ();
 sky130_fd_sc_hd__decap_3 PHY_151 ();
 sky130_fd_sc_hd__decap_3 PHY_152 ();
 sky130_fd_sc_hd__decap_3 PHY_153 ();
 sky130_fd_sc_hd__decap_3 PHY_154 ();
 sky130_fd_sc_hd__decap_3 PHY_155 ();
 sky130_fd_sc_hd__decap_3 PHY_156 ();
 sky130_fd_sc_hd__decap_3 PHY_157 ();
 sky130_fd_sc_hd__decap_3 PHY_158 ();
 sky130_fd_sc_hd__decap_3 PHY_159 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_160 ();
 sky130_fd_sc_hd__decap_3 PHY_161 ();
 sky130_fd_sc_hd__decap_3 PHY_162 ();
 sky130_fd_sc_hd__decap_3 PHY_163 ();
 sky130_fd_sc_hd__decap_3 PHY_164 ();
 sky130_fd_sc_hd__decap_3 PHY_165 ();
 sky130_fd_sc_hd__decap_3 PHY_166 ();
 sky130_fd_sc_hd__decap_3 PHY_167 ();
 sky130_fd_sc_hd__decap_3 PHY_168 ();
 sky130_fd_sc_hd__decap_3 PHY_169 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_170 ();
 sky130_fd_sc_hd__decap_3 PHY_171 ();
 sky130_fd_sc_hd__decap_3 PHY_172 ();
 sky130_fd_sc_hd__decap_3 PHY_173 ();
 sky130_fd_sc_hd__decap_3 PHY_174 ();
 sky130_fd_sc_hd__decap_3 PHY_175 ();
 sky130_fd_sc_hd__decap_3 PHY_176 ();
 sky130_fd_sc_hd__decap_3 PHY_177 ();
 sky130_fd_sc_hd__decap_3 PHY_178 ();
 sky130_fd_sc_hd__decap_3 PHY_179 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_180 ();
 sky130_fd_sc_hd__decap_3 PHY_181 ();
 sky130_fd_sc_hd__decap_3 PHY_182 ();
 sky130_fd_sc_hd__decap_3 PHY_183 ();
 sky130_fd_sc_hd__decap_3 PHY_184 ();
 sky130_fd_sc_hd__decap_3 PHY_185 ();
 sky130_fd_sc_hd__decap_3 PHY_186 ();
 sky130_fd_sc_hd__decap_3 PHY_187 ();
 sky130_fd_sc_hd__decap_3 PHY_188 ();
 sky130_fd_sc_hd__decap_3 PHY_189 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_190 ();
 sky130_fd_sc_hd__decap_3 PHY_191 ();
 sky130_fd_sc_hd__decap_3 PHY_192 ();
 sky130_fd_sc_hd__decap_3 PHY_193 ();
 sky130_fd_sc_hd__decap_3 PHY_194 ();
 sky130_fd_sc_hd__decap_3 PHY_195 ();
 sky130_fd_sc_hd__decap_3 PHY_196 ();
 sky130_fd_sc_hd__decap_3 PHY_197 ();
 sky130_fd_sc_hd__decap_3 PHY_198 ();
 sky130_fd_sc_hd__decap_3 PHY_199 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_200 ();
 sky130_fd_sc_hd__decap_3 PHY_201 ();
 sky130_fd_sc_hd__decap_3 PHY_202 ();
 sky130_fd_sc_hd__decap_3 PHY_203 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_999 ();
 sky130_fd_sc_hd__nand2_1 _0779_ (.A(\read_byte[1] ),
    .B(\read_byte[0] ),
    .Y(_0244_));
 sky130_fd_sc_hd__nor2_1 _0780_ (.A(\read_byte[2] ),
    .B(_0244_),
    .Y(_0245_));
 sky130_fd_sc_hd__inv_2 _0781_ (.A(_0245_),
    .Y(_0246_));
 sky130_fd_sc_hd__nand2_1 _0782_ (.A(_0246_),
    .B(\read_buf[31] ),
    .Y(_0247_));
 sky130_fd_sc_hd__nand2_1 _0783_ (.A(_0245_),
    .B(net6),
    .Y(_0248_));
 sky130_fd_sc_hd__nor2_2 _0784_ (.A(\state[1] ),
    .B(\state[11] ),
    .Y(_0249_));
 sky130_fd_sc_hd__buf_4 _0785_ (.A(_0249_),
    .X(_0250_));
 sky130_fd_sc_hd__a21oi_1 _0786_ (.A1(_0247_),
    .A2(_0248_),
    .B1(_0250_),
    .Y(_0069_));
 sky130_fd_sc_hd__inv_2 _0787_ (.A(\read_byte[1] ),
    .Y(_0251_));
 sky130_fd_sc_hd__inv_2 _0788_ (.A(\read_byte[0] ),
    .Y(_0252_));
 sky130_fd_sc_hd__inv_2 _0789_ (.A(net5),
    .Y(_0253_));
 sky130_fd_sc_hd__or4_1 _0790_ (.A(\read_byte[2] ),
    .B(_0251_),
    .C(_0252_),
    .D(_0253_),
    .X(_0254_));
 sky130_fd_sc_hd__nand2_1 _0791_ (.A(_0246_),
    .B(\read_buf[30] ),
    .Y(_0255_));
 sky130_fd_sc_hd__a21oi_1 _0792_ (.A1(_0254_),
    .A2(_0255_),
    .B1(_0250_),
    .Y(_0068_));
 sky130_fd_sc_hd__inv_2 _0793_ (.A(net4),
    .Y(_0256_));
 sky130_fd_sc_hd__or4_1 _0794_ (.A(\read_byte[2] ),
    .B(_0251_),
    .C(_0252_),
    .D(_0256_),
    .X(_0257_));
 sky130_fd_sc_hd__nand2_1 _0795_ (.A(_0246_),
    .B(\read_buf[29] ),
    .Y(_0258_));
 sky130_fd_sc_hd__a21oi_1 _0796_ (.A1(_0257_),
    .A2(_0258_),
    .B1(_0250_),
    .Y(_0067_));
 sky130_fd_sc_hd__inv_2 _0797_ (.A(net3),
    .Y(_0259_));
 sky130_fd_sc_hd__or4_1 _0798_ (.A(\read_byte[2] ),
    .B(_0251_),
    .C(_0252_),
    .D(_0259_),
    .X(_0260_));
 sky130_fd_sc_hd__nand2_1 _0799_ (.A(_0246_),
    .B(\read_buf[28] ),
    .Y(_0261_));
 sky130_fd_sc_hd__a21oi_1 _0800_ (.A1(_0260_),
    .A2(_0261_),
    .B1(_0250_),
    .Y(_0066_));
 sky130_fd_sc_hd__inv_2 _0801_ (.A(net6),
    .Y(_0262_));
 sky130_fd_sc_hd__or3_1 _0802_ (.A(\read_byte[0] ),
    .B(\read_byte[2] ),
    .C(_0251_),
    .X(_0263_));
 sky130_fd_sc_hd__clkbuf_4 _0803_ (.A(_0263_),
    .X(_0264_));
 sky130_fd_sc_hd__or2_1 _0804_ (.A(_0262_),
    .B(_0264_),
    .X(_0265_));
 sky130_fd_sc_hd__nand2_1 _0805_ (.A(_0264_),
    .B(\read_buf[23] ),
    .Y(_0266_));
 sky130_fd_sc_hd__a21oi_1 _0806_ (.A1(_0265_),
    .A2(_0266_),
    .B1(_0250_),
    .Y(_0065_));
 sky130_fd_sc_hd__or2_1 _0807_ (.A(_0253_),
    .B(_0264_),
    .X(_0267_));
 sky130_fd_sc_hd__nand2_1 _0808_ (.A(_0264_),
    .B(\read_buf[22] ),
    .Y(_0268_));
 sky130_fd_sc_hd__a21oi_1 _0809_ (.A1(_0267_),
    .A2(_0268_),
    .B1(_0250_),
    .Y(_0064_));
 sky130_fd_sc_hd__or2_1 _0810_ (.A(_0256_),
    .B(_0264_),
    .X(_0269_));
 sky130_fd_sc_hd__nand2_1 _0811_ (.A(_0264_),
    .B(\read_buf[21] ),
    .Y(_0270_));
 sky130_fd_sc_hd__a21oi_1 _0812_ (.A1(_0269_),
    .A2(_0270_),
    .B1(_0250_),
    .Y(_0063_));
 sky130_fd_sc_hd__or2_1 _0813_ (.A(_0259_),
    .B(_0264_),
    .X(_0271_));
 sky130_fd_sc_hd__nand2_1 _0814_ (.A(_0264_),
    .B(\read_buf[20] ),
    .Y(_0272_));
 sky130_fd_sc_hd__a21oi_1 _0815_ (.A1(_0271_),
    .A2(_0272_),
    .B1(_0250_),
    .Y(_0062_));
 sky130_fd_sc_hd__or3_1 _0816_ (.A(\read_byte[1] ),
    .B(\read_byte[2] ),
    .C(_0252_),
    .X(_0273_));
 sky130_fd_sc_hd__buf_6 _0817_ (.A(_0273_),
    .X(_0274_));
 sky130_fd_sc_hd__or2_1 _0818_ (.A(_0262_),
    .B(_0274_),
    .X(_0275_));
 sky130_fd_sc_hd__nand2_1 _0819_ (.A(_0274_),
    .B(\read_buf[15] ),
    .Y(_0276_));
 sky130_fd_sc_hd__a21oi_1 _0820_ (.A1(_0275_),
    .A2(_0276_),
    .B1(_0250_),
    .Y(_0061_));
 sky130_fd_sc_hd__or4_1 _0821_ (.A(\read_byte[1] ),
    .B(\read_byte[2] ),
    .C(_0252_),
    .D(_0253_),
    .X(_0277_));
 sky130_fd_sc_hd__nand2_1 _0822_ (.A(_0274_),
    .B(\read_buf[14] ),
    .Y(_0278_));
 sky130_fd_sc_hd__a21oi_1 _0823_ (.A1(_0277_),
    .A2(_0278_),
    .B1(_0250_),
    .Y(_0060_));
 sky130_fd_sc_hd__or4_1 _0824_ (.A(\read_byte[1] ),
    .B(\read_byte[2] ),
    .C(_0252_),
    .D(_0256_),
    .X(_0279_));
 sky130_fd_sc_hd__nand2_1 _0825_ (.A(_0274_),
    .B(\read_buf[13] ),
    .Y(_0280_));
 sky130_fd_sc_hd__a21oi_1 _0826_ (.A1(_0279_),
    .A2(_0280_),
    .B1(_0250_),
    .Y(_0059_));
 sky130_fd_sc_hd__or4_1 _0827_ (.A(\read_byte[1] ),
    .B(\read_byte[2] ),
    .C(_0252_),
    .D(_0259_),
    .X(_0281_));
 sky130_fd_sc_hd__nand2_1 _0828_ (.A(_0274_),
    .B(\read_buf[12] ),
    .Y(_0282_));
 sky130_fd_sc_hd__a21oi_1 _0829_ (.A1(_0281_),
    .A2(_0282_),
    .B1(_0250_),
    .Y(_0058_));
 sky130_fd_sc_hd__or3_1 _0830_ (.A(\read_byte[1] ),
    .B(\read_byte[0] ),
    .C(\read_byte[2] ),
    .X(_0283_));
 sky130_fd_sc_hd__buf_2 _0831_ (.A(_0283_),
    .X(_0284_));
 sky130_fd_sc_hd__or2_1 _0832_ (.A(_0262_),
    .B(_0284_),
    .X(_0285_));
 sky130_fd_sc_hd__nand2_1 _0833_ (.A(_0284_),
    .B(\read_buf[7] ),
    .Y(_0286_));
 sky130_fd_sc_hd__a21oi_1 _0834_ (.A1(_0285_),
    .A2(_0286_),
    .B1(_0250_),
    .Y(_0057_));
 sky130_fd_sc_hd__or2_1 _0835_ (.A(_0253_),
    .B(_0284_),
    .X(_0287_));
 sky130_fd_sc_hd__nand2_1 _0836_ (.A(_0284_),
    .B(\read_buf[6] ),
    .Y(_0288_));
 sky130_fd_sc_hd__a21oi_1 _0837_ (.A1(_0287_),
    .A2(_0288_),
    .B1(_0250_),
    .Y(_0056_));
 sky130_fd_sc_hd__or2_1 _0838_ (.A(_0256_),
    .B(_0284_),
    .X(_0289_));
 sky130_fd_sc_hd__nand2_1 _0839_ (.A(_0284_),
    .B(\read_buf[5] ),
    .Y(_0290_));
 sky130_fd_sc_hd__a21oi_1 _0840_ (.A1(_0289_),
    .A2(_0290_),
    .B1(_0250_),
    .Y(_0055_));
 sky130_fd_sc_hd__or2_1 _0841_ (.A(_0259_),
    .B(_0284_),
    .X(_0291_));
 sky130_fd_sc_hd__nand2_1 _0842_ (.A(_0284_),
    .B(\read_buf[4] ),
    .Y(_0292_));
 sky130_fd_sc_hd__buf_4 _0843_ (.A(_0249_),
    .X(_0293_));
 sky130_fd_sc_hd__a21oi_1 _0844_ (.A1(_0291_),
    .A2(_0292_),
    .B1(_0293_),
    .Y(_0054_));
 sky130_fd_sc_hd__inv_2 _0845_ (.A(\state[9] ),
    .Y(_0294_));
 sky130_fd_sc_hd__or4_1 _0846_ (.A(net50),
    .B(net49),
    .C(net53),
    .D(net52),
    .X(_0295_));
 sky130_fd_sc_hd__or2_1 _0847_ (.A(net39),
    .B(net38),
    .X(_0296_));
 sky130_fd_sc_hd__or3b_1 _0848_ (.A(net37),
    .B(_0296_),
    .C_N(net54),
    .X(_0297_));
 sky130_fd_sc_hd__or4_1 _0849_ (.A(net46),
    .B(net45),
    .C(net48),
    .D(net47),
    .X(_0298_));
 sky130_fd_sc_hd__nor2_1 _0850_ (.A(_0297_),
    .B(_0298_),
    .Y(_0299_));
 sky130_fd_sc_hd__or2_1 _0851_ (.A(net41),
    .B(net42),
    .X(_0300_));
 sky130_fd_sc_hd__nor3_1 _0852_ (.A(net44),
    .B(net43),
    .C(_0300_),
    .Y(_0301_));
 sky130_fd_sc_hd__nand3b_2 _0853_ (.A_N(_0295_),
    .B(_0299_),
    .C(_0301_),
    .Y(_0302_));
 sky130_fd_sc_hd__nand2_1 _0854_ (.A(_0302_),
    .B(net203),
    .Y(_0303_));
 sky130_fd_sc_hd__o21ai_1 _0855_ (.A1(net54),
    .A2(_0294_),
    .B1(_0303_),
    .Y(_0003_));
 sky130_fd_sc_hd__inv_2 _0856_ (.A(net339),
    .Y(_0304_));
 sky130_fd_sc_hd__inv_2 _0857_ (.A(net55),
    .Y(_0305_));
 sky130_fd_sc_hd__nand2_2 _0858_ (.A(_0305_),
    .B(net56),
    .Y(_0306_));
 sky130_fd_sc_hd__buf_6 _0859_ (.A(_0306_),
    .X(_0307_));
 sky130_fd_sc_hd__nand2_1 _0860_ (.A(net332),
    .B(net329),
    .Y(_0308_));
 sky130_fd_sc_hd__nor2_1 _0861_ (.A(net214),
    .B(_0308_),
    .Y(_0309_));
 sky130_fd_sc_hd__clkbuf_8 _0862_ (.A(net342),
    .X(_0310_));
 sky130_fd_sc_hd__nand2_1 _0863_ (.A(_0309_),
    .B(_0310_),
    .Y(_0311_));
 sky130_fd_sc_hd__or3_2 _0864_ (.A(_0304_),
    .B(_0307_),
    .C(_0311_),
    .X(_0312_));
 sky130_fd_sc_hd__inv_2 _0865_ (.A(_0312_),
    .Y(_0313_));
 sky130_fd_sc_hd__or3b_1 _0866_ (.A(net335),
    .B(net205),
    .C_N(net200),
    .X(_0314_));
 sky130_fd_sc_hd__nor2_1 _0867_ (.A(net186),
    .B(net208),
    .Y(_0315_));
 sky130_fd_sc_hd__inv_2 _0868_ (.A(_0315_),
    .Y(_0316_));
 sky130_fd_sc_hd__nor2_1 _0869_ (.A(net189),
    .B(_0316_),
    .Y(_0317_));
 sky130_fd_sc_hd__nand2_1 _0870_ (.A(_0317_),
    .B(net349),
    .Y(_0318_));
 sky130_fd_sc_hd__inv_2 _0871_ (.A(_0318_),
    .Y(_0319_));
 sky130_fd_sc_hd__and3_1 _0872_ (.A(_0319_),
    .B(net63),
    .C(net57),
    .X(_0320_));
 sky130_fd_sc_hd__inv_2 _0873_ (.A(_0310_),
    .Y(_0321_));
 sky130_fd_sc_hd__nor2_1 _0874_ (.A(_0321_),
    .B(_0309_),
    .Y(_0322_));
 sky130_fd_sc_hd__inv_2 _0875_ (.A(net56),
    .Y(_0323_));
 sky130_fd_sc_hd__nand2_2 _0876_ (.A(_0323_),
    .B(net55),
    .Y(_0324_));
 sky130_fd_sc_hd__nand2_4 _0877_ (.A(_0306_),
    .B(_0324_),
    .Y(_0325_));
 sky130_fd_sc_hd__clkbuf_8 _0878_ (.A(_0325_),
    .X(_0326_));
 sky130_fd_sc_hd__nand2_1 _0879_ (.A(_0306_),
    .B(net339),
    .Y(_0327_));
 sky130_fd_sc_hd__nor2_1 _0880_ (.A(_0323_),
    .B(_0327_),
    .Y(_0328_));
 sky130_fd_sc_hd__inv_2 _0881_ (.A(_0328_),
    .Y(_0329_));
 sky130_fd_sc_hd__nand2_1 _0882_ (.A(_0321_),
    .B(net339),
    .Y(_0330_));
 sky130_fd_sc_hd__nand2_1 _0883_ (.A(_0329_),
    .B(_0330_),
    .Y(_0331_));
 sky130_fd_sc_hd__a31o_1 _0884_ (.A1(net339),
    .A2(_0322_),
    .A3(_0326_),
    .B1(_0331_),
    .X(_0332_));
 sky130_fd_sc_hd__a211o_1 _0885_ (.A1(_0313_),
    .A2(_0314_),
    .B1(_0320_),
    .C1(net340),
    .X(_0007_));
 sky130_fd_sc_hd__nor2_4 _0886_ (.A(\state[0] ),
    .B(\state[9] ),
    .Y(net94));
 sky130_fd_sc_hd__inv_2 _0887_ (.A(net94),
    .Y(net64));
 sky130_fd_sc_hd__inv_2 _0888_ (.A(net286),
    .Y(_0333_));
 sky130_fd_sc_hd__inv_2 _0889_ (.A(net327),
    .Y(_0334_));
 sky130_fd_sc_hd__nand2_1 _0890_ (.A(_0334_),
    .B(net192),
    .Y(_0335_));
 sky130_fd_sc_hd__inv_2 _0891_ (.A(net103),
    .Y(_0013_));
 sky130_fd_sc_hd__nor2_1 _0892_ (.A(net177),
    .B(_0013_),
    .Y(_0336_));
 sky130_fd_sc_hd__inv_2 _0893_ (.A(_0336_),
    .Y(_0337_));
 sky130_fd_sc_hd__nor2_1 _0894_ (.A(_0335_),
    .B(_0337_),
    .Y(_0338_));
 sky130_fd_sc_hd__inv_2 _0895_ (.A(net57),
    .Y(_0339_));
 sky130_fd_sc_hd__and3_1 _0896_ (.A(_0319_),
    .B(net63),
    .C(_0339_),
    .X(_0340_));
 sky130_fd_sc_hd__buf_8 _0897_ (.A(net103),
    .X(_0341_));
 sky130_fd_sc_hd__nand2_1 _0898_ (.A(_0340_),
    .B(_0341_),
    .Y(_0342_));
 sky130_fd_sc_hd__o21ai_1 _0899_ (.A1(_0333_),
    .A2(_0338_),
    .B1(_0342_),
    .Y(_0008_));
 sky130_fd_sc_hd__buf_6 _0900_ (.A(_0321_),
    .X(_0343_));
 sky130_fd_sc_hd__buf_4 _0901_ (.A(_0343_),
    .X(_0344_));
 sky130_fd_sc_hd__inv_2 _0902_ (.A(net183),
    .Y(_0345_));
 sky130_fd_sc_hd__nand2_1 _0903_ (.A(_0310_),
    .B(net319),
    .Y(_0346_));
 sky130_fd_sc_hd__inv_2 _0904_ (.A(_0346_),
    .Y(_0347_));
 sky130_fd_sc_hd__nand2_1 _0905_ (.A(_0347_),
    .B(net220),
    .Y(_0348_));
 sky130_fd_sc_hd__nand2_1 _0906_ (.A(_0348_),
    .B(\state[2] ),
    .Y(_0349_));
 sky130_fd_sc_hd__o21ai_1 _0907_ (.A1(_0344_),
    .A2(net184),
    .B1(_0349_),
    .Y(_0004_));
 sky130_fd_sc_hd__inv_2 _0908_ (.A(net348),
    .Y(_0350_));
 sky130_fd_sc_hd__nor2_1 _0909_ (.A(_0350_),
    .B(_0348_),
    .Y(_0351_));
 sky130_fd_sc_hd__inv_2 _0910_ (.A(_0317_),
    .Y(_0352_));
 sky130_fd_sc_hd__nand2_1 _0911_ (.A(_0352_),
    .B(net349),
    .Y(_0353_));
 sky130_fd_sc_hd__inv_2 _0912_ (.A(_0353_),
    .Y(_0354_));
 sky130_fd_sc_hd__nand2_1 _0913_ (.A(_0354_),
    .B(net63),
    .Y(_0355_));
 sky130_fd_sc_hd__inv_2 _0914_ (.A(_0355_),
    .Y(_0356_));
 sky130_fd_sc_hd__a21oi_1 _0915_ (.A1(_0340_),
    .A2(_0013_),
    .B1(_0356_),
    .Y(_0357_));
 sky130_fd_sc_hd__inv_2 _0916_ (.A(net349),
    .Y(_0358_));
 sky130_fd_sc_hd__nor2_1 _0917_ (.A(net63),
    .B(_0358_),
    .Y(_0359_));
 sky130_fd_sc_hd__inv_2 _0918_ (.A(_0359_),
    .Y(_0360_));
 sky130_fd_sc_hd__nand3b_1 _0919_ (.A_N(_0351_),
    .B(_0357_),
    .C(_0360_),
    .Y(_0010_));
 sky130_fd_sc_hd__or2_1 _0920_ (.A(_0314_),
    .B(_0312_),
    .X(_0361_));
 sky130_fd_sc_hd__o31ai_1 _0921_ (.A1(_0304_),
    .A2(_0311_),
    .A3(_0324_),
    .B1(_0361_),
    .Y(_0005_));
 sky130_fd_sc_hd__a21o_1 _0922_ (.A1(_0344_),
    .A2(net183),
    .B1(net110),
    .X(_0006_));
 sky130_fd_sc_hd__inv_2 _0923_ (.A(net337),
    .Y(_0362_));
 sky130_fd_sc_hd__inv_2 _0924_ (.A(word_ready),
    .Y(_0363_));
 sky130_fd_sc_hd__inv_4 _0925_ (.A(_0325_),
    .Y(_0364_));
 sky130_fd_sc_hd__or3_1 _0926_ (.A(net55),
    .B(net56),
    .C(_0274_),
    .X(_0365_));
 sky130_fd_sc_hd__o21ai_2 _0927_ (.A1(_0363_),
    .A2(_0364_),
    .B1(_0365_),
    .Y(_0366_));
 sky130_fd_sc_hd__inv_2 _0928_ (.A(net242),
    .Y(_0367_));
 sky130_fd_sc_hd__o31ai_2 _0929_ (.A1(net228),
    .A2(net345),
    .A3(_0367_),
    .B1(\state[1] ),
    .Y(_0368_));
 sky130_fd_sc_hd__nand2_1 _0930_ (.A(_0338_),
    .B(net286),
    .Y(_0369_));
 sky130_fd_sc_hd__o211ai_1 _0931_ (.A1(_0362_),
    .A2(_0366_),
    .B1(_0368_),
    .C1(net287),
    .Y(_0009_));
 sky130_fd_sc_hd__or2_1 _0932_ (.A(_0363_),
    .B(_0324_),
    .X(_0370_));
 sky130_fd_sc_hd__a21o_1 _0933_ (.A1(_0365_),
    .A2(_0370_),
    .B1(_0362_),
    .X(_0371_));
 sky130_fd_sc_hd__inv_2 _0934_ (.A(\state[1] ),
    .Y(_0372_));
 sky130_fd_sc_hd__or4_1 _0935_ (.A(net228),
    .B(\read_word[0] ),
    .C(_0372_),
    .D(_0367_),
    .X(_0373_));
 sky130_fd_sc_hd__buf_4 _0936_ (.A(net56),
    .X(_0374_));
 sky130_fd_sc_hd__or4_1 _0937_ (.A(net55),
    .B(_0374_),
    .C(_0304_),
    .D(_0344_),
    .X(_0375_));
 sky130_fd_sc_hd__a21oi_1 _0938_ (.A1(net54),
    .A2(\state[9] ),
    .B1(net180),
    .Y(_0376_));
 sky130_fd_sc_hd__and3_1 _0939_ (.A(_0373_),
    .B(_0375_),
    .C(_0376_),
    .X(_0377_));
 sky130_fd_sc_hd__nand2_1 _0940_ (.A(_0371_),
    .B(_0377_),
    .Y(_0011_));
 sky130_fd_sc_hd__and2b_1 _0941_ (.A_N(net350),
    .B(clock_enable),
    .X(_0378_));
 sky130_fd_sc_hd__clkbuf_1 _0942_ (.A(_0378_),
    .X(_0000_));
 sky130_fd_sc_hd__inv_2 _0943_ (.A(net203),
    .Y(_0379_));
 sky130_fd_sc_hd__nor2_1 _0944_ (.A(_0379_),
    .B(_0302_),
    .Y(_0002_));
 sky130_fd_sc_hd__nor2_2 _0945_ (.A(net55),
    .B(_0323_),
    .Y(_0380_));
 sky130_fd_sc_hd__nand2_1 _0946_ (.A(_0380_),
    .B(net337),
    .Y(_0381_));
 sky130_fd_sc_hd__nor2_1 _0947_ (.A(_0363_),
    .B(_0381_),
    .Y(_0001_));
 sky130_fd_sc_hd__inv_2 _0948_ (.A(net335),
    .Y(_0382_));
 sky130_fd_sc_hd__nor2_1 _0949_ (.A(_0306_),
    .B(_0330_),
    .Y(_0383_));
 sky130_fd_sc_hd__a21oi_1 _0950_ (.A1(_0379_),
    .A2(_0304_),
    .B1(_0383_),
    .Y(_0384_));
 sky130_fd_sc_hd__inv_2 _0951_ (.A(_0327_),
    .Y(_0385_));
 sky130_fd_sc_hd__and3_1 _0952_ (.A(_0322_),
    .B(\state[5] ),
    .C(_0380_),
    .X(_0386_));
 sky130_fd_sc_hd__nor2_1 _0953_ (.A(_0385_),
    .B(_0386_),
    .Y(_0387_));
 sky130_fd_sc_hd__nand3_2 _0954_ (.A(_0361_),
    .B(_0384_),
    .C(_0387_),
    .Y(_0388_));
 sky130_fd_sc_hd__a21o_1 _0955_ (.A1(_0313_),
    .A2(_0314_),
    .B1(net335),
    .X(_0389_));
 sky130_fd_sc_hd__o21a_1 _0956_ (.A1(_0382_),
    .A2(_0388_),
    .B1(_0389_),
    .X(_0029_));
 sky130_fd_sc_hd__nor2_1 _0957_ (.A(\write_word[0] ),
    .B(net200),
    .Y(_0390_));
 sky130_fd_sc_hd__nand2_1 _0958_ (.A(\write_word[0] ),
    .B(net200),
    .Y(_0391_));
 sky130_fd_sc_hd__or3b_1 _0959_ (.A(_0304_),
    .B(_0390_),
    .C_N(_0391_),
    .X(_0392_));
 sky130_fd_sc_hd__nand2_1 _0960_ (.A(_0388_),
    .B(net200),
    .Y(_0393_));
 sky130_fd_sc_hd__o21ai_1 _0961_ (.A1(_0392_),
    .A2(_0388_),
    .B1(net201),
    .Y(_0030_));
 sky130_fd_sc_hd__xor2_1 _0962_ (.A(net205),
    .B(_0391_),
    .X(_0394_));
 sky130_fd_sc_hd__or2_1 _0963_ (.A(_0304_),
    .B(_0394_),
    .X(_0395_));
 sky130_fd_sc_hd__nand2_1 _0964_ (.A(_0388_),
    .B(net205),
    .Y(_0396_));
 sky130_fd_sc_hd__o21ai_1 _0965_ (.A1(_0395_),
    .A2(_0388_),
    .B1(net206),
    .Y(_0031_));
 sky130_fd_sc_hd__inv_2 _0966_ (.A(net319),
    .Y(_0397_));
 sky130_fd_sc_hd__nand2_1 _0967_ (.A(_0343_),
    .B(_0397_),
    .Y(_0398_));
 sky130_fd_sc_hd__nor2_1 _0968_ (.A(net203),
    .B(\state[2] ),
    .Y(_0399_));
 sky130_fd_sc_hd__a32o_1 _0969_ (.A1(_0398_),
    .A2(_0346_),
    .A3(\state[2] ),
    .B1(net319),
    .B2(_0399_),
    .X(_0032_));
 sky130_fd_sc_hd__inv_2 _0970_ (.A(net220),
    .Y(_0400_));
 sky130_fd_sc_hd__a21oi_1 _0971_ (.A1(_0400_),
    .A2(_0346_),
    .B1(_0349_),
    .Y(_0401_));
 sky130_fd_sc_hd__a21o_1 _0972_ (.A1(net220),
    .A2(_0399_),
    .B1(_0401_),
    .X(_0033_));
 sky130_fd_sc_hd__nand2_1 _0973_ (.A(_0284_),
    .B(\read_buf[0] ),
    .Y(_0402_));
 sky130_fd_sc_hd__a21oi_1 _0974_ (.A1(_0291_),
    .A2(_0402_),
    .B1(_0293_),
    .Y(_0034_));
 sky130_fd_sc_hd__nand2_1 _0975_ (.A(_0284_),
    .B(\read_buf[1] ),
    .Y(_0403_));
 sky130_fd_sc_hd__a21oi_1 _0976_ (.A1(_0289_),
    .A2(_0403_),
    .B1(_0293_),
    .Y(_0035_));
 sky130_fd_sc_hd__nand2_1 _0977_ (.A(_0284_),
    .B(\read_buf[2] ),
    .Y(_0404_));
 sky130_fd_sc_hd__a21oi_1 _0978_ (.A1(_0287_),
    .A2(_0404_),
    .B1(_0293_),
    .Y(_0036_));
 sky130_fd_sc_hd__nand2_1 _0979_ (.A(_0284_),
    .B(\read_buf[3] ),
    .Y(_0405_));
 sky130_fd_sc_hd__a21oi_1 _0980_ (.A1(_0285_),
    .A2(_0405_),
    .B1(_0293_),
    .Y(_0037_));
 sky130_fd_sc_hd__nand2_1 _0981_ (.A(_0274_),
    .B(\read_buf[8] ),
    .Y(_0406_));
 sky130_fd_sc_hd__a21oi_1 _0982_ (.A1(_0281_),
    .A2(_0406_),
    .B1(_0293_),
    .Y(_0038_));
 sky130_fd_sc_hd__nand2_1 _0983_ (.A(_0274_),
    .B(\read_buf[9] ),
    .Y(_0407_));
 sky130_fd_sc_hd__a21oi_1 _0984_ (.A1(_0279_),
    .A2(_0407_),
    .B1(_0293_),
    .Y(_0039_));
 sky130_fd_sc_hd__nand2_1 _0985_ (.A(_0274_),
    .B(\read_buf[10] ),
    .Y(_0408_));
 sky130_fd_sc_hd__a21oi_1 _0986_ (.A1(_0277_),
    .A2(_0408_),
    .B1(_0293_),
    .Y(_0040_));
 sky130_fd_sc_hd__nand2_1 _0987_ (.A(_0274_),
    .B(\read_buf[11] ),
    .Y(_0409_));
 sky130_fd_sc_hd__a21oi_1 _0988_ (.A1(_0275_),
    .A2(_0409_),
    .B1(_0293_),
    .Y(_0041_));
 sky130_fd_sc_hd__nand2_1 _0989_ (.A(_0264_),
    .B(\read_buf[16] ),
    .Y(_0410_));
 sky130_fd_sc_hd__a21oi_1 _0990_ (.A1(_0271_),
    .A2(_0410_),
    .B1(_0293_),
    .Y(_0042_));
 sky130_fd_sc_hd__nand2_1 _0991_ (.A(_0264_),
    .B(\read_buf[17] ),
    .Y(_0411_));
 sky130_fd_sc_hd__a21oi_1 _0992_ (.A1(_0269_),
    .A2(_0411_),
    .B1(_0293_),
    .Y(_0043_));
 sky130_fd_sc_hd__nand2_1 _0993_ (.A(_0264_),
    .B(\read_buf[18] ),
    .Y(_0412_));
 sky130_fd_sc_hd__a21oi_1 _0994_ (.A1(_0267_),
    .A2(_0412_),
    .B1(_0293_),
    .Y(_0044_));
 sky130_fd_sc_hd__nand2_1 _0995_ (.A(_0264_),
    .B(\read_buf[19] ),
    .Y(_0413_));
 sky130_fd_sc_hd__a21oi_1 _0996_ (.A1(_0265_),
    .A2(_0413_),
    .B1(_0293_),
    .Y(_0045_));
 sky130_fd_sc_hd__nand2_1 _0997_ (.A(_0246_),
    .B(\read_buf[24] ),
    .Y(_0414_));
 sky130_fd_sc_hd__a21oi_1 _0998_ (.A1(_0260_),
    .A2(_0414_),
    .B1(_0293_),
    .Y(_0046_));
 sky130_fd_sc_hd__nand2_1 _0999_ (.A(_0246_),
    .B(\read_buf[25] ),
    .Y(_0415_));
 sky130_fd_sc_hd__a21oi_1 _1000_ (.A1(_0257_),
    .A2(_0415_),
    .B1(_0293_),
    .Y(_0047_));
 sky130_fd_sc_hd__nand2_1 _1001_ (.A(_0246_),
    .B(\read_buf[26] ),
    .Y(_0416_));
 sky130_fd_sc_hd__a21oi_1 _1002_ (.A1(_0254_),
    .A2(_0416_),
    .B1(_0293_),
    .Y(_0048_));
 sky130_fd_sc_hd__nand2_1 _1003_ (.A(_0246_),
    .B(\read_buf[27] ),
    .Y(_0417_));
 sky130_fd_sc_hd__a21oi_1 _1004_ (.A1(_0417_),
    .A2(_0248_),
    .B1(_0249_),
    .Y(_0049_));
 sky130_fd_sc_hd__or3_1 _1005_ (.A(\read_byte[0] ),
    .B(_0249_),
    .C(_0245_),
    .X(_0418_));
 sky130_fd_sc_hd__inv_2 _1006_ (.A(_0418_),
    .Y(_0050_));
 sky130_fd_sc_hd__nand2_1 _1007_ (.A(_0251_),
    .B(_0252_),
    .Y(_0419_));
 sky130_fd_sc_hd__inv_2 _1008_ (.A(_0249_),
    .Y(_0420_));
 sky130_fd_sc_hd__and4_1 _1009_ (.A(_0246_),
    .B(_0244_),
    .C(_0419_),
    .D(_0420_),
    .X(_0421_));
 sky130_fd_sc_hd__clkbuf_1 _1010_ (.A(_0421_),
    .X(_0051_));
 sky130_fd_sc_hd__and3_1 _1011_ (.A(_0420_),
    .B(\read_byte[2] ),
    .C(_0244_),
    .X(_0422_));
 sky130_fd_sc_hd__clkbuf_1 _1012_ (.A(_0422_),
    .X(_0052_));
 sky130_fd_sc_hd__nor2_1 _1013_ (.A(_0250_),
    .B(_0246_),
    .Y(_0053_));
 sky130_fd_sc_hd__inv_2 _1014__1 (.A(clknet_3_1__leaf_clk_i),
    .Y(net109));
 sky130_fd_sc_hd__inv_2 _1015_ (.A(_0341_),
    .Y(_0014_));
 sky130_fd_sc_hd__inv_2 _1016_ (.A(_0341_),
    .Y(_0015_));
 sky130_fd_sc_hd__inv_2 _1017_ (.A(_0341_),
    .Y(_0016_));
 sky130_fd_sc_hd__inv_2 _1018_ (.A(_0341_),
    .Y(_0017_));
 sky130_fd_sc_hd__inv_2 _1019_ (.A(_0341_),
    .Y(_0018_));
 sky130_fd_sc_hd__inv_2 _1020_ (.A(_0341_),
    .Y(_0019_));
 sky130_fd_sc_hd__inv_2 _1021_ (.A(_0341_),
    .Y(_0020_));
 sky130_fd_sc_hd__inv_2 _1022_ (.A(_0341_),
    .Y(_0021_));
 sky130_fd_sc_hd__inv_2 _1023_ (.A(_0341_),
    .Y(_0022_));
 sky130_fd_sc_hd__inv_2 _1024_ (.A(_0341_),
    .Y(_0023_));
 sky130_fd_sc_hd__inv_2 _1025_ (.A(_0341_),
    .Y(_0024_));
 sky130_fd_sc_hd__inv_2 _1026_ (.A(_0341_),
    .Y(_0025_));
 sky130_fd_sc_hd__inv_2 _1027_ (.A(_0341_),
    .Y(_0026_));
 sky130_fd_sc_hd__inv_2 _1028_ (.A(_0341_),
    .Y(_0027_));
 sky130_fd_sc_hd__inv_2 _1029_ (.A(_0341_),
    .Y(_0028_));
 sky130_fd_sc_hd__or2_1 _1030_ (.A(\read_buf[0] ),
    .B(_0326_),
    .X(_0423_));
 sky130_fd_sc_hd__o21ai_1 _1031_ (.A1(\read_buf[24] ),
    .A2(_0364_),
    .B1(_0423_),
    .Y(_0424_));
 sky130_fd_sc_hd__nand2_4 _1032_ (.A(_0366_),
    .B(\state[11] ),
    .Y(_0425_));
 sky130_fd_sc_hd__buf_6 _1033_ (.A(_0425_),
    .X(_0426_));
 sky130_fd_sc_hd__buf_4 _1034_ (.A(_0425_),
    .X(_0427_));
 sky130_fd_sc_hd__nand2_1 _1035_ (.A(_0427_),
    .B(net313),
    .Y(_0428_));
 sky130_fd_sc_hd__o21ai_1 _1036_ (.A1(_0424_),
    .A2(_0426_),
    .B1(net314),
    .Y(_0070_));
 sky130_fd_sc_hd__or2_1 _1037_ (.A(\read_buf[1] ),
    .B(_0326_),
    .X(_0429_));
 sky130_fd_sc_hd__o21ai_1 _1038_ (.A1(\read_buf[25] ),
    .A2(_0364_),
    .B1(_0429_),
    .Y(_0430_));
 sky130_fd_sc_hd__nand2_1 _1039_ (.A(_0427_),
    .B(net271),
    .Y(_0431_));
 sky130_fd_sc_hd__o21ai_1 _1040_ (.A1(_0430_),
    .A2(_0426_),
    .B1(net272),
    .Y(_0071_));
 sky130_fd_sc_hd__or2_1 _1041_ (.A(\read_buf[2] ),
    .B(_0325_),
    .X(_0432_));
 sky130_fd_sc_hd__o21ai_1 _1042_ (.A1(\read_buf[26] ),
    .A2(_0364_),
    .B1(_0432_),
    .Y(_0433_));
 sky130_fd_sc_hd__nand2_1 _1043_ (.A(_0427_),
    .B(net295),
    .Y(_0434_));
 sky130_fd_sc_hd__o21ai_1 _1044_ (.A1(_0433_),
    .A2(_0426_),
    .B1(net296),
    .Y(_0072_));
 sky130_fd_sc_hd__or2_1 _1045_ (.A(\read_buf[3] ),
    .B(_0325_),
    .X(_0435_));
 sky130_fd_sc_hd__o21ai_1 _1046_ (.A1(\read_buf[27] ),
    .A2(_0364_),
    .B1(_0435_),
    .Y(_0436_));
 sky130_fd_sc_hd__nand2_1 _1047_ (.A(_0427_),
    .B(net310),
    .Y(_0437_));
 sky130_fd_sc_hd__o21ai_1 _1048_ (.A1(_0436_),
    .A2(_0426_),
    .B1(net311),
    .Y(_0073_));
 sky130_fd_sc_hd__or2_1 _1049_ (.A(\read_buf[4] ),
    .B(_0325_),
    .X(_0438_));
 sky130_fd_sc_hd__o21ai_1 _1050_ (.A1(\read_buf[28] ),
    .A2(_0364_),
    .B1(_0438_),
    .Y(_0439_));
 sky130_fd_sc_hd__nand2_1 _1051_ (.A(_0427_),
    .B(net280),
    .Y(_0440_));
 sky130_fd_sc_hd__o21ai_1 _1052_ (.A1(_0439_),
    .A2(_0426_),
    .B1(net281),
    .Y(_0074_));
 sky130_fd_sc_hd__or2_1 _1053_ (.A(\read_buf[5] ),
    .B(_0325_),
    .X(_0441_));
 sky130_fd_sc_hd__o21ai_1 _1054_ (.A1(\read_buf[29] ),
    .A2(_0364_),
    .B1(_0441_),
    .Y(_0442_));
 sky130_fd_sc_hd__nand2_1 _1055_ (.A(_0427_),
    .B(net304),
    .Y(_0443_));
 sky130_fd_sc_hd__o21ai_1 _1056_ (.A1(_0442_),
    .A2(_0426_),
    .B1(net305),
    .Y(_0075_));
 sky130_fd_sc_hd__or2_1 _1057_ (.A(\read_buf[6] ),
    .B(_0325_),
    .X(_0444_));
 sky130_fd_sc_hd__o21ai_1 _1058_ (.A1(\read_buf[30] ),
    .A2(_0364_),
    .B1(_0444_),
    .Y(_0445_));
 sky130_fd_sc_hd__nand2_1 _1059_ (.A(_0427_),
    .B(net211),
    .Y(_0446_));
 sky130_fd_sc_hd__o21ai_1 _1060_ (.A1(_0445_),
    .A2(_0426_),
    .B1(net212),
    .Y(_0076_));
 sky130_fd_sc_hd__or2_1 _1061_ (.A(\read_buf[7] ),
    .B(_0325_),
    .X(_0447_));
 sky130_fd_sc_hd__o21ai_1 _1062_ (.A1(\read_buf[31] ),
    .A2(_0364_),
    .B1(_0447_),
    .Y(_0448_));
 sky130_fd_sc_hd__nand2_1 _1063_ (.A(_0427_),
    .B(net262),
    .Y(_0449_));
 sky130_fd_sc_hd__o21ai_1 _1064_ (.A1(_0448_),
    .A2(_0426_),
    .B1(net263),
    .Y(_0077_));
 sky130_fd_sc_hd__buf_4 _1065_ (.A(_0326_),
    .X(_0450_));
 sky130_fd_sc_hd__nand2_1 _1066_ (.A(_0450_),
    .B(\read_buf[16] ),
    .Y(_0451_));
 sky130_fd_sc_hd__nand2_1 _1067_ (.A(_0427_),
    .B(net301),
    .Y(_0452_));
 sky130_fd_sc_hd__o21ai_1 _1068_ (.A1(_0451_),
    .A2(_0426_),
    .B1(net302),
    .Y(_0078_));
 sky130_fd_sc_hd__nand2_1 _1069_ (.A(_0450_),
    .B(\read_buf[17] ),
    .Y(_0453_));
 sky130_fd_sc_hd__nand2_1 _1070_ (.A(_0427_),
    .B(net217),
    .Y(_0454_));
 sky130_fd_sc_hd__o21ai_1 _1071_ (.A1(_0453_),
    .A2(_0426_),
    .B1(net218),
    .Y(_0079_));
 sky130_fd_sc_hd__nand2_1 _1072_ (.A(_0450_),
    .B(\read_buf[18] ),
    .Y(_0455_));
 sky130_fd_sc_hd__nand2_1 _1073_ (.A(_0427_),
    .B(net250),
    .Y(_0456_));
 sky130_fd_sc_hd__o21ai_1 _1074_ (.A1(_0455_),
    .A2(_0426_),
    .B1(net251),
    .Y(_0080_));
 sky130_fd_sc_hd__nand2_1 _1075_ (.A(_0450_),
    .B(\read_buf[19] ),
    .Y(_0457_));
 sky130_fd_sc_hd__nand2_1 _1076_ (.A(_0427_),
    .B(net225),
    .Y(_0458_));
 sky130_fd_sc_hd__o21ai_1 _1077_ (.A1(_0457_),
    .A2(_0426_),
    .B1(net226),
    .Y(_0081_));
 sky130_fd_sc_hd__nand2_1 _1078_ (.A(_0450_),
    .B(\read_buf[20] ),
    .Y(_0459_));
 sky130_fd_sc_hd__nand2_1 _1079_ (.A(_0427_),
    .B(net247),
    .Y(_0460_));
 sky130_fd_sc_hd__o21ai_1 _1080_ (.A1(_0459_),
    .A2(_0426_),
    .B1(net248),
    .Y(_0082_));
 sky130_fd_sc_hd__nand2_1 _1081_ (.A(_0450_),
    .B(\read_buf[21] ),
    .Y(_0461_));
 sky130_fd_sc_hd__nand2_1 _1082_ (.A(_0427_),
    .B(net222),
    .Y(_0462_));
 sky130_fd_sc_hd__o21ai_1 _1083_ (.A1(_0461_),
    .A2(_0426_),
    .B1(net223),
    .Y(_0083_));
 sky130_fd_sc_hd__nand2_1 _1084_ (.A(_0450_),
    .B(\read_buf[22] ),
    .Y(_0463_));
 sky130_fd_sc_hd__nand2_1 _1085_ (.A(_0427_),
    .B(net236),
    .Y(_0464_));
 sky130_fd_sc_hd__o21ai_1 _1086_ (.A1(_0463_),
    .A2(_0426_),
    .B1(net237),
    .Y(_0084_));
 sky130_fd_sc_hd__nand2_1 _1087_ (.A(_0450_),
    .B(\read_buf[23] ),
    .Y(_0465_));
 sky130_fd_sc_hd__nand2_1 _1088_ (.A(_0427_),
    .B(net253),
    .Y(_0466_));
 sky130_fd_sc_hd__o21ai_1 _1089_ (.A1(_0465_),
    .A2(_0426_),
    .B1(net254),
    .Y(_0085_));
 sky130_fd_sc_hd__nand2_1 _1090_ (.A(_0450_),
    .B(\read_buf[8] ),
    .Y(_0467_));
 sky130_fd_sc_hd__buf_6 _1091_ (.A(_0425_),
    .X(_0468_));
 sky130_fd_sc_hd__buf_4 _1092_ (.A(_0425_),
    .X(_0469_));
 sky130_fd_sc_hd__nand2_1 _1093_ (.A(_0469_),
    .B(net244),
    .Y(_0470_));
 sky130_fd_sc_hd__o21ai_1 _1094_ (.A1(_0467_),
    .A2(_0468_),
    .B1(net245),
    .Y(_0086_));
 sky130_fd_sc_hd__nand2_1 _1095_ (.A(_0450_),
    .B(\read_buf[9] ),
    .Y(_0471_));
 sky130_fd_sc_hd__nand2_1 _1096_ (.A(_0469_),
    .B(net233),
    .Y(_0472_));
 sky130_fd_sc_hd__o21ai_1 _1097_ (.A1(_0471_),
    .A2(_0468_),
    .B1(net234),
    .Y(_0087_));
 sky130_fd_sc_hd__nand2_1 _1098_ (.A(_0450_),
    .B(\read_buf[10] ),
    .Y(_0473_));
 sky130_fd_sc_hd__nand2_1 _1099_ (.A(_0469_),
    .B(net256),
    .Y(_0474_));
 sky130_fd_sc_hd__o21ai_1 _1100_ (.A1(_0473_),
    .A2(_0468_),
    .B1(net257),
    .Y(_0088_));
 sky130_fd_sc_hd__nand2_1 _1101_ (.A(_0450_),
    .B(\read_buf[11] ),
    .Y(_0475_));
 sky130_fd_sc_hd__nand2_1 _1102_ (.A(_0469_),
    .B(net230),
    .Y(_0476_));
 sky130_fd_sc_hd__o21ai_1 _1103_ (.A1(_0475_),
    .A2(_0468_),
    .B1(net231),
    .Y(_0089_));
 sky130_fd_sc_hd__nand2_1 _1104_ (.A(_0450_),
    .B(\read_buf[12] ),
    .Y(_0477_));
 sky130_fd_sc_hd__nand2_1 _1105_ (.A(_0469_),
    .B(net274),
    .Y(_0478_));
 sky130_fd_sc_hd__o21ai_1 _1106_ (.A1(_0477_),
    .A2(_0468_),
    .B1(net275),
    .Y(_0090_));
 sky130_fd_sc_hd__nand2_1 _1107_ (.A(_0450_),
    .B(\read_buf[13] ),
    .Y(_0479_));
 sky130_fd_sc_hd__nand2_1 _1108_ (.A(_0469_),
    .B(net259),
    .Y(_0480_));
 sky130_fd_sc_hd__o21ai_1 _1109_ (.A1(_0479_),
    .A2(_0468_),
    .B1(net260),
    .Y(_0091_));
 sky130_fd_sc_hd__nand2_1 _1110_ (.A(_0450_),
    .B(\read_buf[14] ),
    .Y(_0481_));
 sky130_fd_sc_hd__nand2_1 _1111_ (.A(_0469_),
    .B(net292),
    .Y(_0482_));
 sky130_fd_sc_hd__o21ai_1 _1112_ (.A1(_0481_),
    .A2(_0468_),
    .B1(net293),
    .Y(_0092_));
 sky130_fd_sc_hd__nand2_1 _1113_ (.A(_0450_),
    .B(\read_buf[15] ),
    .Y(_0483_));
 sky130_fd_sc_hd__nand2_1 _1114_ (.A(_0469_),
    .B(net277),
    .Y(_0484_));
 sky130_fd_sc_hd__o21ai_1 _1115_ (.A1(_0483_),
    .A2(_0468_),
    .B1(net278),
    .Y(_0093_));
 sky130_fd_sc_hd__nand2_1 _1116_ (.A(_0326_),
    .B(\read_buf[0] ),
    .Y(_0485_));
 sky130_fd_sc_hd__nand2_1 _1117_ (.A(_0469_),
    .B(net239),
    .Y(_0486_));
 sky130_fd_sc_hd__o21ai_1 _1118_ (.A1(_0485_),
    .A2(_0468_),
    .B1(net240),
    .Y(_0094_));
 sky130_fd_sc_hd__nand2_1 _1119_ (.A(_0326_),
    .B(\read_buf[1] ),
    .Y(_0487_));
 sky130_fd_sc_hd__nand2_1 _1120_ (.A(_0469_),
    .B(net316),
    .Y(_0488_));
 sky130_fd_sc_hd__o21ai_1 _1121_ (.A1(_0487_),
    .A2(_0468_),
    .B1(net317),
    .Y(_0095_));
 sky130_fd_sc_hd__nand2_1 _1122_ (.A(_0326_),
    .B(\read_buf[2] ),
    .Y(_0489_));
 sky130_fd_sc_hd__nand2_1 _1123_ (.A(_0469_),
    .B(net268),
    .Y(_0490_));
 sky130_fd_sc_hd__o21ai_1 _1124_ (.A1(_0489_),
    .A2(_0468_),
    .B1(net269),
    .Y(_0096_));
 sky130_fd_sc_hd__nand2_1 _1125_ (.A(_0326_),
    .B(\read_buf[3] ),
    .Y(_0491_));
 sky130_fd_sc_hd__nand2_1 _1126_ (.A(_0469_),
    .B(net289),
    .Y(_0492_));
 sky130_fd_sc_hd__o21ai_1 _1127_ (.A1(_0491_),
    .A2(_0468_),
    .B1(net290),
    .Y(_0097_));
 sky130_fd_sc_hd__nand2_1 _1128_ (.A(_0326_),
    .B(\read_buf[4] ),
    .Y(_0493_));
 sky130_fd_sc_hd__nand2_1 _1129_ (.A(_0469_),
    .B(net298),
    .Y(_0494_));
 sky130_fd_sc_hd__o21ai_1 _1130_ (.A1(_0493_),
    .A2(_0468_),
    .B1(net299),
    .Y(_0098_));
 sky130_fd_sc_hd__nand2_1 _1131_ (.A(_0326_),
    .B(\read_buf[5] ),
    .Y(_0495_));
 sky130_fd_sc_hd__nand2_1 _1132_ (.A(_0469_),
    .B(net283),
    .Y(_0496_));
 sky130_fd_sc_hd__o21ai_1 _1133_ (.A1(_0495_),
    .A2(_0468_),
    .B1(net284),
    .Y(_0099_));
 sky130_fd_sc_hd__nand2_1 _1134_ (.A(_0326_),
    .B(\read_buf[6] ),
    .Y(_0497_));
 sky130_fd_sc_hd__nand2_1 _1135_ (.A(_0469_),
    .B(net307),
    .Y(_0498_));
 sky130_fd_sc_hd__o21ai_1 _1136_ (.A1(_0497_),
    .A2(_0468_),
    .B1(net308),
    .Y(_0100_));
 sky130_fd_sc_hd__nand2_1 _1137_ (.A(_0326_),
    .B(\read_buf[7] ),
    .Y(_0499_));
 sky130_fd_sc_hd__nand2_1 _1138_ (.A(_0469_),
    .B(net324),
    .Y(_0500_));
 sky130_fd_sc_hd__o21ai_1 _1139_ (.A1(_0499_),
    .A2(_0468_),
    .B1(net325),
    .Y(_0101_));
 sky130_fd_sc_hd__inv_2 _1140_ (.A(net329),
    .Y(_0501_));
 sky130_fd_sc_hd__nor2_2 _1141_ (.A(net332),
    .B(_0501_),
    .Y(_0502_));
 sky130_fd_sc_hd__inv_2 _1142_ (.A(net214),
    .Y(_0503_));
 sky130_fd_sc_hd__nor2_1 _1143_ (.A(\state[9] ),
    .B(net339),
    .Y(_0504_));
 sky130_fd_sc_hd__a32o_1 _1144_ (.A1(_0502_),
    .A2(net339),
    .A3(_0503_),
    .B1(word_ready),
    .B2(_0504_),
    .X(_0505_));
 sky130_fd_sc_hd__o21ai_1 _1145_ (.A1(net337),
    .A2(_0504_),
    .B1(_0381_),
    .Y(_0506_));
 sky130_fd_sc_hd__nor2_1 _1146_ (.A(_0383_),
    .B(_0385_),
    .Y(_0507_));
 sky130_fd_sc_hd__nand3_1 _1147_ (.A(_0312_),
    .B(_0506_),
    .C(_0507_),
    .Y(_0508_));
 sky130_fd_sc_hd__mux2_1 _1148_ (.A0(_0505_),
    .A1(net343),
    .S(_0508_),
    .X(_0509_));
 sky130_fd_sc_hd__clkbuf_1 _1149_ (.A(net344),
    .X(_0102_));
 sky130_fd_sc_hd__buf_6 _1150_ (.A(_0307_),
    .X(_0510_));
 sky130_fd_sc_hd__inv_2 _1151_ (.A(net27),
    .Y(_0511_));
 sky130_fd_sc_hd__nand2_1 _1152_ (.A(_0510_),
    .B(_0511_),
    .Y(_0512_));
 sky130_fd_sc_hd__o21ai_1 _1153_ (.A1(net141),
    .A2(_0510_),
    .B1(_0512_),
    .Y(_0513_));
 sky130_fd_sc_hd__buf_4 _1154_ (.A(_0310_),
    .X(_0514_));
 sky130_fd_sc_hd__nand2_1 _1155_ (.A(_0513_),
    .B(_0514_),
    .Y(_0515_));
 sky130_fd_sc_hd__inv_2 _1156_ (.A(net23),
    .Y(_0516_));
 sky130_fd_sc_hd__nand2_1 _1157_ (.A(_0510_),
    .B(_0516_),
    .Y(_0517_));
 sky130_fd_sc_hd__o21ai_1 _1158_ (.A1(net129),
    .A2(_0510_),
    .B1(_0517_),
    .Y(_0518_));
 sky130_fd_sc_hd__nand2_1 _1159_ (.A(_0518_),
    .B(_0344_),
    .Y(_0519_));
 sky130_fd_sc_hd__nand2_1 _1160_ (.A(_0515_),
    .B(_0519_),
    .Y(_0520_));
 sky130_fd_sc_hd__nand2_1 _1161_ (.A(_0520_),
    .B(\write_byte[0] ),
    .Y(_0521_));
 sky130_fd_sc_hd__inv_2 _1162_ (.A(net19),
    .Y(_0522_));
 sky130_fd_sc_hd__nand2_1 _1163_ (.A(_0307_),
    .B(_0522_),
    .Y(_0523_));
 sky130_fd_sc_hd__o21ai_1 _1164_ (.A1(net131),
    .A2(_0510_),
    .B1(_0523_),
    .Y(_0524_));
 sky130_fd_sc_hd__nand2_1 _1165_ (.A(_0524_),
    .B(_0514_),
    .Y(_0525_));
 sky130_fd_sc_hd__inv_2 _1166_ (.A(net14),
    .Y(_0526_));
 sky130_fd_sc_hd__nand2_1 _1167_ (.A(_0307_),
    .B(_0526_),
    .Y(_0527_));
 sky130_fd_sc_hd__o21ai_1 _1168_ (.A1(net139),
    .A2(_0510_),
    .B1(_0527_),
    .Y(_0528_));
 sky130_fd_sc_hd__nand2_1 _1169_ (.A(_0528_),
    .B(_0343_),
    .Y(_0529_));
 sky130_fd_sc_hd__nand2_1 _1170_ (.A(_0525_),
    .B(_0529_),
    .Y(_0530_));
 sky130_fd_sc_hd__nand2_1 _1171_ (.A(_0530_),
    .B(_0501_),
    .Y(_0531_));
 sky130_fd_sc_hd__nand2_1 _1172_ (.A(_0521_),
    .B(_0531_),
    .Y(_0532_));
 sky130_fd_sc_hd__nand2_1 _1173_ (.A(_0532_),
    .B(\write_byte[1] ),
    .Y(_0533_));
 sky130_fd_sc_hd__nand2_1 _1174_ (.A(_0380_),
    .B(net159),
    .Y(_0534_));
 sky130_fd_sc_hd__nand2_1 _1175_ (.A(_0510_),
    .B(net61),
    .Y(_0535_));
 sky130_fd_sc_hd__nand3_1 _1176_ (.A(_0534_),
    .B(_0535_),
    .C(_0343_),
    .Y(_0536_));
 sky130_fd_sc_hd__nand2_1 _1177_ (.A(_0380_),
    .B(net147),
    .Y(_0537_));
 sky130_fd_sc_hd__nand2_1 _1178_ (.A(_0510_),
    .B(net10),
    .Y(_0538_));
 sky130_fd_sc_hd__nand3_1 _1179_ (.A(_0537_),
    .B(_0538_),
    .C(_0310_),
    .Y(_0539_));
 sky130_fd_sc_hd__nand2_1 _1180_ (.A(_0536_),
    .B(_0539_),
    .Y(_0540_));
 sky130_fd_sc_hd__nand2_1 _1181_ (.A(_0540_),
    .B(_0502_),
    .Y(_0541_));
 sky130_fd_sc_hd__nand2_1 _1182_ (.A(_0541_),
    .B(_0503_),
    .Y(_0542_));
 sky130_fd_sc_hd__buf_4 _1183_ (.A(_0307_),
    .X(_0543_));
 sky130_fd_sc_hd__inv_2 _1184_ (.A(net51),
    .Y(_0544_));
 sky130_fd_sc_hd__nand2_1 _1185_ (.A(_0543_),
    .B(_0544_),
    .Y(_0545_));
 sky130_fd_sc_hd__o21ai_1 _1186_ (.A1(net121),
    .A2(_0543_),
    .B1(_0545_),
    .Y(_0546_));
 sky130_fd_sc_hd__nand2_1 _1187_ (.A(_0546_),
    .B(_0514_),
    .Y(_0547_));
 sky130_fd_sc_hd__inv_2 _1188_ (.A(net7),
    .Y(_0548_));
 sky130_fd_sc_hd__nand2_1 _1189_ (.A(_0543_),
    .B(_0548_),
    .Y(_0549_));
 sky130_fd_sc_hd__o21ai_1 _1190_ (.A1(net123),
    .A2(_0543_),
    .B1(_0549_),
    .Y(_0550_));
 sky130_fd_sc_hd__nand2_1 _1191_ (.A(_0550_),
    .B(_0344_),
    .Y(_0551_));
 sky130_fd_sc_hd__nor2_1 _1192_ (.A(net332),
    .B(net329),
    .Y(_0552_));
 sky130_fd_sc_hd__inv_2 _1193_ (.A(_0552_),
    .Y(_0553_));
 sky130_fd_sc_hd__a21oi_1 _1194_ (.A1(_0547_),
    .A2(_0551_),
    .B1(_0553_),
    .Y(_0554_));
 sky130_fd_sc_hd__nor2_1 _1195_ (.A(_0542_),
    .B(_0554_),
    .Y(_0555_));
 sky130_fd_sc_hd__nand2_1 _1196_ (.A(_0533_),
    .B(_0555_),
    .Y(_0556_));
 sky130_fd_sc_hd__nand2_1 _1197_ (.A(_0556_),
    .B(_0326_),
    .Y(_0557_));
 sky130_fd_sc_hd__nand2_1 _1198_ (.A(_0344_),
    .B(net7),
    .Y(_0558_));
 sky130_fd_sc_hd__o211a_1 _1199_ (.A1(_0344_),
    .A2(_0544_),
    .B1(_0558_),
    .C1(_0364_),
    .X(_0559_));
 sky130_fd_sc_hd__nor2_1 _1200_ (.A(_0304_),
    .B(_0559_),
    .Y(_0560_));
 sky130_fd_sc_hd__nand2_1 _1201_ (.A(_0557_),
    .B(_0560_),
    .Y(_0561_));
 sky130_fd_sc_hd__nor2_1 _1202_ (.A(\current_nibble[1] ),
    .B(_0400_),
    .Y(_0562_));
 sky130_fd_sc_hd__mux2_1 _1203_ (.A0(net45),
    .A1(net49),
    .S(_0310_),
    .X(_0563_));
 sky130_fd_sc_hd__and3_1 _1204_ (.A(_0397_),
    .B(net33),
    .C(_0310_),
    .X(_0564_));
 sky130_fd_sc_hd__nand2_1 _1205_ (.A(_0343_),
    .B(net37),
    .Y(_0565_));
 sky130_fd_sc_hd__nand2_1 _1206_ (.A(net42),
    .B(_0310_),
    .Y(_0566_));
 sky130_fd_sc_hd__a21oi_1 _1207_ (.A1(_0565_),
    .A2(_0566_),
    .B1(_0397_),
    .Y(_0567_));
 sky130_fd_sc_hd__o21a_1 _1208_ (.A1(_0564_),
    .A2(_0567_),
    .B1(_0400_),
    .X(_0568_));
 sky130_fd_sc_hd__a21oi_1 _1209_ (.A1(_0562_),
    .A2(_0563_),
    .B1(_0568_),
    .Y(_0569_));
 sky130_fd_sc_hd__nor2_1 _1210_ (.A(\state[5] ),
    .B(\state[8] ),
    .Y(_0570_));
 sky130_fd_sc_hd__nand2_1 _1211_ (.A(_0570_),
    .B(_0350_),
    .Y(_0571_));
 sky130_fd_sc_hd__o211ai_4 _1212_ (.A1(net112),
    .A2(_0571_),
    .B1(net107),
    .C1(_0329_),
    .Y(_0572_));
 sky130_fd_sc_hd__inv_2 _1213_ (.A(_0572_),
    .Y(_0573_));
 sky130_fd_sc_hd__o21a_1 _1214_ (.A1(_0350_),
    .A2(_0569_),
    .B1(_0573_),
    .X(_0574_));
 sky130_fd_sc_hd__nor2_1 _1215_ (.A(net265),
    .B(_0573_),
    .Y(_0575_));
 sky130_fd_sc_hd__a21oi_1 _1216_ (.A1(_0561_),
    .A2(_0574_),
    .B1(net266),
    .Y(_0103_));
 sky130_fd_sc_hd__buf_4 _1217_ (.A(_0305_),
    .X(_0576_));
 sky130_fd_sc_hd__nand3b_1 _1218_ (.A_N(net125),
    .B(_0576_),
    .C(_0374_),
    .Y(_0577_));
 sky130_fd_sc_hd__inv_2 _1219_ (.A(net58),
    .Y(_0578_));
 sky130_fd_sc_hd__nand2_1 _1220_ (.A(_0543_),
    .B(_0578_),
    .Y(_0579_));
 sky130_fd_sc_hd__nand2_1 _1221_ (.A(_0577_),
    .B(_0579_),
    .Y(_0580_));
 sky130_fd_sc_hd__nand2_1 _1222_ (.A(_0580_),
    .B(_0514_),
    .Y(_0581_));
 sky130_fd_sc_hd__inv_2 _1223_ (.A(net18),
    .Y(_0582_));
 sky130_fd_sc_hd__nand2_1 _1224_ (.A(_0543_),
    .B(_0582_),
    .Y(_0583_));
 sky130_fd_sc_hd__inv_2 _1225_ (.A(net161),
    .Y(_0584_));
 sky130_fd_sc_hd__nand3_1 _1226_ (.A(_0576_),
    .B(_0584_),
    .C(_0374_),
    .Y(_0585_));
 sky130_fd_sc_hd__nand2_1 _1227_ (.A(_0583_),
    .B(_0585_),
    .Y(_0586_));
 sky130_fd_sc_hd__nand2_1 _1228_ (.A(_0586_),
    .B(_0344_),
    .Y(_0587_));
 sky130_fd_sc_hd__a21oi_1 _1229_ (.A1(_0581_),
    .A2(_0587_),
    .B1(_0553_),
    .Y(_0588_));
 sky130_fd_sc_hd__nand2_1 _1230_ (.A(_0543_),
    .B(net62),
    .Y(_0589_));
 sky130_fd_sc_hd__nand3_1 _1231_ (.A(_0576_),
    .B(_0374_),
    .C(net155),
    .Y(_0590_));
 sky130_fd_sc_hd__nand3_1 _1232_ (.A(_0589_),
    .B(_0343_),
    .C(_0590_),
    .Y(_0591_));
 sky130_fd_sc_hd__nand2_1 _1233_ (.A(_0543_),
    .B(net11),
    .Y(_0592_));
 sky130_fd_sc_hd__nand3_1 _1234_ (.A(_0576_),
    .B(_0374_),
    .C(net133),
    .Y(_0593_));
 sky130_fd_sc_hd__nand3_1 _1235_ (.A(_0592_),
    .B(_0514_),
    .C(_0593_),
    .Y(_0594_));
 sky130_fd_sc_hd__nand2_1 _1236_ (.A(_0591_),
    .B(_0594_),
    .Y(_0595_));
 sky130_fd_sc_hd__nand2_1 _1237_ (.A(_0595_),
    .B(_0502_),
    .Y(_0596_));
 sky130_fd_sc_hd__nand2_1 _1238_ (.A(_0596_),
    .B(_0503_),
    .Y(_0597_));
 sky130_fd_sc_hd__nor2_1 _1239_ (.A(_0588_),
    .B(_0597_),
    .Y(_0598_));
 sky130_fd_sc_hd__nand3b_1 _1240_ (.A_N(net115),
    .B(_0576_),
    .C(_0374_),
    .Y(_0599_));
 sky130_fd_sc_hd__inv_2 _1241_ (.A(net28),
    .Y(_0600_));
 sky130_fd_sc_hd__nand2_1 _1242_ (.A(_0307_),
    .B(_0600_),
    .Y(_0601_));
 sky130_fd_sc_hd__nand2_1 _1243_ (.A(_0599_),
    .B(_0601_),
    .Y(_0602_));
 sky130_fd_sc_hd__nand2_1 _1244_ (.A(_0602_),
    .B(_0514_),
    .Y(_0603_));
 sky130_fd_sc_hd__inv_2 _1245_ (.A(net24),
    .Y(_0604_));
 sky130_fd_sc_hd__nand2_1 _1246_ (.A(_0307_),
    .B(_0604_),
    .Y(_0605_));
 sky130_fd_sc_hd__inv_2 _1247_ (.A(net171),
    .Y(_0606_));
 sky130_fd_sc_hd__nand3_1 _1248_ (.A(_0576_),
    .B(_0606_),
    .C(_0374_),
    .Y(_0607_));
 sky130_fd_sc_hd__nand2_1 _1249_ (.A(_0605_),
    .B(_0607_),
    .Y(_0608_));
 sky130_fd_sc_hd__nand2_1 _1250_ (.A(_0608_),
    .B(_0343_),
    .Y(_0609_));
 sky130_fd_sc_hd__nand2_1 _1251_ (.A(_0603_),
    .B(_0609_),
    .Y(_0610_));
 sky130_fd_sc_hd__nand2_1 _1252_ (.A(_0610_),
    .B(\write_byte[0] ),
    .Y(_0611_));
 sky130_fd_sc_hd__inv_2 _1253_ (.A(net20),
    .Y(_0612_));
 sky130_fd_sc_hd__nand2_1 _1254_ (.A(_0307_),
    .B(_0612_),
    .Y(_0613_));
 sky130_fd_sc_hd__inv_2 _1255_ (.A(net169),
    .Y(_0614_));
 sky130_fd_sc_hd__nand3_1 _1256_ (.A(_0576_),
    .B(_0614_),
    .C(_0374_),
    .Y(_0615_));
 sky130_fd_sc_hd__nand2_1 _1257_ (.A(_0613_),
    .B(_0615_),
    .Y(_0616_));
 sky130_fd_sc_hd__nand2_1 _1258_ (.A(_0616_),
    .B(_0514_),
    .Y(_0617_));
 sky130_fd_sc_hd__inv_2 _1259_ (.A(net15),
    .Y(_0618_));
 sky130_fd_sc_hd__nand2_1 _1260_ (.A(_0307_),
    .B(_0618_),
    .Y(_0619_));
 sky130_fd_sc_hd__inv_2 _1261_ (.A(net165),
    .Y(_0620_));
 sky130_fd_sc_hd__nand3_1 _1262_ (.A(_0576_),
    .B(_0620_),
    .C(_0374_),
    .Y(_0621_));
 sky130_fd_sc_hd__nand2_1 _1263_ (.A(_0619_),
    .B(_0621_),
    .Y(_0622_));
 sky130_fd_sc_hd__nand2_1 _1264_ (.A(_0622_),
    .B(_0343_),
    .Y(_0623_));
 sky130_fd_sc_hd__nand2_1 _1265_ (.A(_0617_),
    .B(_0623_),
    .Y(_0624_));
 sky130_fd_sc_hd__nand2_1 _1266_ (.A(_0624_),
    .B(_0501_),
    .Y(_0625_));
 sky130_fd_sc_hd__nand2_1 _1267_ (.A(_0611_),
    .B(_0625_),
    .Y(_0626_));
 sky130_fd_sc_hd__nand2_1 _1268_ (.A(_0626_),
    .B(\write_byte[1] ),
    .Y(_0627_));
 sky130_fd_sc_hd__nand2_1 _1269_ (.A(_0598_),
    .B(_0627_),
    .Y(_0628_));
 sky130_fd_sc_hd__nand2_1 _1270_ (.A(_0628_),
    .B(_0326_),
    .Y(_0629_));
 sky130_fd_sc_hd__nand2_1 _1271_ (.A(_0344_),
    .B(net18),
    .Y(_0630_));
 sky130_fd_sc_hd__o211a_1 _1272_ (.A1(_0344_),
    .A2(_0578_),
    .B1(_0630_),
    .C1(_0364_),
    .X(_0631_));
 sky130_fd_sc_hd__nor2_1 _1273_ (.A(_0304_),
    .B(_0631_),
    .Y(_0632_));
 sky130_fd_sc_hd__nand2_1 _1274_ (.A(_0629_),
    .B(_0632_),
    .Y(_0633_));
 sky130_fd_sc_hd__mux2_1 _1275_ (.A0(net38),
    .A1(net43),
    .S(_0310_),
    .X(_0634_));
 sky130_fd_sc_hd__nand2_1 _1276_ (.A(_0634_),
    .B(\current_nibble[1] ),
    .Y(_0635_));
 sky130_fd_sc_hd__or3b_1 _1277_ (.A(_0343_),
    .B(\current_nibble[1] ),
    .C_N(net34),
    .X(_0636_));
 sky130_fd_sc_hd__nand2_1 _1278_ (.A(_0635_),
    .B(_0636_),
    .Y(_0637_));
 sky130_fd_sc_hd__nand2_1 _1279_ (.A(_0637_),
    .B(_0400_),
    .Y(_0638_));
 sky130_fd_sc_hd__mux2_1 _1280_ (.A0(net46),
    .A1(net50),
    .S(_0310_),
    .X(_0639_));
 sky130_fd_sc_hd__nand2_1 _1281_ (.A(_0639_),
    .B(_0562_),
    .Y(_0640_));
 sky130_fd_sc_hd__nand2_1 _1282_ (.A(_0638_),
    .B(_0640_),
    .Y(_0641_));
 sky130_fd_sc_hd__or2_1 _1283_ (.A(_0514_),
    .B(_0571_),
    .X(_0642_));
 sky130_fd_sc_hd__a21boi_1 _1284_ (.A1(_0641_),
    .A2(\state[2] ),
    .B1_N(_0642_),
    .Y(_0643_));
 sky130_fd_sc_hd__nand2_1 _1285_ (.A(_0633_),
    .B(_0643_),
    .Y(_0644_));
 sky130_fd_sc_hd__nand2_1 _1286_ (.A(_0644_),
    .B(_0573_),
    .Y(_0645_));
 sky130_fd_sc_hd__nand2_1 _1287_ (.A(_0572_),
    .B(net194),
    .Y(_0646_));
 sky130_fd_sc_hd__nand2_1 _1288_ (.A(_0645_),
    .B(net195),
    .Y(_0104_));
 sky130_fd_sc_hd__inv_2 _1289_ (.A(net30),
    .Y(_0647_));
 sky130_fd_sc_hd__nand2_1 _1290_ (.A(_0510_),
    .B(_0647_),
    .Y(_0648_));
 sky130_fd_sc_hd__o21ai_1 _1291_ (.A1(net143),
    .A2(_0510_),
    .B1(_0648_),
    .Y(_0649_));
 sky130_fd_sc_hd__nand2_1 _1292_ (.A(_0649_),
    .B(_0514_),
    .Y(_0650_));
 sky130_fd_sc_hd__inv_2 _1293_ (.A(net25),
    .Y(_0651_));
 sky130_fd_sc_hd__nand2_1 _1294_ (.A(_0307_),
    .B(_0651_),
    .Y(_0652_));
 sky130_fd_sc_hd__o21ai_1 _1295_ (.A1(net135),
    .A2(_0510_),
    .B1(_0652_),
    .Y(_0653_));
 sky130_fd_sc_hd__nand2_1 _1296_ (.A(_0653_),
    .B(_0343_),
    .Y(_0654_));
 sky130_fd_sc_hd__nand2_1 _1297_ (.A(_0650_),
    .B(_0654_),
    .Y(_0655_));
 sky130_fd_sc_hd__nand2_1 _1298_ (.A(_0655_),
    .B(\write_byte[0] ),
    .Y(_0656_));
 sky130_fd_sc_hd__inv_2 _1299_ (.A(net21),
    .Y(_0657_));
 sky130_fd_sc_hd__nand2_1 _1300_ (.A(_0307_),
    .B(_0657_),
    .Y(_0658_));
 sky130_fd_sc_hd__o21ai_1 _1301_ (.A1(net149),
    .A2(_0510_),
    .B1(_0658_),
    .Y(_0659_));
 sky130_fd_sc_hd__nand2_1 _1302_ (.A(_0659_),
    .B(_0514_),
    .Y(_0660_));
 sky130_fd_sc_hd__inv_2 _1303_ (.A(net16),
    .Y(_0661_));
 sky130_fd_sc_hd__nand2_1 _1304_ (.A(_0307_),
    .B(_0661_),
    .Y(_0662_));
 sky130_fd_sc_hd__o21ai_1 _1305_ (.A1(net137),
    .A2(_0510_),
    .B1(_0662_),
    .Y(_0663_));
 sky130_fd_sc_hd__nand2_1 _1306_ (.A(_0663_),
    .B(_0343_),
    .Y(_0664_));
 sky130_fd_sc_hd__nand2_1 _1307_ (.A(_0660_),
    .B(_0664_),
    .Y(_0665_));
 sky130_fd_sc_hd__nand2_1 _1308_ (.A(_0665_),
    .B(_0501_),
    .Y(_0666_));
 sky130_fd_sc_hd__nand2_1 _1309_ (.A(_0656_),
    .B(_0666_),
    .Y(_0667_));
 sky130_fd_sc_hd__nand2_1 _1310_ (.A(_0667_),
    .B(\write_byte[1] ),
    .Y(_0668_));
 sky130_fd_sc_hd__nand2_1 _1311_ (.A(_0380_),
    .B(net153),
    .Y(_0669_));
 sky130_fd_sc_hd__nand2_1 _1312_ (.A(_0510_),
    .B(net8),
    .Y(_0670_));
 sky130_fd_sc_hd__nand3_1 _1313_ (.A(_0669_),
    .B(_0670_),
    .C(_0343_),
    .Y(_0671_));
 sky130_fd_sc_hd__nand2_1 _1314_ (.A(_0380_),
    .B(net127),
    .Y(_0672_));
 sky130_fd_sc_hd__nand2_1 _1315_ (.A(_0510_),
    .B(net12),
    .Y(_0673_));
 sky130_fd_sc_hd__nand3_1 _1316_ (.A(_0672_),
    .B(_0673_),
    .C(_0310_),
    .Y(_0674_));
 sky130_fd_sc_hd__nand2_1 _1317_ (.A(_0671_),
    .B(_0674_),
    .Y(_0675_));
 sky130_fd_sc_hd__nand2_1 _1318_ (.A(_0675_),
    .B(_0502_),
    .Y(_0676_));
 sky130_fd_sc_hd__nand2_1 _1319_ (.A(_0676_),
    .B(_0503_),
    .Y(_0677_));
 sky130_fd_sc_hd__inv_2 _1320_ (.A(net59),
    .Y(_0678_));
 sky130_fd_sc_hd__nand2_1 _1321_ (.A(_0543_),
    .B(_0678_),
    .Y(_0679_));
 sky130_fd_sc_hd__o21ai_1 _1322_ (.A1(net117),
    .A2(_0543_),
    .B1(_0679_),
    .Y(_0680_));
 sky130_fd_sc_hd__nand2_1 _1323_ (.A(_0680_),
    .B(_0514_),
    .Y(_0681_));
 sky130_fd_sc_hd__inv_2 _1324_ (.A(net29),
    .Y(_0682_));
 sky130_fd_sc_hd__nand2_1 _1325_ (.A(_0543_),
    .B(_0682_),
    .Y(_0683_));
 sky130_fd_sc_hd__o21ai_1 _1326_ (.A1(net145),
    .A2(_0543_),
    .B1(_0683_),
    .Y(_0684_));
 sky130_fd_sc_hd__nand2_1 _1327_ (.A(_0684_),
    .B(_0344_),
    .Y(_0685_));
 sky130_fd_sc_hd__a21oi_1 _1328_ (.A1(_0681_),
    .A2(_0685_),
    .B1(_0553_),
    .Y(_0686_));
 sky130_fd_sc_hd__nor2_1 _1329_ (.A(_0677_),
    .B(_0686_),
    .Y(_0687_));
 sky130_fd_sc_hd__nand2_1 _1330_ (.A(_0668_),
    .B(_0687_),
    .Y(_0688_));
 sky130_fd_sc_hd__nand2_1 _1331_ (.A(_0688_),
    .B(_0326_),
    .Y(_0689_));
 sky130_fd_sc_hd__nand2_1 _1332_ (.A(_0344_),
    .B(net29),
    .Y(_0690_));
 sky130_fd_sc_hd__o211a_1 _1333_ (.A1(_0344_),
    .A2(_0678_),
    .B1(_0690_),
    .C1(_0364_),
    .X(_0691_));
 sky130_fd_sc_hd__nor2_1 _1334_ (.A(_0304_),
    .B(_0691_),
    .Y(_0692_));
 sky130_fd_sc_hd__nand2_1 _1335_ (.A(_0689_),
    .B(_0692_),
    .Y(_0693_));
 sky130_fd_sc_hd__mux2_1 _1336_ (.A0(net47),
    .A1(net52),
    .S(_0310_),
    .X(_0694_));
 sky130_fd_sc_hd__a21oi_1 _1337_ (.A1(_0694_),
    .A2(_0397_),
    .B1(_0400_),
    .Y(_0695_));
 sky130_fd_sc_hd__a22o_1 _1338_ (.A1(_0343_),
    .A2(net39),
    .B1(net35),
    .B2(_0397_),
    .X(_0696_));
 sky130_fd_sc_hd__a21o_1 _1339_ (.A1(_0696_),
    .A2(_0398_),
    .B1(net220),
    .X(_0697_));
 sky130_fd_sc_hd__nand2_1 _1340_ (.A(_0697_),
    .B(\state[2] ),
    .Y(_0698_));
 sky130_fd_sc_hd__o21ai_1 _1341_ (.A1(_0695_),
    .A2(_0698_),
    .B1(_0573_),
    .Y(_0699_));
 sky130_fd_sc_hd__inv_2 _1342_ (.A(_0699_),
    .Y(_0700_));
 sky130_fd_sc_hd__nor2_1 _1343_ (.A(net321),
    .B(_0573_),
    .Y(_0701_));
 sky130_fd_sc_hd__a21oi_1 _1344_ (.A1(_0693_),
    .A2(_0700_),
    .B1(net322),
    .Y(_0105_));
 sky130_fd_sc_hd__nand3b_1 _1345_ (.A_N(net113),
    .B(_0576_),
    .C(_0374_),
    .Y(_0702_));
 sky130_fd_sc_hd__inv_2 _1346_ (.A(net60),
    .Y(_0703_));
 sky130_fd_sc_hd__nand2_1 _1347_ (.A(_0543_),
    .B(_0703_),
    .Y(_0704_));
 sky130_fd_sc_hd__nand2_1 _1348_ (.A(_0702_),
    .B(_0704_),
    .Y(_0705_));
 sky130_fd_sc_hd__nand2_1 _1349_ (.A(_0705_),
    .B(_0514_),
    .Y(_0706_));
 sky130_fd_sc_hd__inv_2 _1350_ (.A(net40),
    .Y(_0707_));
 sky130_fd_sc_hd__nand2_1 _1351_ (.A(_0543_),
    .B(_0707_),
    .Y(_0708_));
 sky130_fd_sc_hd__inv_2 _1352_ (.A(net175),
    .Y(_0709_));
 sky130_fd_sc_hd__nand3_1 _1353_ (.A(_0576_),
    .B(_0709_),
    .C(_0374_),
    .Y(_0710_));
 sky130_fd_sc_hd__nand2_1 _1354_ (.A(_0708_),
    .B(_0710_),
    .Y(_0711_));
 sky130_fd_sc_hd__nand2_1 _1355_ (.A(_0711_),
    .B(_0344_),
    .Y(_0712_));
 sky130_fd_sc_hd__a21oi_1 _1356_ (.A1(_0706_),
    .A2(_0712_),
    .B1(_0553_),
    .Y(_0713_));
 sky130_fd_sc_hd__nand2_1 _1357_ (.A(_0543_),
    .B(net9),
    .Y(_0714_));
 sky130_fd_sc_hd__nand3_1 _1358_ (.A(_0576_),
    .B(_0374_),
    .C(net151),
    .Y(_0715_));
 sky130_fd_sc_hd__nand3_1 _1359_ (.A(_0714_),
    .B(_0343_),
    .C(_0715_),
    .Y(_0716_));
 sky130_fd_sc_hd__nand2_1 _1360_ (.A(_0510_),
    .B(net13),
    .Y(_0717_));
 sky130_fd_sc_hd__nand3_1 _1361_ (.A(_0576_),
    .B(_0374_),
    .C(net157),
    .Y(_0718_));
 sky130_fd_sc_hd__nand3_1 _1362_ (.A(_0717_),
    .B(_0310_),
    .C(_0718_),
    .Y(_0719_));
 sky130_fd_sc_hd__nand2_1 _1363_ (.A(_0716_),
    .B(_0719_),
    .Y(_0720_));
 sky130_fd_sc_hd__nand2_1 _1364_ (.A(_0720_),
    .B(_0502_),
    .Y(_0721_));
 sky130_fd_sc_hd__nand2_1 _1365_ (.A(_0721_),
    .B(_0503_),
    .Y(_0722_));
 sky130_fd_sc_hd__nor2_1 _1366_ (.A(_0713_),
    .B(_0722_),
    .Y(_0723_));
 sky130_fd_sc_hd__nand3b_1 _1367_ (.A_N(net119),
    .B(_0576_),
    .C(_0374_),
    .Y(_0724_));
 sky130_fd_sc_hd__inv_2 _1368_ (.A(net31),
    .Y(_0725_));
 sky130_fd_sc_hd__nand2_1 _1369_ (.A(_0307_),
    .B(_0725_),
    .Y(_0726_));
 sky130_fd_sc_hd__nand2_1 _1370_ (.A(_0724_),
    .B(_0726_),
    .Y(_0727_));
 sky130_fd_sc_hd__nand2_1 _1371_ (.A(_0727_),
    .B(_0514_),
    .Y(_0728_));
 sky130_fd_sc_hd__inv_2 _1372_ (.A(net26),
    .Y(_0729_));
 sky130_fd_sc_hd__nand2_1 _1373_ (.A(_0307_),
    .B(_0729_),
    .Y(_0730_));
 sky130_fd_sc_hd__inv_2 _1374_ (.A(net163),
    .Y(_0731_));
 sky130_fd_sc_hd__nand3_1 _1375_ (.A(_0576_),
    .B(_0731_),
    .C(_0374_),
    .Y(_0732_));
 sky130_fd_sc_hd__nand2_1 _1376_ (.A(_0730_),
    .B(_0732_),
    .Y(_0733_));
 sky130_fd_sc_hd__nand2_1 _1377_ (.A(_0733_),
    .B(_0343_),
    .Y(_0734_));
 sky130_fd_sc_hd__nand2_1 _1378_ (.A(_0728_),
    .B(_0734_),
    .Y(_0735_));
 sky130_fd_sc_hd__nand2_1 _1379_ (.A(_0735_),
    .B(\write_byte[0] ),
    .Y(_0736_));
 sky130_fd_sc_hd__inv_2 _1380_ (.A(net22),
    .Y(_0737_));
 sky130_fd_sc_hd__nand2_1 _1381_ (.A(_0307_),
    .B(_0737_),
    .Y(_0738_));
 sky130_fd_sc_hd__inv_2 _1382_ (.A(net173),
    .Y(_0739_));
 sky130_fd_sc_hd__nand3_1 _1383_ (.A(_0576_),
    .B(_0739_),
    .C(_0374_),
    .Y(_0740_));
 sky130_fd_sc_hd__nand2_1 _1384_ (.A(_0738_),
    .B(_0740_),
    .Y(_0741_));
 sky130_fd_sc_hd__nand2_1 _1385_ (.A(_0741_),
    .B(_0514_),
    .Y(_0742_));
 sky130_fd_sc_hd__inv_2 _1386_ (.A(net17),
    .Y(_0743_));
 sky130_fd_sc_hd__nand2_1 _1387_ (.A(_0307_),
    .B(_0743_),
    .Y(_0744_));
 sky130_fd_sc_hd__inv_2 _1388_ (.A(net167),
    .Y(_0745_));
 sky130_fd_sc_hd__nand3_1 _1389_ (.A(_0576_),
    .B(_0745_),
    .C(net56),
    .Y(_0746_));
 sky130_fd_sc_hd__nand2_1 _1390_ (.A(_0744_),
    .B(_0746_),
    .Y(_0747_));
 sky130_fd_sc_hd__nand2_1 _1391_ (.A(_0747_),
    .B(_0343_),
    .Y(_0748_));
 sky130_fd_sc_hd__nand2_1 _1392_ (.A(_0742_),
    .B(_0748_),
    .Y(_0749_));
 sky130_fd_sc_hd__nand2_1 _1393_ (.A(_0749_),
    .B(_0501_),
    .Y(_0750_));
 sky130_fd_sc_hd__nand2_1 _1394_ (.A(_0736_),
    .B(_0750_),
    .Y(_0751_));
 sky130_fd_sc_hd__nand2_1 _1395_ (.A(_0751_),
    .B(\write_byte[1] ),
    .Y(_0752_));
 sky130_fd_sc_hd__nand2_1 _1396_ (.A(_0723_),
    .B(_0752_),
    .Y(_0753_));
 sky130_fd_sc_hd__nand2_1 _1397_ (.A(_0753_),
    .B(_0326_),
    .Y(_0754_));
 sky130_fd_sc_hd__nand2_1 _1398_ (.A(_0344_),
    .B(net40),
    .Y(_0755_));
 sky130_fd_sc_hd__o211a_1 _1399_ (.A1(_0344_),
    .A2(_0703_),
    .B1(_0755_),
    .C1(_0364_),
    .X(_0756_));
 sky130_fd_sc_hd__nor2_1 _1400_ (.A(_0304_),
    .B(_0756_),
    .Y(_0757_));
 sky130_fd_sc_hd__nand2_1 _1401_ (.A(_0754_),
    .B(_0757_),
    .Y(_0758_));
 sky130_fd_sc_hd__mux2_1 _1402_ (.A0(net41),
    .A1(net44),
    .S(_0310_),
    .X(_0759_));
 sky130_fd_sc_hd__nand2_1 _1403_ (.A(_0759_),
    .B(\current_nibble[1] ),
    .Y(_0760_));
 sky130_fd_sc_hd__mux2_1 _1404_ (.A0(net32),
    .A1(net36),
    .S(_0310_),
    .X(_0761_));
 sky130_fd_sc_hd__nand2_1 _1405_ (.A(_0761_),
    .B(_0397_),
    .Y(_0762_));
 sky130_fd_sc_hd__nand2_1 _1406_ (.A(_0760_),
    .B(_0762_),
    .Y(_0763_));
 sky130_fd_sc_hd__nand2_1 _1407_ (.A(_0763_),
    .B(_0400_),
    .Y(_0764_));
 sky130_fd_sc_hd__mux2_1 _1408_ (.A0(net48),
    .A1(net53),
    .S(_0310_),
    .X(_0765_));
 sky130_fd_sc_hd__nand2_1 _1409_ (.A(_0765_),
    .B(_0562_),
    .Y(_0766_));
 sky130_fd_sc_hd__nand2_1 _1410_ (.A(_0764_),
    .B(_0766_),
    .Y(_0767_));
 sky130_fd_sc_hd__nor2_1 _1411_ (.A(net57),
    .B(_0642_),
    .Y(_0768_));
 sky130_fd_sc_hd__a21oi_1 _1412_ (.A1(_0767_),
    .A2(\state[2] ),
    .B1(_0768_),
    .Y(_0769_));
 sky130_fd_sc_hd__nand2_1 _1413_ (.A(_0758_),
    .B(_0769_),
    .Y(_0770_));
 sky130_fd_sc_hd__nand2_1 _1414_ (.A(_0770_),
    .B(_0573_),
    .Y(_0771_));
 sky130_fd_sc_hd__nand2_1 _1415_ (.A(_0572_),
    .B(net197),
    .Y(_0772_));
 sky130_fd_sc_hd__nand2_1 _1416_ (.A(_0771_),
    .B(net198),
    .Y(_0106_));
 sky130_fd_sc_hd__and4b_1 _1417_ (.A_N(_0570_),
    .B(_0507_),
    .C(net107),
    .D(_0360_),
    .X(_0773_));
 sky130_fd_sc_hd__nor2_1 _1418_ (.A(_0386_),
    .B(_0340_),
    .Y(_0774_));
 sky130_fd_sc_hd__nand3_2 _1419_ (.A(_0773_),
    .B(_0774_),
    .C(_0355_),
    .Y(_0775_));
 sky130_fd_sc_hd__buf_4 _1420_ (.A(_0775_),
    .X(_0776_));
 sky130_fd_sc_hd__buf_4 _1421_ (.A(_0775_),
    .X(_0777_));
 sky130_fd_sc_hd__nand2_1 _1422_ (.A(_0777_),
    .B(net123),
    .Y(_0778_));
 sky130_fd_sc_hd__o21ai_1 _1423_ (.A1(_0548_),
    .A2(_0776_),
    .B1(net124),
    .Y(_0107_));
 sky130_fd_sc_hd__nand2_1 _1424_ (.A(_0777_),
    .B(net161),
    .Y(_0153_));
 sky130_fd_sc_hd__o21ai_1 _1425_ (.A1(_0582_),
    .A2(_0776_),
    .B1(net162),
    .Y(_0108_));
 sky130_fd_sc_hd__nand2_1 _1426_ (.A(_0777_),
    .B(net145),
    .Y(_0154_));
 sky130_fd_sc_hd__o21ai_1 _1427_ (.A1(_0682_),
    .A2(_0776_),
    .B1(net146),
    .Y(_0109_));
 sky130_fd_sc_hd__nand2_1 _1428_ (.A(_0777_),
    .B(net175),
    .Y(_0155_));
 sky130_fd_sc_hd__o21ai_1 _1429_ (.A1(_0707_),
    .A2(_0776_),
    .B1(net176),
    .Y(_0110_));
 sky130_fd_sc_hd__nand2_1 _1430_ (.A(_0777_),
    .B(net121),
    .Y(_0156_));
 sky130_fd_sc_hd__o21ai_1 _1431_ (.A1(_0544_),
    .A2(_0776_),
    .B1(net122),
    .Y(_0111_));
 sky130_fd_sc_hd__nand2_1 _1432_ (.A(_0777_),
    .B(net125),
    .Y(_0157_));
 sky130_fd_sc_hd__o21ai_1 _1433_ (.A1(_0578_),
    .A2(_0776_),
    .B1(net126),
    .Y(_0112_));
 sky130_fd_sc_hd__nand2_1 _1434_ (.A(_0777_),
    .B(net117),
    .Y(_0158_));
 sky130_fd_sc_hd__o21ai_1 _1435_ (.A1(_0678_),
    .A2(_0776_),
    .B1(net118),
    .Y(_0113_));
 sky130_fd_sc_hd__nand2_1 _1436_ (.A(_0777_),
    .B(net113),
    .Y(_0159_));
 sky130_fd_sc_hd__o21ai_1 _1437_ (.A1(_0703_),
    .A2(_0776_),
    .B1(net114),
    .Y(_0114_));
 sky130_fd_sc_hd__inv_2 _1438_ (.A(net61),
    .Y(_0160_));
 sky130_fd_sc_hd__nand2_1 _1439_ (.A(_0777_),
    .B(net159),
    .Y(_0161_));
 sky130_fd_sc_hd__o21ai_1 _1440_ (.A1(_0160_),
    .A2(_0776_),
    .B1(net160),
    .Y(_0115_));
 sky130_fd_sc_hd__inv_2 _1441_ (.A(net62),
    .Y(_0162_));
 sky130_fd_sc_hd__nand2_1 _1442_ (.A(_0777_),
    .B(net155),
    .Y(_0163_));
 sky130_fd_sc_hd__o21ai_1 _1443_ (.A1(_0162_),
    .A2(_0776_),
    .B1(net156),
    .Y(_0116_));
 sky130_fd_sc_hd__inv_2 _1444_ (.A(net8),
    .Y(_0164_));
 sky130_fd_sc_hd__nand2_1 _1445_ (.A(_0777_),
    .B(net153),
    .Y(_0165_));
 sky130_fd_sc_hd__o21ai_1 _1446_ (.A1(_0164_),
    .A2(_0776_),
    .B1(net154),
    .Y(_0117_));
 sky130_fd_sc_hd__inv_2 _1447_ (.A(net9),
    .Y(_0166_));
 sky130_fd_sc_hd__nand2_1 _1448_ (.A(_0777_),
    .B(net151),
    .Y(_0167_));
 sky130_fd_sc_hd__o21ai_1 _1449_ (.A1(_0166_),
    .A2(_0776_),
    .B1(net152),
    .Y(_0118_));
 sky130_fd_sc_hd__inv_2 _1450_ (.A(net10),
    .Y(_0168_));
 sky130_fd_sc_hd__nand2_1 _1451_ (.A(_0777_),
    .B(net147),
    .Y(_0169_));
 sky130_fd_sc_hd__o21ai_1 _1452_ (.A1(_0168_),
    .A2(_0776_),
    .B1(net148),
    .Y(_0119_));
 sky130_fd_sc_hd__inv_2 _1453_ (.A(net11),
    .Y(_0170_));
 sky130_fd_sc_hd__nand2_1 _1454_ (.A(_0777_),
    .B(net133),
    .Y(_0171_));
 sky130_fd_sc_hd__o21ai_1 _1455_ (.A1(_0170_),
    .A2(_0776_),
    .B1(net134),
    .Y(_0120_));
 sky130_fd_sc_hd__inv_2 _1456_ (.A(net12),
    .Y(_0172_));
 sky130_fd_sc_hd__nand2_1 _1457_ (.A(_0777_),
    .B(net127),
    .Y(_0173_));
 sky130_fd_sc_hd__o21ai_1 _1458_ (.A1(_0172_),
    .A2(_0776_),
    .B1(net128),
    .Y(_0121_));
 sky130_fd_sc_hd__inv_2 _1459_ (.A(net13),
    .Y(_0174_));
 sky130_fd_sc_hd__nand2_1 _1460_ (.A(_0777_),
    .B(net157),
    .Y(_0175_));
 sky130_fd_sc_hd__o21ai_1 _1461_ (.A1(_0174_),
    .A2(_0776_),
    .B1(net158),
    .Y(_0122_));
 sky130_fd_sc_hd__buf_4 _1462_ (.A(_0775_),
    .X(_0176_));
 sky130_fd_sc_hd__buf_4 _1463_ (.A(_0775_),
    .X(_0177_));
 sky130_fd_sc_hd__nand2_1 _1464_ (.A(_0177_),
    .B(net139),
    .Y(_0178_));
 sky130_fd_sc_hd__o21ai_1 _1465_ (.A1(_0526_),
    .A2(_0176_),
    .B1(net140),
    .Y(_0123_));
 sky130_fd_sc_hd__nand2_1 _1466_ (.A(_0177_),
    .B(net165),
    .Y(_0179_));
 sky130_fd_sc_hd__o21ai_1 _1467_ (.A1(_0618_),
    .A2(_0176_),
    .B1(net166),
    .Y(_0124_));
 sky130_fd_sc_hd__nand2_1 _1468_ (.A(_0177_),
    .B(net137),
    .Y(_0180_));
 sky130_fd_sc_hd__o21ai_1 _1469_ (.A1(_0661_),
    .A2(_0176_),
    .B1(net138),
    .Y(_0125_));
 sky130_fd_sc_hd__nand2_1 _1470_ (.A(_0177_),
    .B(net167),
    .Y(_0181_));
 sky130_fd_sc_hd__o21ai_1 _1471_ (.A1(_0743_),
    .A2(_0176_),
    .B1(net168),
    .Y(_0126_));
 sky130_fd_sc_hd__nand2_1 _1472_ (.A(_0177_),
    .B(net131),
    .Y(_0182_));
 sky130_fd_sc_hd__o21ai_1 _1473_ (.A1(_0522_),
    .A2(_0176_),
    .B1(net132),
    .Y(_0127_));
 sky130_fd_sc_hd__nand2_1 _1474_ (.A(_0177_),
    .B(net169),
    .Y(_0183_));
 sky130_fd_sc_hd__o21ai_1 _1475_ (.A1(_0612_),
    .A2(_0176_),
    .B1(net170),
    .Y(_0128_));
 sky130_fd_sc_hd__nand2_1 _1476_ (.A(_0177_),
    .B(net149),
    .Y(_0184_));
 sky130_fd_sc_hd__o21ai_1 _1477_ (.A1(_0657_),
    .A2(_0176_),
    .B1(net150),
    .Y(_0129_));
 sky130_fd_sc_hd__nand2_1 _1478_ (.A(_0177_),
    .B(net173),
    .Y(_0185_));
 sky130_fd_sc_hd__o21ai_1 _1479_ (.A1(_0737_),
    .A2(_0176_),
    .B1(net174),
    .Y(_0130_));
 sky130_fd_sc_hd__nand2_1 _1480_ (.A(_0177_),
    .B(net129),
    .Y(_0186_));
 sky130_fd_sc_hd__o21ai_1 _1481_ (.A1(_0516_),
    .A2(_0176_),
    .B1(net130),
    .Y(_0131_));
 sky130_fd_sc_hd__nand2_1 _1482_ (.A(_0177_),
    .B(net171),
    .Y(_0187_));
 sky130_fd_sc_hd__o21ai_1 _1483_ (.A1(_0604_),
    .A2(_0176_),
    .B1(net172),
    .Y(_0132_));
 sky130_fd_sc_hd__nand2_1 _1484_ (.A(_0177_),
    .B(net135),
    .Y(_0188_));
 sky130_fd_sc_hd__o21ai_1 _1485_ (.A1(_0651_),
    .A2(_0176_),
    .B1(net136),
    .Y(_0133_));
 sky130_fd_sc_hd__nand2_1 _1486_ (.A(_0177_),
    .B(net163),
    .Y(_0189_));
 sky130_fd_sc_hd__o21ai_1 _1487_ (.A1(_0729_),
    .A2(_0176_),
    .B1(net164),
    .Y(_0134_));
 sky130_fd_sc_hd__nand2_1 _1488_ (.A(_0177_),
    .B(net141),
    .Y(_0190_));
 sky130_fd_sc_hd__o21ai_1 _1489_ (.A1(_0511_),
    .A2(_0176_),
    .B1(net142),
    .Y(_0135_));
 sky130_fd_sc_hd__nand2_1 _1490_ (.A(_0177_),
    .B(net115),
    .Y(_0191_));
 sky130_fd_sc_hd__o21ai_1 _1491_ (.A1(_0600_),
    .A2(_0176_),
    .B1(net116),
    .Y(_0136_));
 sky130_fd_sc_hd__nand2_1 _1492_ (.A(_0177_),
    .B(net143),
    .Y(_0192_));
 sky130_fd_sc_hd__o21ai_1 _1493_ (.A1(_0647_),
    .A2(_0176_),
    .B1(net144),
    .Y(_0137_));
 sky130_fd_sc_hd__nand2_1 _1494_ (.A(_0177_),
    .B(net119),
    .Y(_0193_));
 sky130_fd_sc_hd__o21ai_1 _1495_ (.A1(_0725_),
    .A2(_0176_),
    .B1(net120),
    .Y(_0138_));
 sky130_fd_sc_hd__nor2_1 _1496_ (.A(net180),
    .B(net64),
    .Y(_0194_));
 sky130_fd_sc_hd__o21a_1 _1497_ (.A1(net112),
    .A2(net352),
    .B1(net181),
    .X(_0139_));
 sky130_fd_sc_hd__and3_1 _1498_ (.A(_0304_),
    .B(_0350_),
    .C(_0345_),
    .X(_0195_));
 sky130_fd_sc_hd__a21o_1 _1499_ (.A1(_0195_),
    .A2(_0379_),
    .B1(_0328_),
    .X(_0196_));
 sky130_fd_sc_hd__nand2_1 _1500_ (.A(_0385_),
    .B(_0324_),
    .Y(_0197_));
 sky130_fd_sc_hd__a211oi_1 _1501_ (.A1(_0514_),
    .A2(_0197_),
    .B1(_0195_),
    .C1(_0196_),
    .Y(_0198_));
 sky130_fd_sc_hd__a21o_1 _1502_ (.A1(_0514_),
    .A2(_0196_),
    .B1(_0198_),
    .X(_0140_));
 sky130_fd_sc_hd__nand2_1 _1503_ (.A(_0337_),
    .B(net286),
    .Y(_0199_));
 sky130_fd_sc_hd__o21ai_1 _1504_ (.A1(net203),
    .A2(net286),
    .B1(_0199_),
    .Y(_0200_));
 sky130_fd_sc_hd__or2_1 _1505_ (.A(_0333_),
    .B(_0200_),
    .X(_0201_));
 sky130_fd_sc_hd__inv_2 _1506_ (.A(_0201_),
    .Y(_0202_));
 sky130_fd_sc_hd__mux2_1 _1507_ (.A0(_0202_),
    .A1(_0200_),
    .S(net327),
    .X(_0203_));
 sky130_fd_sc_hd__clkbuf_1 _1508_ (.A(_0203_),
    .X(_0141_));
 sky130_fd_sc_hd__or2_1 _1509_ (.A(net192),
    .B(_0334_),
    .X(_0204_));
 sky130_fd_sc_hd__nand2_1 _1510_ (.A(_0204_),
    .B(_0335_),
    .Y(_0205_));
 sky130_fd_sc_hd__a22o_1 _1511_ (.A1(net192),
    .A2(_0200_),
    .B1(_0202_),
    .B2(_0205_),
    .X(_0142_));
 sky130_fd_sc_hd__nor2_1 _1512_ (.A(_0359_),
    .B(_0320_),
    .Y(_0206_));
 sky130_fd_sc_hd__o2111ai_1 _1513_ (.A1(\state[6] ),
    .A2(\state[8] ),
    .B1(_0199_),
    .C1(_0206_),
    .D1(_0357_),
    .Y(_0207_));
 sky130_fd_sc_hd__and2_1 _1514_ (.A(_0013_),
    .B(net177),
    .X(_0208_));
 sky130_fd_sc_hd__o22a_1 _1515_ (.A1(\state[6] ),
    .A2(\state[8] ),
    .B1(_0208_),
    .B2(_0199_),
    .X(_0209_));
 sky130_fd_sc_hd__nand2_1 _1516_ (.A(_0206_),
    .B(_0209_),
    .Y(_0210_));
 sky130_fd_sc_hd__a21o_1 _1517_ (.A1(_0340_),
    .A2(_0013_),
    .B1(_0356_),
    .X(_0211_));
 sky130_fd_sc_hd__o21ai_1 _1518_ (.A1(_0210_),
    .A2(_0211_),
    .B1(net177),
    .Y(_0212_));
 sky130_fd_sc_hd__nand2_1 _1519_ (.A(_0207_),
    .B(net178),
    .Y(_0143_));
 sky130_fd_sc_hd__nor2_1 _1520_ (.A(\state[8] ),
    .B(_0339_),
    .Y(_0213_));
 sky130_fd_sc_hd__inv_2 _1521_ (.A(_0213_),
    .Y(_0214_));
 sky130_fd_sc_hd__o21a_1 _1522_ (.A1(net208),
    .A2(_0353_),
    .B1(_0214_),
    .X(_0215_));
 sky130_fd_sc_hd__a21oi_1 _1523_ (.A1(\state[8] ),
    .A2(_0350_),
    .B1(_0351_),
    .Y(_0216_));
 sky130_fd_sc_hd__nand3b_2 _1524_ (.A_N(_0216_),
    .B(_0206_),
    .C(_0342_),
    .Y(_0217_));
 sky130_fd_sc_hd__nand2_1 _1525_ (.A(_0217_),
    .B(net208),
    .Y(_0218_));
 sky130_fd_sc_hd__o21ai_1 _1526_ (.A1(_0215_),
    .A2(_0217_),
    .B1(net209),
    .Y(_0144_));
 sky130_fd_sc_hd__nand2_1 _1527_ (.A(net186),
    .B(\latency_count[0] ),
    .Y(_0219_));
 sky130_fd_sc_hd__a21o_1 _1528_ (.A1(_0316_),
    .A2(_0219_),
    .B1(_0358_),
    .X(_0220_));
 sky130_fd_sc_hd__a21o_1 _1529_ (.A1(_0214_),
    .A2(_0220_),
    .B1(_0217_),
    .X(_0221_));
 sky130_fd_sc_hd__nand2_1 _1530_ (.A(_0217_),
    .B(net186),
    .Y(_0222_));
 sky130_fd_sc_hd__nand2_1 _1531_ (.A(_0221_),
    .B(net187),
    .Y(_0145_));
 sky130_fd_sc_hd__nand2_1 _1532_ (.A(_0316_),
    .B(net189),
    .Y(_0223_));
 sky130_fd_sc_hd__a21o_1 _1533_ (.A1(_0354_),
    .A2(_0223_),
    .B1(_0213_),
    .X(_0224_));
 sky130_fd_sc_hd__nand2_1 _1534_ (.A(_0217_),
    .B(net189),
    .Y(_0225_));
 sky130_fd_sc_hd__o21ai_1 _1535_ (.A1(_0224_),
    .A2(_0217_),
    .B1(net190),
    .Y(_0146_));
 sky130_fd_sc_hd__o21ai_1 _1536_ (.A1(_0379_),
    .A2(\state[1] ),
    .B1(_0368_),
    .Y(_0226_));
 sky130_fd_sc_hd__nand2_1 _1537_ (.A(_0226_),
    .B(net345),
    .Y(_0227_));
 sky130_fd_sc_hd__or2b_1 _1538_ (.A(net345),
    .B_N(_0368_),
    .X(_0228_));
 sky130_fd_sc_hd__and2_1 _1539_ (.A(net346),
    .B(_0228_),
    .X(_0229_));
 sky130_fd_sc_hd__clkbuf_1 _1540_ (.A(net347),
    .X(_0147_));
 sky130_fd_sc_hd__nand2_1 _1541_ (.A(\read_word[0] ),
    .B(net242),
    .Y(_0230_));
 sky130_fd_sc_hd__inv_2 _1542_ (.A(_0230_),
    .Y(_0231_));
 sky130_fd_sc_hd__o21ai_1 _1543_ (.A1(_0372_),
    .A2(_0231_),
    .B1(_0226_),
    .Y(_0232_));
 sky130_fd_sc_hd__a21boi_1 _1544_ (.A1(_0367_),
    .A2(_0227_),
    .B1_N(_0232_),
    .Y(_0148_));
 sky130_fd_sc_hd__nor2_1 _1545_ (.A(net228),
    .B(_0372_),
    .Y(_0233_));
 sky130_fd_sc_hd__a22o_1 _1546_ (.A1(_0231_),
    .A2(_0233_),
    .B1(_0232_),
    .B2(net228),
    .X(_0149_));
 sky130_fd_sc_hd__nand2_1 _1547_ (.A(_0501_),
    .B(\state[5] ),
    .Y(_0234_));
 sky130_fd_sc_hd__o211a_1 _1548_ (.A1(_0330_),
    .A2(_0324_),
    .B1(_0197_),
    .C1(_0384_),
    .X(_0235_));
 sky130_fd_sc_hd__nand2_2 _1549_ (.A(_0361_),
    .B(_0235_),
    .Y(_0236_));
 sky130_fd_sc_hd__nand2_1 _1550_ (.A(_0236_),
    .B(net329),
    .Y(_0237_));
 sky130_fd_sc_hd__o21ai_1 _1551_ (.A1(_0234_),
    .A2(_0236_),
    .B1(net330),
    .Y(_0150_));
 sky130_fd_sc_hd__or3b_1 _1552_ (.A(_0304_),
    .B(_0552_),
    .C_N(_0308_),
    .X(_0238_));
 sky130_fd_sc_hd__nand2_1 _1553_ (.A(_0236_),
    .B(net332),
    .Y(_0239_));
 sky130_fd_sc_hd__o21ai_1 _1554_ (.A1(_0238_),
    .A2(_0236_),
    .B1(net333),
    .Y(_0151_));
 sky130_fd_sc_hd__nand2_1 _1555_ (.A(_0309_),
    .B(_0543_),
    .Y(_0240_));
 sky130_fd_sc_hd__nand2_1 _1556_ (.A(_0308_),
    .B(net214),
    .Y(_0241_));
 sky130_fd_sc_hd__a21o_1 _1557_ (.A1(_0240_),
    .A2(_0241_),
    .B1(_0304_),
    .X(_0242_));
 sky130_fd_sc_hd__nand2_1 _1558_ (.A(_0236_),
    .B(net214),
    .Y(_0243_));
 sky130_fd_sc_hd__o21ai_1 _1559_ (.A1(_0242_),
    .A2(_0236_),
    .B1(net215),
    .Y(_0152_));
 sky130_fd_sc_hd__dfstp_1 _1560_ (.CLK(clknet_3_6__leaf_clk_i),
    .D(net204),
    .SET_B(net106),
    .Q(\state[0] ));
 sky130_fd_sc_hd__dfrtp_2 _1561_ (.CLK(clknet_3_6__leaf_clk_i),
    .D(_0001_),
    .RESET_B(net106),
    .Q(\state[1] ));
 sky130_fd_sc_hd__dfrtp_4 _1562_ (.CLK(clknet_3_7__leaf_clk_i),
    .D(net185),
    .RESET_B(net106),
    .Q(\state[2] ));
 sky130_fd_sc_hd__dfrtp_1 _1563_ (.CLK(clknet_3_6__leaf_clk_i),
    .D(_0005_),
    .RESET_B(net106),
    .Q(\state[3] ));
 sky130_fd_sc_hd__dfrtp_1 _1564_ (.CLK(clknet_3_6__leaf_clk_i),
    .D(net111),
    .RESET_B(net106),
    .Q(\state[4] ));
 sky130_fd_sc_hd__dfrtp_1 _1565_ (.CLK(clknet_3_6__leaf_clk_i),
    .D(net341),
    .RESET_B(net107),
    .Q(\state[5] ));
 sky130_fd_sc_hd__dfrtp_1 _1566_ (.CLK(clknet_3_3__leaf_clk_i),
    .D(net328),
    .RESET_B(net106),
    .Q(\state[6] ));
 sky130_fd_sc_hd__dfrtp_1 _1567_ (.CLK(clknet_3_6__leaf_clk_i),
    .D(_0002_),
    .RESET_B(net106),
    .Q(\state[7] ));
 sky130_fd_sc_hd__dfrtp_2 _1568_ (.CLK(clknet_3_1__leaf_clk_i),
    .D(_0010_),
    .RESET_B(net107),
    .Q(\state[8] ));
 sky130_fd_sc_hd__dfrtp_4 _1569_ (.CLK(clknet_3_6__leaf_clk_i),
    .D(net338),
    .RESET_B(net106),
    .Q(\state[9] ));
 sky130_fd_sc_hd__dfrtp_1 _1570_ (.CLK(clknet_3_6__leaf_clk_i),
    .D(net112),
    .RESET_B(net106),
    .Q(\state[10] ));
 sky130_fd_sc_hd__dfrtp_2 _1571_ (.CLK(clknet_3_6__leaf_clk_i),
    .D(net288),
    .RESET_B(net106),
    .Q(\state[11] ));
 sky130_fd_sc_hd__dfrtp_1 _1572_ (.CLK(clknet_3_4__leaf_clk_i),
    .D(net336),
    .RESET_B(net107),
    .Q(\write_word[0] ));
 sky130_fd_sc_hd__dfrtp_1 _1573_ (.CLK(clknet_3_4__leaf_clk_i),
    .D(net202),
    .RESET_B(net107),
    .Q(\write_word[1] ));
 sky130_fd_sc_hd__dfrtp_1 _1574_ (.CLK(clknet_3_4__leaf_clk_i),
    .D(net207),
    .RESET_B(net107),
    .Q(\write_word[2] ));
 sky130_fd_sc_hd__dfrtp_2 _1575_ (.CLK(clknet_3_7__leaf_clk_i),
    .D(net320),
    .RESET_B(net106),
    .Q(\current_nibble[1] ));
 sky130_fd_sc_hd__dfrtp_1 _1576_ (.CLK(clknet_3_6__leaf_clk_i),
    .D(net221),
    .RESET_B(net106),
    .Q(\current_nibble[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1577_ (.CLK(net103),
    .D(_0034_),
    .Q(\read_buf[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1578_ (.CLK(net103),
    .D(_0035_),
    .Q(\read_buf[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1579_ (.CLK(net103),
    .D(_0036_),
    .Q(\read_buf[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1580_ (.CLK(net103),
    .D(_0037_),
    .Q(\read_buf[3] ));
 sky130_fd_sc_hd__dfxtp_1 _1581_ (.CLK(net103),
    .D(_0038_),
    .Q(\read_buf[8] ));
 sky130_fd_sc_hd__dfxtp_1 _1582_ (.CLK(net2),
    .D(_0039_),
    .Q(\read_buf[9] ));
 sky130_fd_sc_hd__dfxtp_1 _1583_ (.CLK(net2),
    .D(_0040_),
    .Q(\read_buf[10] ));
 sky130_fd_sc_hd__dfxtp_1 _1584_ (.CLK(net2),
    .D(_0041_),
    .Q(\read_buf[11] ));
 sky130_fd_sc_hd__dfxtp_1 _1585_ (.CLK(net103),
    .D(_0042_),
    .Q(\read_buf[16] ));
 sky130_fd_sc_hd__dfxtp_1 _1586_ (.CLK(net103),
    .D(_0043_),
    .Q(\read_buf[17] ));
 sky130_fd_sc_hd__dfxtp_1 _1587_ (.CLK(net103),
    .D(_0044_),
    .Q(\read_buf[18] ));
 sky130_fd_sc_hd__dfxtp_1 _1588_ (.CLK(net103),
    .D(_0045_),
    .Q(\read_buf[19] ));
 sky130_fd_sc_hd__dfxtp_1 _1589_ (.CLK(net103),
    .D(_0046_),
    .Q(\read_buf[24] ));
 sky130_fd_sc_hd__dfxtp_1 _1590_ (.CLK(net103),
    .D(_0047_),
    .Q(\read_buf[25] ));
 sky130_fd_sc_hd__dfxtp_1 _1591_ (.CLK(net103),
    .D(_0048_),
    .Q(\read_buf[26] ));
 sky130_fd_sc_hd__dfxtp_1 _1592_ (.CLK(net103),
    .D(_0049_),
    .Q(\read_buf[27] ));
 sky130_fd_sc_hd__dfxtp_1 _1593_ (.CLK(net103),
    .D(_0050_),
    .Q(\read_byte[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1594_ (.CLK(net2),
    .D(_0051_),
    .Q(\read_byte[1] ));
 sky130_fd_sc_hd__dfxtp_2 _1595_ (.CLK(net2),
    .D(_0052_),
    .Q(\read_byte[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1596_ (.CLK(net2),
    .D(_0053_),
    .Q(word_ready));
 sky130_fd_sc_hd__dfrtp_4 _1597_ (.CLK(net109),
    .D(_0000_),
    .RESET_B(net107),
    .Q(net63));
 sky130_fd_sc_hd__dfxtp_1 _1598_ (.CLK(_0013_),
    .D(_0054_),
    .Q(\read_buf[4] ));
 sky130_fd_sc_hd__dfxtp_1 _1599_ (.CLK(_0014_),
    .D(_0055_),
    .Q(\read_buf[5] ));
 sky130_fd_sc_hd__dfxtp_1 _1600_ (.CLK(_0015_),
    .D(_0056_),
    .Q(\read_buf[6] ));
 sky130_fd_sc_hd__dfxtp_1 _1601_ (.CLK(_0016_),
    .D(_0057_),
    .Q(\read_buf[7] ));
 sky130_fd_sc_hd__dfxtp_1 _1602_ (.CLK(_0017_),
    .D(_0058_),
    .Q(\read_buf[12] ));
 sky130_fd_sc_hd__dfxtp_1 _1603_ (.CLK(_0018_),
    .D(_0059_),
    .Q(\read_buf[13] ));
 sky130_fd_sc_hd__dfxtp_1 _1604_ (.CLK(_0019_),
    .D(_0060_),
    .Q(\read_buf[14] ));
 sky130_fd_sc_hd__dfxtp_1 _1605_ (.CLK(_0020_),
    .D(_0061_),
    .Q(\read_buf[15] ));
 sky130_fd_sc_hd__dfxtp_1 _1606_ (.CLK(_0021_),
    .D(_0062_),
    .Q(\read_buf[20] ));
 sky130_fd_sc_hd__dfxtp_1 _1607_ (.CLK(_0022_),
    .D(_0063_),
    .Q(\read_buf[21] ));
 sky130_fd_sc_hd__dfxtp_1 _1608_ (.CLK(_0023_),
    .D(_0064_),
    .Q(\read_buf[22] ));
 sky130_fd_sc_hd__dfxtp_1 _1609_ (.CLK(_0024_),
    .D(_0065_),
    .Q(\read_buf[23] ));
 sky130_fd_sc_hd__dfxtp_1 _1610_ (.CLK(_0025_),
    .D(_0066_),
    .Q(\read_buf[28] ));
 sky130_fd_sc_hd__dfxtp_1 _1611_ (.CLK(_0026_),
    .D(_0067_),
    .Q(\read_buf[29] ));
 sky130_fd_sc_hd__dfxtp_1 _1612_ (.CLK(_0027_),
    .D(_0068_),
    .Q(\read_buf[30] ));
 sky130_fd_sc_hd__dfxtp_1 _1613_ (.CLK(_0028_),
    .D(_0069_),
    .Q(\read_buf[31] ));
 sky130_fd_sc_hd__dfrtp_2 _1614_ (.CLK(clknet_3_0__leaf_clk_i),
    .D(net315),
    .RESET_B(net104),
    .Q(net69));
 sky130_fd_sc_hd__dfrtp_2 _1615_ (.CLK(clknet_3_0__leaf_clk_i),
    .D(net273),
    .RESET_B(net104),
    .Q(net80));
 sky130_fd_sc_hd__dfrtp_2 _1616_ (.CLK(clknet_3_0__leaf_clk_i),
    .D(net297),
    .RESET_B(net104),
    .Q(net91));
 sky130_fd_sc_hd__dfrtp_2 _1617_ (.CLK(clknet_3_1__leaf_clk_i),
    .D(net312),
    .RESET_B(net104),
    .Q(net96));
 sky130_fd_sc_hd__dfrtp_2 _1618_ (.CLK(clknet_3_1__leaf_clk_i),
    .D(net282),
    .RESET_B(net104),
    .Q(net97));
 sky130_fd_sc_hd__dfrtp_1 _1619_ (.CLK(clknet_3_0__leaf_clk_i),
    .D(net306),
    .RESET_B(net104),
    .Q(net98));
 sky130_fd_sc_hd__dfrtp_1 _1620_ (.CLK(clknet_3_0__leaf_clk_i),
    .D(net213),
    .RESET_B(net104),
    .Q(net99));
 sky130_fd_sc_hd__dfrtp_2 _1621_ (.CLK(clknet_3_1__leaf_clk_i),
    .D(net264),
    .RESET_B(net104),
    .Q(net100));
 sky130_fd_sc_hd__dfrtp_1 _1622_ (.CLK(clknet_3_0__leaf_clk_i),
    .D(net303),
    .RESET_B(net104),
    .Q(net101));
 sky130_fd_sc_hd__dfrtp_1 _1623_ (.CLK(clknet_3_0__leaf_clk_i),
    .D(net219),
    .RESET_B(net104),
    .Q(net102));
 sky130_fd_sc_hd__dfrtp_1 _1624_ (.CLK(clknet_3_0__leaf_clk_i),
    .D(net252),
    .RESET_B(net104),
    .Q(net70));
 sky130_fd_sc_hd__dfrtp_1 _1625_ (.CLK(clknet_3_0__leaf_clk_i),
    .D(net227),
    .RESET_B(net104),
    .Q(net71));
 sky130_fd_sc_hd__dfrtp_1 _1626_ (.CLK(clknet_3_0__leaf_clk_i),
    .D(net249),
    .RESET_B(net104),
    .Q(net72));
 sky130_fd_sc_hd__dfrtp_1 _1627_ (.CLK(clknet_3_0__leaf_clk_i),
    .D(net224),
    .RESET_B(net104),
    .Q(net73));
 sky130_fd_sc_hd__dfrtp_1 _1628_ (.CLK(clknet_3_0__leaf_clk_i),
    .D(net238),
    .RESET_B(net104),
    .Q(net74));
 sky130_fd_sc_hd__dfrtp_1 _1629_ (.CLK(clknet_3_2__leaf_clk_i),
    .D(net255),
    .RESET_B(net104),
    .Q(net75));
 sky130_fd_sc_hd__dfrtp_1 _1630_ (.CLK(clknet_3_2__leaf_clk_i),
    .D(net246),
    .RESET_B(net105),
    .Q(net76));
 sky130_fd_sc_hd__dfrtp_1 _1631_ (.CLK(clknet_3_3__leaf_clk_i),
    .D(net235),
    .RESET_B(net105),
    .Q(net77));
 sky130_fd_sc_hd__dfrtp_1 _1632_ (.CLK(clknet_3_2__leaf_clk_i),
    .D(net258),
    .RESET_B(net105),
    .Q(net78));
 sky130_fd_sc_hd__dfrtp_1 _1633_ (.CLK(clknet_3_2__leaf_clk_i),
    .D(net232),
    .RESET_B(net105),
    .Q(net79));
 sky130_fd_sc_hd__dfrtp_1 _1634_ (.CLK(clknet_3_2__leaf_clk_i),
    .D(net276),
    .RESET_B(net105),
    .Q(net81));
 sky130_fd_sc_hd__dfrtp_1 _1635_ (.CLK(clknet_3_2__leaf_clk_i),
    .D(net261),
    .RESET_B(net105),
    .Q(net82));
 sky130_fd_sc_hd__dfrtp_1 _1636_ (.CLK(clknet_3_2__leaf_clk_i),
    .D(net294),
    .RESET_B(net105),
    .Q(net83));
 sky130_fd_sc_hd__dfrtp_1 _1637_ (.CLK(clknet_3_2__leaf_clk_i),
    .D(net279),
    .RESET_B(net105),
    .Q(net84));
 sky130_fd_sc_hd__dfrtp_2 _1638_ (.CLK(clknet_3_2__leaf_clk_i),
    .D(net241),
    .RESET_B(net105),
    .Q(net85));
 sky130_fd_sc_hd__dfrtp_1 _1639_ (.CLK(clknet_3_2__leaf_clk_i),
    .D(net318),
    .RESET_B(net105),
    .Q(net86));
 sky130_fd_sc_hd__dfrtp_2 _1640_ (.CLK(clknet_3_2__leaf_clk_i),
    .D(net270),
    .RESET_B(net105),
    .Q(net87));
 sky130_fd_sc_hd__dfrtp_2 _1641_ (.CLK(clknet_3_3__leaf_clk_i),
    .D(net291),
    .RESET_B(net105),
    .Q(net88));
 sky130_fd_sc_hd__dfrtp_2 _1642_ (.CLK(clknet_3_3__leaf_clk_i),
    .D(net300),
    .RESET_B(net105),
    .Q(net89));
 sky130_fd_sc_hd__dfrtp_2 _1643_ (.CLK(clknet_3_2__leaf_clk_i),
    .D(net285),
    .RESET_B(net105),
    .Q(net90));
 sky130_fd_sc_hd__dfrtp_2 _1644_ (.CLK(clknet_3_2__leaf_clk_i),
    .D(net309),
    .RESET_B(net105),
    .Q(net92));
 sky130_fd_sc_hd__dfrtp_4 _1645_ (.CLK(clknet_3_3__leaf_clk_i),
    .D(net326),
    .RESET_B(net105),
    .Q(net93));
 sky130_fd_sc_hd__dfrtp_4 _1646_ (.CLK(clknet_3_3__leaf_clk_i),
    .D(_0102_),
    .RESET_B(net106),
    .Q(net95));
 sky130_fd_sc_hd__dfxtp_2 _1647_ (.CLK(clknet_3_4__leaf_clk_i),
    .D(net267),
    .Q(net65));
 sky130_fd_sc_hd__dfxtp_1 _1648_ (.CLK(clknet_3_4__leaf_clk_i),
    .D(net196),
    .Q(net66));
 sky130_fd_sc_hd__dfxtp_1 _1649_ (.CLK(clknet_3_4__leaf_clk_i),
    .D(net323),
    .Q(net67));
 sky130_fd_sc_hd__dfxtp_1 _1650_ (.CLK(clknet_3_4__leaf_clk_i),
    .D(net199),
    .Q(net68));
 sky130_fd_sc_hd__dfxtp_1 _1651_ (.CLK(clknet_3_4__leaf_clk_i),
    .D(_0107_),
    .Q(\write_buf[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1652_ (.CLK(clknet_3_5__leaf_clk_i),
    .D(_0108_),
    .Q(\write_buf[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1653_ (.CLK(clknet_3_4__leaf_clk_i),
    .D(_0109_),
    .Q(\write_buf[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1654_ (.CLK(clknet_3_5__leaf_clk_i),
    .D(_0110_),
    .Q(\write_buf[3] ));
 sky130_fd_sc_hd__dfxtp_1 _1655_ (.CLK(clknet_3_4__leaf_clk_i),
    .D(_0111_),
    .Q(\write_buf[4] ));
 sky130_fd_sc_hd__dfxtp_1 _1656_ (.CLK(clknet_3_5__leaf_clk_i),
    .D(_0112_),
    .Q(\write_buf[5] ));
 sky130_fd_sc_hd__dfxtp_1 _1657_ (.CLK(clknet_3_4__leaf_clk_i),
    .D(_0113_),
    .Q(\write_buf[6] ));
 sky130_fd_sc_hd__dfxtp_1 _1658_ (.CLK(clknet_3_5__leaf_clk_i),
    .D(_0114_),
    .Q(\write_buf[7] ));
 sky130_fd_sc_hd__dfxtp_1 _1659_ (.CLK(clknet_3_5__leaf_clk_i),
    .D(_0115_),
    .Q(\write_buf[8] ));
 sky130_fd_sc_hd__dfxtp_1 _1660_ (.CLK(clknet_3_5__leaf_clk_i),
    .D(_0116_),
    .Q(\write_buf[9] ));
 sky130_fd_sc_hd__dfxtp_1 _1661_ (.CLK(clknet_3_5__leaf_clk_i),
    .D(_0117_),
    .Q(\write_buf[10] ));
 sky130_fd_sc_hd__dfxtp_1 _1662_ (.CLK(clknet_3_5__leaf_clk_i),
    .D(_0118_),
    .Q(\write_buf[11] ));
 sky130_fd_sc_hd__dfxtp_1 _1663_ (.CLK(clknet_3_5__leaf_clk_i),
    .D(_0119_),
    .Q(\write_buf[12] ));
 sky130_fd_sc_hd__dfxtp_1 _1664_ (.CLK(clknet_3_5__leaf_clk_i),
    .D(_0120_),
    .Q(\write_buf[13] ));
 sky130_fd_sc_hd__dfxtp_1 _1665_ (.CLK(clknet_3_5__leaf_clk_i),
    .D(_0121_),
    .Q(\write_buf[14] ));
 sky130_fd_sc_hd__dfxtp_1 _1666_ (.CLK(clknet_3_5__leaf_clk_i),
    .D(_0122_),
    .Q(\write_buf[15] ));
 sky130_fd_sc_hd__dfxtp_1 _1667_ (.CLK(clknet_3_5__leaf_clk_i),
    .D(_0123_),
    .Q(\write_buf[16] ));
 sky130_fd_sc_hd__dfxtp_1 _1668_ (.CLK(clknet_3_5__leaf_clk_i),
    .D(_0124_),
    .Q(\write_buf[17] ));
 sky130_fd_sc_hd__dfxtp_1 _1669_ (.CLK(clknet_3_5__leaf_clk_i),
    .D(_0125_),
    .Q(\write_buf[18] ));
 sky130_fd_sc_hd__dfxtp_1 _1670_ (.CLK(clknet_3_7__leaf_clk_i),
    .D(_0126_),
    .Q(\write_buf[19] ));
 sky130_fd_sc_hd__dfxtp_1 _1671_ (.CLK(clknet_3_5__leaf_clk_i),
    .D(_0127_),
    .Q(\write_buf[20] ));
 sky130_fd_sc_hd__dfxtp_1 _1672_ (.CLK(clknet_3_7__leaf_clk_i),
    .D(_0128_),
    .Q(\write_buf[21] ));
 sky130_fd_sc_hd__dfxtp_1 _1673_ (.CLK(clknet_3_7__leaf_clk_i),
    .D(_0129_),
    .Q(\write_buf[22] ));
 sky130_fd_sc_hd__dfxtp_1 _1674_ (.CLK(clknet_3_7__leaf_clk_i),
    .D(_0130_),
    .Q(\write_buf[23] ));
 sky130_fd_sc_hd__dfxtp_1 _1675_ (.CLK(clknet_3_7__leaf_clk_i),
    .D(_0131_),
    .Q(\write_buf[24] ));
 sky130_fd_sc_hd__dfxtp_1 _1676_ (.CLK(clknet_3_7__leaf_clk_i),
    .D(_0132_),
    .Q(\write_buf[25] ));
 sky130_fd_sc_hd__dfxtp_1 _1677_ (.CLK(clknet_3_7__leaf_clk_i),
    .D(_0133_),
    .Q(\write_buf[26] ));
 sky130_fd_sc_hd__dfxtp_1 _1678_ (.CLK(clknet_3_7__leaf_clk_i),
    .D(_0134_),
    .Q(\write_buf[27] ));
 sky130_fd_sc_hd__dfxtp_1 _1679_ (.CLK(clknet_3_7__leaf_clk_i),
    .D(_0135_),
    .Q(\write_buf[28] ));
 sky130_fd_sc_hd__dfxtp_1 _1680_ (.CLK(clknet_3_7__leaf_clk_i),
    .D(_0136_),
    .Q(\write_buf[29] ));
 sky130_fd_sc_hd__dfxtp_1 _1681_ (.CLK(clknet_3_7__leaf_clk_i),
    .D(_0137_),
    .Q(\write_buf[30] ));
 sky130_fd_sc_hd__dfxtp_1 _1682_ (.CLK(clknet_3_7__leaf_clk_i),
    .D(_0138_),
    .Q(\write_buf[31] ));
 sky130_fd_sc_hd__dfrtp_1 _1683_ (.CLK(clknet_3_7__leaf_clk_i),
    .D(net182),
    .RESET_B(net107),
    .Q(clock_enable));
 sky130_fd_sc_hd__dfrtp_1 _1684_ (.CLK(clknet_3_7__leaf_clk_i),
    .D(_0140_),
    .RESET_B(net107),
    .Q(\current_nibble[0] ));
 sky130_fd_sc_hd__dfrtp_1 _1685_ (.CLK(clknet_3_3__leaf_clk_i),
    .D(_0141_),
    .RESET_B(net1),
    .Q(\pre_cycle[0] ));
 sky130_fd_sc_hd__dfrtp_1 _1686_ (.CLK(clknet_3_6__leaf_clk_i),
    .D(net193),
    .RESET_B(net106),
    .Q(\pre_cycle[1] ));
 sky130_fd_sc_hd__dfrtp_1 _1687_ (.CLK(clknet_3_3__leaf_clk_i),
    .D(net179),
    .RESET_B(net1),
    .Q(current_dqsm));
 sky130_fd_sc_hd__dfrtp_1 _1688_ (.CLK(clknet_3_1__leaf_clk_i),
    .D(net210),
    .RESET_B(net1),
    .Q(\latency_count[0] ));
 sky130_fd_sc_hd__dfrtp_1 _1689_ (.CLK(clknet_3_1__leaf_clk_i),
    .D(net188),
    .RESET_B(net1),
    .Q(\latency_count[1] ));
 sky130_fd_sc_hd__dfrtp_1 _1690_ (.CLK(clknet_3_1__leaf_clk_i),
    .D(net191),
    .RESET_B(net107),
    .Q(\latency_count[2] ));
 sky130_fd_sc_hd__dfrtp_1 _1691_ (.CLK(clknet_3_6__leaf_clk_i),
    .D(_0147_),
    .RESET_B(net106),
    .Q(\read_word[0] ));
 sky130_fd_sc_hd__dfrtp_1 _1692_ (.CLK(clknet_3_6__leaf_clk_i),
    .D(net243),
    .RESET_B(net106),
    .Q(\read_word[1] ));
 sky130_fd_sc_hd__dfrtp_1 _1693_ (.CLK(clknet_3_6__leaf_clk_i),
    .D(net229),
    .RESET_B(net107),
    .Q(\read_word[2] ));
 sky130_fd_sc_hd__dfrtp_1 _1694_ (.CLK(clknet_3_7__leaf_clk_i),
    .D(net331),
    .RESET_B(net107),
    .Q(\write_byte[0] ));
 sky130_fd_sc_hd__dfrtp_1 _1695_ (.CLK(clknet_3_5__leaf_clk_i),
    .D(net334),
    .RESET_B(net107),
    .Q(\write_byte[1] ));
 sky130_fd_sc_hd__dfrtp_1 _1696_ (.CLK(clknet_3_4__leaf_clk_i),
    .D(net216),
    .RESET_B(net107),
    .Q(\write_byte[2] ));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk_i (.A(clk_i),
    .X(clknet_0_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_0__f_clk_i (.A(clknet_0_clk_i),
    .X(clknet_3_0__leaf_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_1__f_clk_i (.A(clknet_0_clk_i),
    .X(clknet_3_1__leaf_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_2__f_clk_i (.A(clknet_0_clk_i),
    .X(clknet_3_2__leaf_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_3__f_clk_i (.A(clknet_0_clk_i),
    .X(clknet_3_3__leaf_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_4__f_clk_i (.A(clknet_0_clk_i),
    .X(clknet_3_4__leaf_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_5__f_clk_i (.A(clknet_0_clk_i),
    .X(clknet_3_5__leaf_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_6__f_clk_i (.A(clknet_0_clk_i),
    .X(clknet_3_6__leaf_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_7__f_clk_i (.A(clknet_0_clk_i),
    .X(clknet_3_7__leaf_clk_i));
 sky130_fd_sc_hd__buf_4 fanout103 (.A(net2),
    .X(net103));
 sky130_fd_sc_hd__clkbuf_8 fanout104 (.A(net1),
    .X(net104));
 sky130_fd_sc_hd__clkbuf_8 fanout105 (.A(net1),
    .X(net105));
 sky130_fd_sc_hd__clkbuf_8 fanout106 (.A(net107),
    .X(net106));
 sky130_fd_sc_hd__buf_6 fanout107 (.A(net1),
    .X(net107));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1 (.A(\state[7] ),
    .X(net110));
 sky130_fd_sc_hd__dlygate4sd3_1 hold10 (.A(\write_buf[31] ),
    .X(net119));
 sky130_fd_sc_hd__dlygate4sd3_1 hold100 (.A(_0218_),
    .X(net209));
 sky130_fd_sc_hd__dlygate4sd3_1 hold101 (.A(_0144_),
    .X(net210));
 sky130_fd_sc_hd__dlygate4sd3_1 hold102 (.A(net99),
    .X(net211));
 sky130_fd_sc_hd__dlygate4sd3_1 hold103 (.A(_0446_),
    .X(net212));
 sky130_fd_sc_hd__dlygate4sd3_1 hold104 (.A(_0076_),
    .X(net213));
 sky130_fd_sc_hd__buf_1 hold105 (.A(\write_byte[2] ),
    .X(net214));
 sky130_fd_sc_hd__dlygate4sd3_1 hold106 (.A(_0243_),
    .X(net215));
 sky130_fd_sc_hd__dlygate4sd3_1 hold107 (.A(_0152_),
    .X(net216));
 sky130_fd_sc_hd__dlygate4sd3_1 hold108 (.A(net102),
    .X(net217));
 sky130_fd_sc_hd__dlygate4sd3_1 hold109 (.A(_0454_),
    .X(net218));
 sky130_fd_sc_hd__dlygate4sd3_1 hold11 (.A(_0193_),
    .X(net120));
 sky130_fd_sc_hd__dlygate4sd3_1 hold110 (.A(_0079_),
    .X(net219));
 sky130_fd_sc_hd__buf_1 hold111 (.A(\current_nibble[2] ),
    .X(net220));
 sky130_fd_sc_hd__dlygate4sd3_1 hold112 (.A(_0033_),
    .X(net221));
 sky130_fd_sc_hd__dlygate4sd3_1 hold113 (.A(net73),
    .X(net222));
 sky130_fd_sc_hd__dlygate4sd3_1 hold114 (.A(_0462_),
    .X(net223));
 sky130_fd_sc_hd__dlygate4sd3_1 hold115 (.A(_0083_),
    .X(net224));
 sky130_fd_sc_hd__dlygate4sd3_1 hold116 (.A(net71),
    .X(net225));
 sky130_fd_sc_hd__dlygate4sd3_1 hold117 (.A(_0458_),
    .X(net226));
 sky130_fd_sc_hd__dlygate4sd3_1 hold118 (.A(_0081_),
    .X(net227));
 sky130_fd_sc_hd__buf_1 hold119 (.A(\read_word[2] ),
    .X(net228));
 sky130_fd_sc_hd__dlygate4sd3_1 hold12 (.A(\write_buf[4] ),
    .X(net121));
 sky130_fd_sc_hd__dlygate4sd3_1 hold120 (.A(_0149_),
    .X(net229));
 sky130_fd_sc_hd__dlygate4sd3_1 hold121 (.A(net79),
    .X(net230));
 sky130_fd_sc_hd__dlygate4sd3_1 hold122 (.A(_0476_),
    .X(net231));
 sky130_fd_sc_hd__dlygate4sd3_1 hold123 (.A(_0089_),
    .X(net232));
 sky130_fd_sc_hd__dlygate4sd3_1 hold124 (.A(net77),
    .X(net233));
 sky130_fd_sc_hd__dlygate4sd3_1 hold125 (.A(_0472_),
    .X(net234));
 sky130_fd_sc_hd__dlygate4sd3_1 hold126 (.A(_0087_),
    .X(net235));
 sky130_fd_sc_hd__dlygate4sd3_1 hold127 (.A(net74),
    .X(net236));
 sky130_fd_sc_hd__dlygate4sd3_1 hold128 (.A(_0464_),
    .X(net237));
 sky130_fd_sc_hd__dlygate4sd3_1 hold129 (.A(_0084_),
    .X(net238));
 sky130_fd_sc_hd__dlygate4sd3_1 hold13 (.A(_0156_),
    .X(net122));
 sky130_fd_sc_hd__dlygate4sd3_1 hold130 (.A(net85),
    .X(net239));
 sky130_fd_sc_hd__dlygate4sd3_1 hold131 (.A(_0486_),
    .X(net240));
 sky130_fd_sc_hd__dlygate4sd3_1 hold132 (.A(_0094_),
    .X(net241));
 sky130_fd_sc_hd__dlygate4sd3_1 hold133 (.A(\read_word[1] ),
    .X(net242));
 sky130_fd_sc_hd__dlygate4sd3_1 hold134 (.A(_0148_),
    .X(net243));
 sky130_fd_sc_hd__dlygate4sd3_1 hold135 (.A(net76),
    .X(net244));
 sky130_fd_sc_hd__dlygate4sd3_1 hold136 (.A(_0470_),
    .X(net245));
 sky130_fd_sc_hd__dlygate4sd3_1 hold137 (.A(_0086_),
    .X(net246));
 sky130_fd_sc_hd__dlygate4sd3_1 hold138 (.A(net72),
    .X(net247));
 sky130_fd_sc_hd__dlygate4sd3_1 hold139 (.A(_0460_),
    .X(net248));
 sky130_fd_sc_hd__dlygate4sd3_1 hold14 (.A(\write_buf[0] ),
    .X(net123));
 sky130_fd_sc_hd__dlygate4sd3_1 hold140 (.A(_0082_),
    .X(net249));
 sky130_fd_sc_hd__dlygate4sd3_1 hold141 (.A(net70),
    .X(net250));
 sky130_fd_sc_hd__dlygate4sd3_1 hold142 (.A(_0456_),
    .X(net251));
 sky130_fd_sc_hd__dlygate4sd3_1 hold143 (.A(_0080_),
    .X(net252));
 sky130_fd_sc_hd__dlygate4sd3_1 hold144 (.A(net75),
    .X(net253));
 sky130_fd_sc_hd__dlygate4sd3_1 hold145 (.A(_0466_),
    .X(net254));
 sky130_fd_sc_hd__dlygate4sd3_1 hold146 (.A(_0085_),
    .X(net255));
 sky130_fd_sc_hd__dlygate4sd3_1 hold147 (.A(net78),
    .X(net256));
 sky130_fd_sc_hd__dlygate4sd3_1 hold148 (.A(_0474_),
    .X(net257));
 sky130_fd_sc_hd__dlygate4sd3_1 hold149 (.A(_0088_),
    .X(net258));
 sky130_fd_sc_hd__dlygate4sd3_1 hold15 (.A(_0778_),
    .X(net124));
 sky130_fd_sc_hd__dlygate4sd3_1 hold150 (.A(net82),
    .X(net259));
 sky130_fd_sc_hd__dlygate4sd3_1 hold151 (.A(_0480_),
    .X(net260));
 sky130_fd_sc_hd__dlygate4sd3_1 hold152 (.A(_0091_),
    .X(net261));
 sky130_fd_sc_hd__dlygate4sd3_1 hold153 (.A(net100),
    .X(net262));
 sky130_fd_sc_hd__dlygate4sd3_1 hold154 (.A(_0449_),
    .X(net263));
 sky130_fd_sc_hd__dlygate4sd3_1 hold155 (.A(_0077_),
    .X(net264));
 sky130_fd_sc_hd__dlygate4sd3_1 hold156 (.A(net65),
    .X(net265));
 sky130_fd_sc_hd__dlygate4sd3_1 hold157 (.A(_0575_),
    .X(net266));
 sky130_fd_sc_hd__dlygate4sd3_1 hold158 (.A(_0103_),
    .X(net267));
 sky130_fd_sc_hd__dlygate4sd3_1 hold159 (.A(net87),
    .X(net268));
 sky130_fd_sc_hd__dlygate4sd3_1 hold16 (.A(\write_buf[5] ),
    .X(net125));
 sky130_fd_sc_hd__dlygate4sd3_1 hold160 (.A(_0490_),
    .X(net269));
 sky130_fd_sc_hd__dlygate4sd3_1 hold161 (.A(_0096_),
    .X(net270));
 sky130_fd_sc_hd__dlygate4sd3_1 hold162 (.A(net80),
    .X(net271));
 sky130_fd_sc_hd__dlygate4sd3_1 hold163 (.A(_0431_),
    .X(net272));
 sky130_fd_sc_hd__dlygate4sd3_1 hold164 (.A(_0071_),
    .X(net273));
 sky130_fd_sc_hd__dlygate4sd3_1 hold165 (.A(net81),
    .X(net274));
 sky130_fd_sc_hd__dlygate4sd3_1 hold166 (.A(_0478_),
    .X(net275));
 sky130_fd_sc_hd__dlygate4sd3_1 hold167 (.A(_0090_),
    .X(net276));
 sky130_fd_sc_hd__dlygate4sd3_1 hold168 (.A(net84),
    .X(net277));
 sky130_fd_sc_hd__dlygate4sd3_1 hold169 (.A(_0484_),
    .X(net278));
 sky130_fd_sc_hd__dlygate4sd3_1 hold17 (.A(_0157_),
    .X(net126));
 sky130_fd_sc_hd__dlygate4sd3_1 hold170 (.A(_0093_),
    .X(net279));
 sky130_fd_sc_hd__dlygate4sd3_1 hold171 (.A(net97),
    .X(net280));
 sky130_fd_sc_hd__dlygate4sd3_1 hold172 (.A(_0440_),
    .X(net281));
 sky130_fd_sc_hd__dlygate4sd3_1 hold173 (.A(_0074_),
    .X(net282));
 sky130_fd_sc_hd__dlygate4sd3_1 hold174 (.A(net90),
    .X(net283));
 sky130_fd_sc_hd__dlygate4sd3_1 hold175 (.A(_0496_),
    .X(net284));
 sky130_fd_sc_hd__dlygate4sd3_1 hold176 (.A(_0099_),
    .X(net285));
 sky130_fd_sc_hd__buf_1 hold177 (.A(\state[6] ),
    .X(net286));
 sky130_fd_sc_hd__dlygate4sd3_1 hold178 (.A(_0369_),
    .X(net287));
 sky130_fd_sc_hd__dlygate4sd3_1 hold179 (.A(_0009_),
    .X(net288));
 sky130_fd_sc_hd__dlygate4sd3_1 hold18 (.A(\write_buf[14] ),
    .X(net127));
 sky130_fd_sc_hd__dlygate4sd3_1 hold180 (.A(net88),
    .X(net289));
 sky130_fd_sc_hd__dlygate4sd3_1 hold181 (.A(_0492_),
    .X(net290));
 sky130_fd_sc_hd__dlygate4sd3_1 hold182 (.A(_0097_),
    .X(net291));
 sky130_fd_sc_hd__dlygate4sd3_1 hold183 (.A(net83),
    .X(net292));
 sky130_fd_sc_hd__dlygate4sd3_1 hold184 (.A(_0482_),
    .X(net293));
 sky130_fd_sc_hd__dlygate4sd3_1 hold185 (.A(_0092_),
    .X(net294));
 sky130_fd_sc_hd__dlygate4sd3_1 hold186 (.A(net91),
    .X(net295));
 sky130_fd_sc_hd__dlygate4sd3_1 hold187 (.A(_0434_),
    .X(net296));
 sky130_fd_sc_hd__dlygate4sd3_1 hold188 (.A(_0072_),
    .X(net297));
 sky130_fd_sc_hd__dlygate4sd3_1 hold189 (.A(net89),
    .X(net298));
 sky130_fd_sc_hd__dlygate4sd3_1 hold19 (.A(_0173_),
    .X(net128));
 sky130_fd_sc_hd__dlygate4sd3_1 hold190 (.A(_0494_),
    .X(net299));
 sky130_fd_sc_hd__dlygate4sd3_1 hold191 (.A(_0098_),
    .X(net300));
 sky130_fd_sc_hd__dlygate4sd3_1 hold192 (.A(net101),
    .X(net301));
 sky130_fd_sc_hd__dlygate4sd3_1 hold193 (.A(_0452_),
    .X(net302));
 sky130_fd_sc_hd__dlygate4sd3_1 hold194 (.A(_0078_),
    .X(net303));
 sky130_fd_sc_hd__dlygate4sd3_1 hold195 (.A(net98),
    .X(net304));
 sky130_fd_sc_hd__dlygate4sd3_1 hold196 (.A(_0443_),
    .X(net305));
 sky130_fd_sc_hd__dlygate4sd3_1 hold197 (.A(_0075_),
    .X(net306));
 sky130_fd_sc_hd__dlygate4sd3_1 hold198 (.A(net92),
    .X(net307));
 sky130_fd_sc_hd__dlygate4sd3_1 hold199 (.A(_0498_),
    .X(net308));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(_0006_),
    .X(net111));
 sky130_fd_sc_hd__dlygate4sd3_1 hold20 (.A(\write_buf[24] ),
    .X(net129));
 sky130_fd_sc_hd__dlygate4sd3_1 hold200 (.A(_0100_),
    .X(net309));
 sky130_fd_sc_hd__dlygate4sd3_1 hold201 (.A(net96),
    .X(net310));
 sky130_fd_sc_hd__dlygate4sd3_1 hold202 (.A(_0437_),
    .X(net311));
 sky130_fd_sc_hd__dlygate4sd3_1 hold203 (.A(_0073_),
    .X(net312));
 sky130_fd_sc_hd__dlygate4sd3_1 hold204 (.A(net69),
    .X(net313));
 sky130_fd_sc_hd__dlygate4sd3_1 hold205 (.A(_0428_),
    .X(net314));
 sky130_fd_sc_hd__dlygate4sd3_1 hold206 (.A(_0070_),
    .X(net315));
 sky130_fd_sc_hd__dlygate4sd3_1 hold207 (.A(net86),
    .X(net316));
 sky130_fd_sc_hd__dlygate4sd3_1 hold208 (.A(_0488_),
    .X(net317));
 sky130_fd_sc_hd__dlygate4sd3_1 hold209 (.A(_0095_),
    .X(net318));
 sky130_fd_sc_hd__dlygate4sd3_1 hold21 (.A(_0186_),
    .X(net130));
 sky130_fd_sc_hd__buf_1 hold210 (.A(\current_nibble[1] ),
    .X(net319));
 sky130_fd_sc_hd__dlygate4sd3_1 hold211 (.A(_0032_),
    .X(net320));
 sky130_fd_sc_hd__dlygate4sd3_1 hold212 (.A(net67),
    .X(net321));
 sky130_fd_sc_hd__dlygate4sd3_1 hold213 (.A(_0701_),
    .X(net322));
 sky130_fd_sc_hd__dlygate4sd3_1 hold214 (.A(_0105_),
    .X(net323));
 sky130_fd_sc_hd__dlygate4sd3_1 hold215 (.A(net93),
    .X(net324));
 sky130_fd_sc_hd__dlygate4sd3_1 hold216 (.A(_0500_),
    .X(net325));
 sky130_fd_sc_hd__dlygate4sd3_1 hold217 (.A(_0101_),
    .X(net326));
 sky130_fd_sc_hd__dlygate4sd3_1 hold218 (.A(\pre_cycle[0] ),
    .X(net327));
 sky130_fd_sc_hd__dlygate4sd3_1 hold219 (.A(_0008_),
    .X(net328));
 sky130_fd_sc_hd__dlygate4sd3_1 hold22 (.A(\write_buf[20] ),
    .X(net131));
 sky130_fd_sc_hd__buf_1 hold220 (.A(\write_byte[0] ),
    .X(net329));
 sky130_fd_sc_hd__dlygate4sd3_1 hold221 (.A(_0237_),
    .X(net330));
 sky130_fd_sc_hd__dlygate4sd3_1 hold222 (.A(_0150_),
    .X(net331));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold223 (.A(\write_byte[1] ),
    .X(net332));
 sky130_fd_sc_hd__dlygate4sd3_1 hold224 (.A(_0239_),
    .X(net333));
 sky130_fd_sc_hd__dlygate4sd3_1 hold225 (.A(_0151_),
    .X(net334));
 sky130_fd_sc_hd__buf_1 hold226 (.A(\write_word[0] ),
    .X(net335));
 sky130_fd_sc_hd__dlygate4sd3_1 hold227 (.A(_0029_),
    .X(net336));
 sky130_fd_sc_hd__buf_1 hold228 (.A(\state[11] ),
    .X(net337));
 sky130_fd_sc_hd__dlygate4sd3_1 hold229 (.A(_0011_),
    .X(net338));
 sky130_fd_sc_hd__dlygate4sd3_1 hold23 (.A(_0182_),
    .X(net132));
 sky130_fd_sc_hd__clkbuf_2 hold230 (.A(\state[5] ),
    .X(net339));
 sky130_fd_sc_hd__dlygate4sd3_1 hold231 (.A(_0332_),
    .X(net340));
 sky130_fd_sc_hd__dlygate4sd3_1 hold232 (.A(_0007_),
    .X(net341));
 sky130_fd_sc_hd__dlygate4sd3_1 hold233 (.A(\current_nibble[0] ),
    .X(net342));
 sky130_fd_sc_hd__dlygate4sd3_1 hold234 (.A(net95),
    .X(net343));
 sky130_fd_sc_hd__dlygate4sd3_1 hold235 (.A(_0509_),
    .X(net344));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold236 (.A(\read_word[0] ),
    .X(net345));
 sky130_fd_sc_hd__dlygate4sd3_1 hold237 (.A(_0227_),
    .X(net346));
 sky130_fd_sc_hd__dlygate4sd3_1 hold238 (.A(_0229_),
    .X(net347));
 sky130_fd_sc_hd__dlygate4sd3_1 hold239 (.A(\state[2] ),
    .X(net348));
 sky130_fd_sc_hd__dlygate4sd3_1 hold24 (.A(\write_buf[13] ),
    .X(net133));
 sky130_fd_sc_hd__buf_1 hold240 (.A(\state[8] ),
    .X(net349));
 sky130_fd_sc_hd__dlygate4sd3_1 hold241 (.A(net63),
    .X(net350));
 sky130_fd_sc_hd__dlygate4sd3_1 hold242 (.A(\state[4] ),
    .X(net351));
 sky130_fd_sc_hd__dlygate4sd3_1 hold243 (.A(clock_enable),
    .X(net352));
 sky130_fd_sc_hd__dlygate4sd3_1 hold25 (.A(_0171_),
    .X(net134));
 sky130_fd_sc_hd__dlygate4sd3_1 hold26 (.A(\write_buf[26] ),
    .X(net135));
 sky130_fd_sc_hd__dlygate4sd3_1 hold27 (.A(_0188_),
    .X(net136));
 sky130_fd_sc_hd__dlygate4sd3_1 hold28 (.A(\write_buf[18] ),
    .X(net137));
 sky130_fd_sc_hd__dlygate4sd3_1 hold29 (.A(_0180_),
    .X(net138));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold3 (.A(net351),
    .X(net112));
 sky130_fd_sc_hd__dlygate4sd3_1 hold30 (.A(\write_buf[16] ),
    .X(net139));
 sky130_fd_sc_hd__dlygate4sd3_1 hold31 (.A(_0178_),
    .X(net140));
 sky130_fd_sc_hd__dlygate4sd3_1 hold32 (.A(\write_buf[28] ),
    .X(net141));
 sky130_fd_sc_hd__dlygate4sd3_1 hold33 (.A(_0190_),
    .X(net142));
 sky130_fd_sc_hd__dlygate4sd3_1 hold34 (.A(\write_buf[30] ),
    .X(net143));
 sky130_fd_sc_hd__dlygate4sd3_1 hold35 (.A(_0192_),
    .X(net144));
 sky130_fd_sc_hd__dlygate4sd3_1 hold36 (.A(\write_buf[2] ),
    .X(net145));
 sky130_fd_sc_hd__dlygate4sd3_1 hold37 (.A(_0154_),
    .X(net146));
 sky130_fd_sc_hd__dlygate4sd3_1 hold38 (.A(\write_buf[12] ),
    .X(net147));
 sky130_fd_sc_hd__dlygate4sd3_1 hold39 (.A(_0169_),
    .X(net148));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4 (.A(\write_buf[7] ),
    .X(net113));
 sky130_fd_sc_hd__dlygate4sd3_1 hold40 (.A(\write_buf[22] ),
    .X(net149));
 sky130_fd_sc_hd__dlygate4sd3_1 hold41 (.A(_0184_),
    .X(net150));
 sky130_fd_sc_hd__dlygate4sd3_1 hold42 (.A(\write_buf[11] ),
    .X(net151));
 sky130_fd_sc_hd__dlygate4sd3_1 hold43 (.A(_0167_),
    .X(net152));
 sky130_fd_sc_hd__dlygate4sd3_1 hold44 (.A(\write_buf[10] ),
    .X(net153));
 sky130_fd_sc_hd__dlygate4sd3_1 hold45 (.A(_0165_),
    .X(net154));
 sky130_fd_sc_hd__dlygate4sd3_1 hold46 (.A(\write_buf[9] ),
    .X(net155));
 sky130_fd_sc_hd__dlygate4sd3_1 hold47 (.A(_0163_),
    .X(net156));
 sky130_fd_sc_hd__dlygate4sd3_1 hold48 (.A(\write_buf[15] ),
    .X(net157));
 sky130_fd_sc_hd__dlygate4sd3_1 hold49 (.A(_0175_),
    .X(net158));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5 (.A(_0159_),
    .X(net114));
 sky130_fd_sc_hd__dlygate4sd3_1 hold50 (.A(\write_buf[8] ),
    .X(net159));
 sky130_fd_sc_hd__dlygate4sd3_1 hold51 (.A(_0161_),
    .X(net160));
 sky130_fd_sc_hd__dlygate4sd3_1 hold52 (.A(\write_buf[1] ),
    .X(net161));
 sky130_fd_sc_hd__dlygate4sd3_1 hold53 (.A(_0153_),
    .X(net162));
 sky130_fd_sc_hd__dlygate4sd3_1 hold54 (.A(\write_buf[27] ),
    .X(net163));
 sky130_fd_sc_hd__dlygate4sd3_1 hold55 (.A(_0189_),
    .X(net164));
 sky130_fd_sc_hd__dlygate4sd3_1 hold56 (.A(\write_buf[17] ),
    .X(net165));
 sky130_fd_sc_hd__dlygate4sd3_1 hold57 (.A(_0179_),
    .X(net166));
 sky130_fd_sc_hd__dlygate4sd3_1 hold58 (.A(\write_buf[19] ),
    .X(net167));
 sky130_fd_sc_hd__dlygate4sd3_1 hold59 (.A(_0181_),
    .X(net168));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6 (.A(\write_buf[29] ),
    .X(net115));
 sky130_fd_sc_hd__dlygate4sd3_1 hold60 (.A(\write_buf[21] ),
    .X(net169));
 sky130_fd_sc_hd__dlygate4sd3_1 hold61 (.A(_0183_),
    .X(net170));
 sky130_fd_sc_hd__dlygate4sd3_1 hold62 (.A(\write_buf[25] ),
    .X(net171));
 sky130_fd_sc_hd__dlygate4sd3_1 hold63 (.A(_0187_),
    .X(net172));
 sky130_fd_sc_hd__dlygate4sd3_1 hold64 (.A(\write_buf[23] ),
    .X(net173));
 sky130_fd_sc_hd__dlygate4sd3_1 hold65 (.A(_0185_),
    .X(net174));
 sky130_fd_sc_hd__dlygate4sd3_1 hold66 (.A(\write_buf[3] ),
    .X(net175));
 sky130_fd_sc_hd__dlygate4sd3_1 hold67 (.A(_0155_),
    .X(net176));
 sky130_fd_sc_hd__dlygate4sd3_1 hold68 (.A(current_dqsm),
    .X(net177));
 sky130_fd_sc_hd__dlygate4sd3_1 hold69 (.A(_0212_),
    .X(net178));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7 (.A(_0191_),
    .X(net116));
 sky130_fd_sc_hd__dlygate4sd3_1 hold70 (.A(_0143_),
    .X(net179));
 sky130_fd_sc_hd__dlygate4sd3_1 hold71 (.A(\state[3] ),
    .X(net180));
 sky130_fd_sc_hd__dlygate4sd3_1 hold72 (.A(_0194_),
    .X(net181));
 sky130_fd_sc_hd__dlygate4sd3_1 hold73 (.A(_0139_),
    .X(net182));
 sky130_fd_sc_hd__dlygate4sd3_1 hold74 (.A(\state[10] ),
    .X(net183));
 sky130_fd_sc_hd__dlygate4sd3_1 hold75 (.A(_0345_),
    .X(net184));
 sky130_fd_sc_hd__dlygate4sd3_1 hold76 (.A(_0004_),
    .X(net185));
 sky130_fd_sc_hd__dlygate4sd3_1 hold77 (.A(\latency_count[1] ),
    .X(net186));
 sky130_fd_sc_hd__dlygate4sd3_1 hold78 (.A(_0222_),
    .X(net187));
 sky130_fd_sc_hd__dlygate4sd3_1 hold79 (.A(_0145_),
    .X(net188));
 sky130_fd_sc_hd__dlygate4sd3_1 hold8 (.A(\write_buf[6] ),
    .X(net117));
 sky130_fd_sc_hd__dlygate4sd3_1 hold80 (.A(\latency_count[2] ),
    .X(net189));
 sky130_fd_sc_hd__dlygate4sd3_1 hold81 (.A(_0225_),
    .X(net190));
 sky130_fd_sc_hd__dlygate4sd3_1 hold82 (.A(_0146_),
    .X(net191));
 sky130_fd_sc_hd__dlygate4sd3_1 hold83 (.A(\pre_cycle[1] ),
    .X(net192));
 sky130_fd_sc_hd__dlygate4sd3_1 hold84 (.A(_0142_),
    .X(net193));
 sky130_fd_sc_hd__dlygate4sd3_1 hold85 (.A(net66),
    .X(net194));
 sky130_fd_sc_hd__dlygate4sd3_1 hold86 (.A(_0646_),
    .X(net195));
 sky130_fd_sc_hd__dlygate4sd3_1 hold87 (.A(_0104_),
    .X(net196));
 sky130_fd_sc_hd__dlygate4sd3_1 hold88 (.A(net68),
    .X(net197));
 sky130_fd_sc_hd__dlygate4sd3_1 hold89 (.A(_0772_),
    .X(net198));
 sky130_fd_sc_hd__dlygate4sd3_1 hold9 (.A(_0158_),
    .X(net118));
 sky130_fd_sc_hd__dlygate4sd3_1 hold90 (.A(_0106_),
    .X(net199));
 sky130_fd_sc_hd__buf_1 hold91 (.A(\write_word[1] ),
    .X(net200));
 sky130_fd_sc_hd__dlygate4sd3_1 hold92 (.A(_0393_),
    .X(net201));
 sky130_fd_sc_hd__dlygate4sd3_1 hold93 (.A(_0030_),
    .X(net202));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold94 (.A(\state[0] ),
    .X(net203));
 sky130_fd_sc_hd__dlygate4sd3_1 hold95 (.A(_0003_),
    .X(net204));
 sky130_fd_sc_hd__buf_1 hold96 (.A(\write_word[2] ),
    .X(net205));
 sky130_fd_sc_hd__dlygate4sd3_1 hold97 (.A(_0396_),
    .X(net206));
 sky130_fd_sc_hd__dlygate4sd3_1 hold98 (.A(_0031_),
    .X(net207));
 sky130_fd_sc_hd__dlygate4sd3_1 hold99 (.A(\latency_count[0] ),
    .X(net208));
 sky130_fd_sc_hd__clkbuf_8 input1 (.A(nrst_i),
    .X(net1));
 sky130_fd_sc_hd__buf_1 input10 (.A(sport_i[12]),
    .X(net10));
 sky130_fd_sc_hd__buf_1 input11 (.A(sport_i[13]),
    .X(net11));
 sky130_fd_sc_hd__buf_1 input12 (.A(sport_i[14]),
    .X(net12));
 sky130_fd_sc_hd__buf_1 input13 (.A(sport_i[15]),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_1 input14 (.A(sport_i[16]),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_1 input15 (.A(sport_i[17]),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_1 input16 (.A(sport_i[18]),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_1 input17 (.A(sport_i[19]),
    .X(net17));
 sky130_fd_sc_hd__buf_1 input18 (.A(sport_i[1]),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_1 input19 (.A(sport_i[20]),
    .X(net19));
 sky130_fd_sc_hd__buf_2 input2 (.A(spi_dqsm_i),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 input20 (.A(sport_i[21]),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_1 input21 (.A(sport_i[22]),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_1 input22 (.A(sport_i[23]),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_1 input23 (.A(sport_i[24]),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_1 input24 (.A(sport_i[25]),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_1 input25 (.A(sport_i[26]),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_1 input26 (.A(sport_i[27]),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_1 input27 (.A(sport_i[28]),
    .X(net27));
 sky130_fd_sc_hd__clkbuf_1 input28 (.A(sport_i[29]),
    .X(net28));
 sky130_fd_sc_hd__buf_1 input29 (.A(sport_i[2]),
    .X(net29));
 sky130_fd_sc_hd__dlymetal6s2s_1 input3 (.A(spi_miso_i[0]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_1 input30 (.A(sport_i[30]),
    .X(net30));
 sky130_fd_sc_hd__clkbuf_1 input31 (.A(sport_i[31]),
    .X(net31));
 sky130_fd_sc_hd__clkbuf_1 input32 (.A(sport_i[32]),
    .X(net32));
 sky130_fd_sc_hd__clkbuf_1 input33 (.A(sport_i[33]),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_1 input34 (.A(sport_i[34]),
    .X(net34));
 sky130_fd_sc_hd__clkbuf_1 input35 (.A(sport_i[35]),
    .X(net35));
 sky130_fd_sc_hd__clkbuf_1 input36 (.A(sport_i[36]),
    .X(net36));
 sky130_fd_sc_hd__clkbuf_1 input37 (.A(sport_i[37]),
    .X(net37));
 sky130_fd_sc_hd__clkbuf_1 input38 (.A(sport_i[38]),
    .X(net38));
 sky130_fd_sc_hd__buf_1 input39 (.A(sport_i[39]),
    .X(net39));
 sky130_fd_sc_hd__clkbuf_2 input4 (.A(spi_miso_i[1]),
    .X(net4));
 sky130_fd_sc_hd__buf_1 input40 (.A(sport_i[3]),
    .X(net40));
 sky130_fd_sc_hd__clkbuf_1 input41 (.A(sport_i[40]),
    .X(net41));
 sky130_fd_sc_hd__clkbuf_1 input42 (.A(sport_i[41]),
    .X(net42));
 sky130_fd_sc_hd__buf_1 input43 (.A(sport_i[42]),
    .X(net43));
 sky130_fd_sc_hd__buf_1 input44 (.A(sport_i[43]),
    .X(net44));
 sky130_fd_sc_hd__clkbuf_1 input45 (.A(sport_i[44]),
    .X(net45));
 sky130_fd_sc_hd__clkbuf_1 input46 (.A(sport_i[45]),
    .X(net46));
 sky130_fd_sc_hd__clkbuf_1 input47 (.A(sport_i[46]),
    .X(net47));
 sky130_fd_sc_hd__clkbuf_1 input48 (.A(sport_i[47]),
    .X(net48));
 sky130_fd_sc_hd__clkbuf_1 input49 (.A(sport_i[48]),
    .X(net49));
 sky130_fd_sc_hd__buf_2 input5 (.A(spi_miso_i[2]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_1 input50 (.A(sport_i[49]),
    .X(net50));
 sky130_fd_sc_hd__buf_1 input51 (.A(sport_i[4]),
    .X(net51));
 sky130_fd_sc_hd__buf_1 input52 (.A(sport_i[50]),
    .X(net52));
 sky130_fd_sc_hd__buf_1 input53 (.A(sport_i[51]),
    .X(net53));
 sky130_fd_sc_hd__clkbuf_2 input54 (.A(sport_i[52]),
    .X(net54));
 sky130_fd_sc_hd__clkbuf_4 input55 (.A(sport_i[54]),
    .X(net55));
 sky130_fd_sc_hd__clkbuf_4 input56 (.A(sport_i[55]),
    .X(net56));
 sky130_fd_sc_hd__buf_2 input57 (.A(sport_i[56]),
    .X(net57));
 sky130_fd_sc_hd__clkbuf_1 input58 (.A(sport_i[5]),
    .X(net58));
 sky130_fd_sc_hd__clkbuf_1 input59 (.A(sport_i[6]),
    .X(net59));
 sky130_fd_sc_hd__buf_2 input6 (.A(spi_miso_i[3]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_1 input60 (.A(sport_i[7]),
    .X(net60));
 sky130_fd_sc_hd__buf_1 input61 (.A(sport_i[8]),
    .X(net61));
 sky130_fd_sc_hd__buf_1 input62 (.A(sport_i[9]),
    .X(net62));
 sky130_fd_sc_hd__buf_1 input7 (.A(sport_i[0]),
    .X(net7));
 sky130_fd_sc_hd__buf_1 input8 (.A(sport_i[10]),
    .X(net8));
 sky130_fd_sc_hd__buf_1 input9 (.A(sport_i[11]),
    .X(net9));
 sky130_fd_sc_hd__buf_12 output100 (.A(net100),
    .X(sport_o[7]));
 sky130_fd_sc_hd__buf_12 output101 (.A(net101),
    .X(sport_o[8]));
 sky130_fd_sc_hd__buf_12 output102 (.A(net102),
    .X(sport_o[9]));
 sky130_fd_sc_hd__buf_12 output63 (.A(net63),
    .X(spi_clk_o));
 sky130_fd_sc_hd__buf_12 output64 (.A(net64),
    .X(spi_cs_o));
 sky130_fd_sc_hd__buf_12 output65 (.A(net65),
    .X(spi_mosi_o[0]));
 sky130_fd_sc_hd__buf_12 output66 (.A(net66),
    .X(spi_mosi_o[1]));
 sky130_fd_sc_hd__buf_12 output67 (.A(net67),
    .X(spi_mosi_o[2]));
 sky130_fd_sc_hd__buf_12 output68 (.A(net68),
    .X(spi_mosi_o[3]));
 sky130_fd_sc_hd__buf_12 output69 (.A(net69),
    .X(sport_o[0]));
 sky130_fd_sc_hd__buf_12 output70 (.A(net70),
    .X(sport_o[10]));
 sky130_fd_sc_hd__buf_12 output71 (.A(net71),
    .X(sport_o[11]));
 sky130_fd_sc_hd__buf_12 output72 (.A(net72),
    .X(sport_o[12]));
 sky130_fd_sc_hd__buf_12 output73 (.A(net73),
    .X(sport_o[13]));
 sky130_fd_sc_hd__buf_12 output74 (.A(net74),
    .X(sport_o[14]));
 sky130_fd_sc_hd__buf_12 output75 (.A(net75),
    .X(sport_o[15]));
 sky130_fd_sc_hd__buf_12 output76 (.A(net76),
    .X(sport_o[16]));
 sky130_fd_sc_hd__buf_12 output77 (.A(net77),
    .X(sport_o[17]));
 sky130_fd_sc_hd__buf_12 output78 (.A(net78),
    .X(sport_o[18]));
 sky130_fd_sc_hd__buf_12 output79 (.A(net79),
    .X(sport_o[19]));
 sky130_fd_sc_hd__buf_12 output80 (.A(net80),
    .X(sport_o[1]));
 sky130_fd_sc_hd__buf_12 output81 (.A(net81),
    .X(sport_o[20]));
 sky130_fd_sc_hd__buf_12 output82 (.A(net82),
    .X(sport_o[21]));
 sky130_fd_sc_hd__buf_12 output83 (.A(net83),
    .X(sport_o[22]));
 sky130_fd_sc_hd__buf_12 output84 (.A(net84),
    .X(sport_o[23]));
 sky130_fd_sc_hd__buf_12 output85 (.A(net85),
    .X(sport_o[24]));
 sky130_fd_sc_hd__buf_12 output86 (.A(net86),
    .X(sport_o[25]));
 sky130_fd_sc_hd__buf_12 output87 (.A(net87),
    .X(sport_o[26]));
 sky130_fd_sc_hd__buf_12 output88 (.A(net88),
    .X(sport_o[27]));
 sky130_fd_sc_hd__buf_12 output89 (.A(net89),
    .X(sport_o[28]));
 sky130_fd_sc_hd__buf_12 output90 (.A(net90),
    .X(sport_o[29]));
 sky130_fd_sc_hd__buf_12 output91 (.A(net91),
    .X(sport_o[2]));
 sky130_fd_sc_hd__buf_12 output92 (.A(net92),
    .X(sport_o[30]));
 sky130_fd_sc_hd__buf_12 output93 (.A(net93),
    .X(sport_o[31]));
 sky130_fd_sc_hd__buf_12 output94 (.A(net94),
    .X(sport_o[32]));
 sky130_fd_sc_hd__buf_12 output95 (.A(net95),
    .X(sport_o[33]));
 sky130_fd_sc_hd__buf_12 output96 (.A(net96),
    .X(sport_o[3]));
 sky130_fd_sc_hd__buf_12 output97 (.A(net97),
    .X(sport_o[4]));
 sky130_fd_sc_hd__buf_12 output98 (.A(net98),
    .X(sport_o[5]));
 sky130_fd_sc_hd__buf_12 output99 (.A(net99),
    .X(sport_o[6]));
 sky130_fd_sc_hd__conb_1 spi_mem_m_108 (.LO(net108));
 assign spi_dqsm_o = net108;
endmodule

