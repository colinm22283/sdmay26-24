VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO spi_mem_m
  CLASS BLOCK ;
  FOREIGN spi_mem_m ;
  ORIGIN 0.000 0.000 ;
  SIZE 300.000 BY 300.000 ;
  PIN clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met2 ;
        RECT 74.610 296.000 74.890 300.000 ;
    END
  END clk_i
  PIN nrst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met2 ;
        RECT 224.570 296.000 224.850 300.000 ;
    END
  END nrst_i
  PIN spi_clk_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 12.970 0.000 13.250 4.000 ;
    END
  END spi_clk_o
  PIN spi_cs_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 37.810 0.000 38.090 4.000 ;
    END
  END spi_cs_o
  PIN spi_dqsm_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 62.650 0.000 62.930 4.000 ;
    END
  END spi_dqsm_i
  PIN spi_dqsm_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.490 0.000 87.770 4.000 ;
    END
  END spi_dqsm_o
  PIN spi_miso_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 112.330 0.000 112.610 4.000 ;
    END
  END spi_miso_i[0]
  PIN spi_miso_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 162.010 0.000 162.290 4.000 ;
    END
  END spi_miso_i[1]
  PIN spi_miso_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 211.690 0.000 211.970 4.000 ;
    END
  END spi_miso_i[2]
  PIN spi_miso_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 261.370 0.000 261.650 4.000 ;
    END
  END spi_miso_i[3]
  PIN spi_mosi_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 137.170 0.000 137.450 4.000 ;
    END
  END spi_mosi_o[0]
  PIN spi_mosi_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 186.850 0.000 187.130 4.000 ;
    END
  END spi_mosi_o[1]
  PIN spi_mosi_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 236.530 0.000 236.810 4.000 ;
    END
  END spi_mosi_o[2]
  PIN spi_mosi_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 286.210 0.000 286.490 4.000 ;
    END
  END spi_mosi_o[3]
  PIN sport_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 35.400 300.000 36.000 ;
    END
  END sport_i[0]
  PIN sport_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 76.200 300.000 76.800 ;
    END
  END sport_i[10]
  PIN sport_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 80.280 300.000 80.880 ;
    END
  END sport_i[11]
  PIN sport_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 84.360 300.000 84.960 ;
    END
  END sport_i[12]
  PIN sport_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 88.440 300.000 89.040 ;
    END
  END sport_i[13]
  PIN sport_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 92.520 300.000 93.120 ;
    END
  END sport_i[14]
  PIN sport_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 96.600 300.000 97.200 ;
    END
  END sport_i[15]
  PIN sport_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 100.680 300.000 101.280 ;
    END
  END sport_i[16]
  PIN sport_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 104.760 300.000 105.360 ;
    END
  END sport_i[17]
  PIN sport_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 108.840 300.000 109.440 ;
    END
  END sport_i[18]
  PIN sport_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 112.920 300.000 113.520 ;
    END
  END sport_i[19]
  PIN sport_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 39.480 300.000 40.080 ;
    END
  END sport_i[1]
  PIN sport_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 117.000 300.000 117.600 ;
    END
  END sport_i[20]
  PIN sport_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 121.080 300.000 121.680 ;
    END
  END sport_i[21]
  PIN sport_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 125.160 300.000 125.760 ;
    END
  END sport_i[22]
  PIN sport_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 129.240 300.000 129.840 ;
    END
  END sport_i[23]
  PIN sport_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 133.320 300.000 133.920 ;
    END
  END sport_i[24]
  PIN sport_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 137.400 300.000 138.000 ;
    END
  END sport_i[25]
  PIN sport_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 141.480 300.000 142.080 ;
    END
  END sport_i[26]
  PIN sport_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 145.560 300.000 146.160 ;
    END
  END sport_i[27]
  PIN sport_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 149.640 300.000 150.240 ;
    END
  END sport_i[28]
  PIN sport_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 153.720 300.000 154.320 ;
    END
  END sport_i[29]
  PIN sport_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 43.560 300.000 44.160 ;
    END
  END sport_i[2]
  PIN sport_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 157.800 300.000 158.400 ;
    END
  END sport_i[30]
  PIN sport_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 161.880 300.000 162.480 ;
    END
  END sport_i[31]
  PIN sport_i[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 165.960 300.000 166.560 ;
    END
  END sport_i[32]
  PIN sport_i[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 170.040 300.000 170.640 ;
    END
  END sport_i[33]
  PIN sport_i[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 174.120 300.000 174.720 ;
    END
  END sport_i[34]
  PIN sport_i[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 178.200 300.000 178.800 ;
    END
  END sport_i[35]
  PIN sport_i[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 182.280 300.000 182.880 ;
    END
  END sport_i[36]
  PIN sport_i[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 186.360 300.000 186.960 ;
    END
  END sport_i[37]
  PIN sport_i[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 190.440 300.000 191.040 ;
    END
  END sport_i[38]
  PIN sport_i[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 194.520 300.000 195.120 ;
    END
  END sport_i[39]
  PIN sport_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 47.640 300.000 48.240 ;
    END
  END sport_i[3]
  PIN sport_i[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 198.600 300.000 199.200 ;
    END
  END sport_i[40]
  PIN sport_i[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 202.680 300.000 203.280 ;
    END
  END sport_i[41]
  PIN sport_i[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 206.760 300.000 207.360 ;
    END
  END sport_i[42]
  PIN sport_i[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 210.840 300.000 211.440 ;
    END
  END sport_i[43]
  PIN sport_i[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 214.920 300.000 215.520 ;
    END
  END sport_i[44]
  PIN sport_i[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 219.000 300.000 219.600 ;
    END
  END sport_i[45]
  PIN sport_i[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 223.080 300.000 223.680 ;
    END
  END sport_i[46]
  PIN sport_i[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 227.160 300.000 227.760 ;
    END
  END sport_i[47]
  PIN sport_i[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 231.240 300.000 231.840 ;
    END
  END sport_i[48]
  PIN sport_i[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 235.320 300.000 235.920 ;
    END
  END sport_i[49]
  PIN sport_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 51.720 300.000 52.320 ;
    END
  END sport_i[4]
  PIN sport_i[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 239.400 300.000 240.000 ;
    END
  END sport_i[50]
  PIN sport_i[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 243.480 300.000 244.080 ;
    END
  END sport_i[51]
  PIN sport_i[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 296.000 247.560 300.000 248.160 ;
    END
  END sport_i[52]
  PIN sport_i[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 251.640 300.000 252.240 ;
    END
  END sport_i[53]
  PIN sport_i[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 296.000 255.720 300.000 256.320 ;
    END
  END sport_i[54]
  PIN sport_i[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 296.000 259.800 300.000 260.400 ;
    END
  END sport_i[55]
  PIN sport_i[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 296.000 263.880 300.000 264.480 ;
    END
  END sport_i[56]
  PIN sport_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 55.800 300.000 56.400 ;
    END
  END sport_i[5]
  PIN sport_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 59.880 300.000 60.480 ;
    END
  END sport_i[6]
  PIN sport_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 63.960 300.000 64.560 ;
    END
  END sport_i[7]
  PIN sport_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 68.040 300.000 68.640 ;
    END
  END sport_i[8]
  PIN sport_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 296.000 72.120 300.000 72.720 ;
    END
  END sport_i[9]
  PIN sport_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 15.000 4.000 15.600 ;
    END
  END sport_o[0]
  PIN sport_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 96.600 4.000 97.200 ;
    END
  END sport_o[10]
  PIN sport_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 104.760 4.000 105.360 ;
    END
  END sport_o[11]
  PIN sport_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 112.920 4.000 113.520 ;
    END
  END sport_o[12]
  PIN sport_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 121.080 4.000 121.680 ;
    END
  END sport_o[13]
  PIN sport_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 129.240 4.000 129.840 ;
    END
  END sport_o[14]
  PIN sport_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 137.400 4.000 138.000 ;
    END
  END sport_o[15]
  PIN sport_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 145.560 4.000 146.160 ;
    END
  END sport_o[16]
  PIN sport_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 153.720 4.000 154.320 ;
    END
  END sport_o[17]
  PIN sport_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 161.880 4.000 162.480 ;
    END
  END sport_o[18]
  PIN sport_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 170.040 4.000 170.640 ;
    END
  END sport_o[19]
  PIN sport_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 23.160 4.000 23.760 ;
    END
  END sport_o[1]
  PIN sport_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 178.200 4.000 178.800 ;
    END
  END sport_o[20]
  PIN sport_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 186.360 4.000 186.960 ;
    END
  END sport_o[21]
  PIN sport_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 194.520 4.000 195.120 ;
    END
  END sport_o[22]
  PIN sport_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 202.680 4.000 203.280 ;
    END
  END sport_o[23]
  PIN sport_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 210.840 4.000 211.440 ;
    END
  END sport_o[24]
  PIN sport_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 219.000 4.000 219.600 ;
    END
  END sport_o[25]
  PIN sport_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 227.160 4.000 227.760 ;
    END
  END sport_o[26]
  PIN sport_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 235.320 4.000 235.920 ;
    END
  END sport_o[27]
  PIN sport_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 243.480 4.000 244.080 ;
    END
  END sport_o[28]
  PIN sport_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 251.640 4.000 252.240 ;
    END
  END sport_o[29]
  PIN sport_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 31.320 4.000 31.920 ;
    END
  END sport_o[2]
  PIN sport_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 259.800 4.000 260.400 ;
    END
  END sport_o[30]
  PIN sport_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 267.960 4.000 268.560 ;
    END
  END sport_o[31]
  PIN sport_o[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 276.120 4.000 276.720 ;
    END
  END sport_o[32]
  PIN sport_o[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 284.280 4.000 284.880 ;
    END
  END sport_o[33]
  PIN sport_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 39.480 4.000 40.080 ;
    END
  END sport_o[3]
  PIN sport_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 47.640 4.000 48.240 ;
    END
  END sport_o[4]
  PIN sport_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 55.800 4.000 56.400 ;
    END
  END sport_o[5]
  PIN sport_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 63.960 4.000 64.560 ;
    END
  END sport_o[6]
  PIN sport_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 72.120 4.000 72.720 ;
    END
  END sport_o[7]
  PIN sport_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 80.280 4.000 80.880 ;
    END
  END sport_o[8]
  PIN sport_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 88.440 4.000 89.040 ;
    END
  END sport_o[9]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 288.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 288.560 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 288.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 288.560 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 294.400 288.405 ;
      LAYER met1 ;
        RECT 4.670 9.900 296.170 288.560 ;
      LAYER met2 ;
        RECT 4.690 295.720 74.330 296.000 ;
        RECT 75.170 295.720 224.290 296.000 ;
        RECT 225.130 295.720 296.140 296.000 ;
        RECT 4.690 4.280 296.140 295.720 ;
        RECT 4.690 3.670 12.690 4.280 ;
        RECT 13.530 3.670 37.530 4.280 ;
        RECT 38.370 3.670 62.370 4.280 ;
        RECT 63.210 3.670 87.210 4.280 ;
        RECT 88.050 3.670 112.050 4.280 ;
        RECT 112.890 3.670 136.890 4.280 ;
        RECT 137.730 3.670 161.730 4.280 ;
        RECT 162.570 3.670 186.570 4.280 ;
        RECT 187.410 3.670 211.410 4.280 ;
        RECT 212.250 3.670 236.250 4.280 ;
        RECT 237.090 3.670 261.090 4.280 ;
        RECT 261.930 3.670 285.930 4.280 ;
        RECT 286.770 3.670 296.140 4.280 ;
      LAYER met3 ;
        RECT 3.990 285.280 296.000 288.485 ;
        RECT 4.400 283.880 296.000 285.280 ;
        RECT 3.990 277.120 296.000 283.880 ;
        RECT 4.400 275.720 296.000 277.120 ;
        RECT 3.990 268.960 296.000 275.720 ;
        RECT 4.400 267.560 296.000 268.960 ;
        RECT 3.990 264.880 296.000 267.560 ;
        RECT 3.990 263.480 295.600 264.880 ;
        RECT 3.990 260.800 296.000 263.480 ;
        RECT 4.400 259.400 295.600 260.800 ;
        RECT 3.990 256.720 296.000 259.400 ;
        RECT 3.990 255.320 295.600 256.720 ;
        RECT 3.990 252.640 296.000 255.320 ;
        RECT 4.400 251.240 295.600 252.640 ;
        RECT 3.990 248.560 296.000 251.240 ;
        RECT 3.990 247.160 295.600 248.560 ;
        RECT 3.990 244.480 296.000 247.160 ;
        RECT 4.400 243.080 295.600 244.480 ;
        RECT 3.990 240.400 296.000 243.080 ;
        RECT 3.990 239.000 295.600 240.400 ;
        RECT 3.990 236.320 296.000 239.000 ;
        RECT 4.400 234.920 295.600 236.320 ;
        RECT 3.990 232.240 296.000 234.920 ;
        RECT 3.990 230.840 295.600 232.240 ;
        RECT 3.990 228.160 296.000 230.840 ;
        RECT 4.400 226.760 295.600 228.160 ;
        RECT 3.990 224.080 296.000 226.760 ;
        RECT 3.990 222.680 295.600 224.080 ;
        RECT 3.990 220.000 296.000 222.680 ;
        RECT 4.400 218.600 295.600 220.000 ;
        RECT 3.990 215.920 296.000 218.600 ;
        RECT 3.990 214.520 295.600 215.920 ;
        RECT 3.990 211.840 296.000 214.520 ;
        RECT 4.400 210.440 295.600 211.840 ;
        RECT 3.990 207.760 296.000 210.440 ;
        RECT 3.990 206.360 295.600 207.760 ;
        RECT 3.990 203.680 296.000 206.360 ;
        RECT 4.400 202.280 295.600 203.680 ;
        RECT 3.990 199.600 296.000 202.280 ;
        RECT 3.990 198.200 295.600 199.600 ;
        RECT 3.990 195.520 296.000 198.200 ;
        RECT 4.400 194.120 295.600 195.520 ;
        RECT 3.990 191.440 296.000 194.120 ;
        RECT 3.990 190.040 295.600 191.440 ;
        RECT 3.990 187.360 296.000 190.040 ;
        RECT 4.400 185.960 295.600 187.360 ;
        RECT 3.990 183.280 296.000 185.960 ;
        RECT 3.990 181.880 295.600 183.280 ;
        RECT 3.990 179.200 296.000 181.880 ;
        RECT 4.400 177.800 295.600 179.200 ;
        RECT 3.990 175.120 296.000 177.800 ;
        RECT 3.990 173.720 295.600 175.120 ;
        RECT 3.990 171.040 296.000 173.720 ;
        RECT 4.400 169.640 295.600 171.040 ;
        RECT 3.990 166.960 296.000 169.640 ;
        RECT 3.990 165.560 295.600 166.960 ;
        RECT 3.990 162.880 296.000 165.560 ;
        RECT 4.400 161.480 295.600 162.880 ;
        RECT 3.990 158.800 296.000 161.480 ;
        RECT 3.990 157.400 295.600 158.800 ;
        RECT 3.990 154.720 296.000 157.400 ;
        RECT 4.400 153.320 295.600 154.720 ;
        RECT 3.990 150.640 296.000 153.320 ;
        RECT 3.990 149.240 295.600 150.640 ;
        RECT 3.990 146.560 296.000 149.240 ;
        RECT 4.400 145.160 295.600 146.560 ;
        RECT 3.990 142.480 296.000 145.160 ;
        RECT 3.990 141.080 295.600 142.480 ;
        RECT 3.990 138.400 296.000 141.080 ;
        RECT 4.400 137.000 295.600 138.400 ;
        RECT 3.990 134.320 296.000 137.000 ;
        RECT 3.990 132.920 295.600 134.320 ;
        RECT 3.990 130.240 296.000 132.920 ;
        RECT 4.400 128.840 295.600 130.240 ;
        RECT 3.990 126.160 296.000 128.840 ;
        RECT 3.990 124.760 295.600 126.160 ;
        RECT 3.990 122.080 296.000 124.760 ;
        RECT 4.400 120.680 295.600 122.080 ;
        RECT 3.990 118.000 296.000 120.680 ;
        RECT 3.990 116.600 295.600 118.000 ;
        RECT 3.990 113.920 296.000 116.600 ;
        RECT 4.400 112.520 295.600 113.920 ;
        RECT 3.990 109.840 296.000 112.520 ;
        RECT 3.990 108.440 295.600 109.840 ;
        RECT 3.990 105.760 296.000 108.440 ;
        RECT 4.400 104.360 295.600 105.760 ;
        RECT 3.990 101.680 296.000 104.360 ;
        RECT 3.990 100.280 295.600 101.680 ;
        RECT 3.990 97.600 296.000 100.280 ;
        RECT 4.400 96.200 295.600 97.600 ;
        RECT 3.990 93.520 296.000 96.200 ;
        RECT 3.990 92.120 295.600 93.520 ;
        RECT 3.990 89.440 296.000 92.120 ;
        RECT 4.400 88.040 295.600 89.440 ;
        RECT 3.990 85.360 296.000 88.040 ;
        RECT 3.990 83.960 295.600 85.360 ;
        RECT 3.990 81.280 296.000 83.960 ;
        RECT 4.400 79.880 295.600 81.280 ;
        RECT 3.990 77.200 296.000 79.880 ;
        RECT 3.990 75.800 295.600 77.200 ;
        RECT 3.990 73.120 296.000 75.800 ;
        RECT 4.400 71.720 295.600 73.120 ;
        RECT 3.990 69.040 296.000 71.720 ;
        RECT 3.990 67.640 295.600 69.040 ;
        RECT 3.990 64.960 296.000 67.640 ;
        RECT 4.400 63.560 295.600 64.960 ;
        RECT 3.990 60.880 296.000 63.560 ;
        RECT 3.990 59.480 295.600 60.880 ;
        RECT 3.990 56.800 296.000 59.480 ;
        RECT 4.400 55.400 295.600 56.800 ;
        RECT 3.990 52.720 296.000 55.400 ;
        RECT 3.990 51.320 295.600 52.720 ;
        RECT 3.990 48.640 296.000 51.320 ;
        RECT 4.400 47.240 295.600 48.640 ;
        RECT 3.990 44.560 296.000 47.240 ;
        RECT 3.990 43.160 295.600 44.560 ;
        RECT 3.990 40.480 296.000 43.160 ;
        RECT 4.400 39.080 295.600 40.480 ;
        RECT 3.990 36.400 296.000 39.080 ;
        RECT 3.990 35.000 295.600 36.400 ;
        RECT 3.990 32.320 296.000 35.000 ;
        RECT 4.400 30.920 296.000 32.320 ;
        RECT 3.990 24.160 296.000 30.920 ;
        RECT 4.400 22.760 296.000 24.160 ;
        RECT 3.990 16.000 296.000 22.760 ;
        RECT 4.400 14.600 296.000 16.000 ;
        RECT 3.990 10.715 296.000 14.600 ;
      LAYER met4 ;
        RECT 248.695 91.975 251.040 146.025 ;
        RECT 253.440 91.975 256.385 146.025 ;
  END
END spi_mem_m
END LIBRARY

