// This is the unpowered netlist.
module wavg_pipe_m (clk_i,
    mstream_i,
    nrst_i,
    sstream_o,
    mstream_o,
    sstream_i,
    t0x,
    t0y,
    t1x,
    t1y,
    t2x,
    t2y,
    v0z,
    v1z,
    v2z);
 input clk_i;
 input mstream_i;
 input nrst_i;
 output sstream_o;
 output [115:0] mstream_o;
 input [115:0] sstream_i;
 input [31:0] t0x;
 input [31:0] t0y;
 input [31:0] t1x;
 input [31:0] t1y;
 input [31:0] t2x;
 input [31:0] t2y;
 input [31:0] v0z;
 input [31:0] v1z;
 input [31:0] v2z;

 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire _05356_;
 wire _05357_;
 wire _05358_;
 wire _05359_;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire _05373_;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05377_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire _05383_;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire _05387_;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire _05411_;
 wire _05412_;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire _05420_;
 wire _05421_;
 wire _05422_;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire _05429_;
 wire _05430_;
 wire _05431_;
 wire _05432_;
 wire _05433_;
 wire _05434_;
 wire _05435_;
 wire _05436_;
 wire _05437_;
 wire _05438_;
 wire _05439_;
 wire _05440_;
 wire _05441_;
 wire _05442_;
 wire _05443_;
 wire _05444_;
 wire _05445_;
 wire _05446_;
 wire _05447_;
 wire _05448_;
 wire _05449_;
 wire _05450_;
 wire _05451_;
 wire _05452_;
 wire _05453_;
 wire _05454_;
 wire _05455_;
 wire _05456_;
 wire _05457_;
 wire _05458_;
 wire _05459_;
 wire _05460_;
 wire _05461_;
 wire _05462_;
 wire _05463_;
 wire _05464_;
 wire _05465_;
 wire _05466_;
 wire _05467_;
 wire _05468_;
 wire _05469_;
 wire _05470_;
 wire _05471_;
 wire _05472_;
 wire _05473_;
 wire _05474_;
 wire _05475_;
 wire _05476_;
 wire _05477_;
 wire _05478_;
 wire _05479_;
 wire _05480_;
 wire _05481_;
 wire _05482_;
 wire _05483_;
 wire _05484_;
 wire _05485_;
 wire _05486_;
 wire _05487_;
 wire _05488_;
 wire _05489_;
 wire _05490_;
 wire _05491_;
 wire _05492_;
 wire _05493_;
 wire _05494_;
 wire _05495_;
 wire _05496_;
 wire _05497_;
 wire _05498_;
 wire _05499_;
 wire _05500_;
 wire _05501_;
 wire _05502_;
 wire _05503_;
 wire _05504_;
 wire _05505_;
 wire _05506_;
 wire _05507_;
 wire _05508_;
 wire _05509_;
 wire _05510_;
 wire _05511_;
 wire _05512_;
 wire _05513_;
 wire _05514_;
 wire _05515_;
 wire _05516_;
 wire _05517_;
 wire _05518_;
 wire _05519_;
 wire _05520_;
 wire _05521_;
 wire _05522_;
 wire _05523_;
 wire _05524_;
 wire _05525_;
 wire _05526_;
 wire _05527_;
 wire _05528_;
 wire _05529_;
 wire _05530_;
 wire _05531_;
 wire _05532_;
 wire _05533_;
 wire _05534_;
 wire _05535_;
 wire _05536_;
 wire _05537_;
 wire _05538_;
 wire _05539_;
 wire _05540_;
 wire _05541_;
 wire _05542_;
 wire _05543_;
 wire _05544_;
 wire _05545_;
 wire _05546_;
 wire _05547_;
 wire _05548_;
 wire _05549_;
 wire _05550_;
 wire _05551_;
 wire _05552_;
 wire _05553_;
 wire _05554_;
 wire _05555_;
 wire _05556_;
 wire _05557_;
 wire _05558_;
 wire _05559_;
 wire _05560_;
 wire _05561_;
 wire _05562_;
 wire _05563_;
 wire _05564_;
 wire _05565_;
 wire _05566_;
 wire _05567_;
 wire _05568_;
 wire _05569_;
 wire _05570_;
 wire _05571_;
 wire _05572_;
 wire _05573_;
 wire _05574_;
 wire _05575_;
 wire _05576_;
 wire _05577_;
 wire _05578_;
 wire _05579_;
 wire _05580_;
 wire _05581_;
 wire _05582_;
 wire _05583_;
 wire _05584_;
 wire _05585_;
 wire _05586_;
 wire _05587_;
 wire _05588_;
 wire _05589_;
 wire _05590_;
 wire _05591_;
 wire _05592_;
 wire _05593_;
 wire _05594_;
 wire _05595_;
 wire _05596_;
 wire _05597_;
 wire _05598_;
 wire _05599_;
 wire _05600_;
 wire _05601_;
 wire _05602_;
 wire _05603_;
 wire _05604_;
 wire _05605_;
 wire _05606_;
 wire _05607_;
 wire _05608_;
 wire _05609_;
 wire _05610_;
 wire _05611_;
 wire _05612_;
 wire _05613_;
 wire _05614_;
 wire _05615_;
 wire _05616_;
 wire _05617_;
 wire _05618_;
 wire _05619_;
 wire _05620_;
 wire _05621_;
 wire _05622_;
 wire _05623_;
 wire _05624_;
 wire _05625_;
 wire _05626_;
 wire _05627_;
 wire _05628_;
 wire _05629_;
 wire _05630_;
 wire _05631_;
 wire _05632_;
 wire _05633_;
 wire _05634_;
 wire _05635_;
 wire _05636_;
 wire _05637_;
 wire _05638_;
 wire _05639_;
 wire _05640_;
 wire _05641_;
 wire _05642_;
 wire _05643_;
 wire _05644_;
 wire _05645_;
 wire _05646_;
 wire _05647_;
 wire _05648_;
 wire _05649_;
 wire _05650_;
 wire _05651_;
 wire _05652_;
 wire _05653_;
 wire _05654_;
 wire _05655_;
 wire _05656_;
 wire _05657_;
 wire _05658_;
 wire _05659_;
 wire _05660_;
 wire _05661_;
 wire _05662_;
 wire _05663_;
 wire _05664_;
 wire _05665_;
 wire _05666_;
 wire _05667_;
 wire _05668_;
 wire _05669_;
 wire _05670_;
 wire _05671_;
 wire _05672_;
 wire _05673_;
 wire _05674_;
 wire _05675_;
 wire _05676_;
 wire _05677_;
 wire _05678_;
 wire _05679_;
 wire _05680_;
 wire _05681_;
 wire _05682_;
 wire _05683_;
 wire _05684_;
 wire _05685_;
 wire _05686_;
 wire _05687_;
 wire _05688_;
 wire _05689_;
 wire _05690_;
 wire _05691_;
 wire _05692_;
 wire _05693_;
 wire _05694_;
 wire _05695_;
 wire _05696_;
 wire _05697_;
 wire _05698_;
 wire _05699_;
 wire _05700_;
 wire _05701_;
 wire _05702_;
 wire _05703_;
 wire _05704_;
 wire _05705_;
 wire _05706_;
 wire _05707_;
 wire _05708_;
 wire _05709_;
 wire _05710_;
 wire _05711_;
 wire _05712_;
 wire _05713_;
 wire _05714_;
 wire _05715_;
 wire _05716_;
 wire _05717_;
 wire _05718_;
 wire _05719_;
 wire _05720_;
 wire _05721_;
 wire _05722_;
 wire _05723_;
 wire _05724_;
 wire _05725_;
 wire _05726_;
 wire _05727_;
 wire _05728_;
 wire _05729_;
 wire _05730_;
 wire _05731_;
 wire _05732_;
 wire _05733_;
 wire _05734_;
 wire _05735_;
 wire _05736_;
 wire _05737_;
 wire _05738_;
 wire _05739_;
 wire _05740_;
 wire _05741_;
 wire _05742_;
 wire _05743_;
 wire _05744_;
 wire _05745_;
 wire _05746_;
 wire _05747_;
 wire _05748_;
 wire _05749_;
 wire _05750_;
 wire _05751_;
 wire _05752_;
 wire _05753_;
 wire _05754_;
 wire _05755_;
 wire _05756_;
 wire _05757_;
 wire _05758_;
 wire _05759_;
 wire _05760_;
 wire _05761_;
 wire _05762_;
 wire _05763_;
 wire _05764_;
 wire _05765_;
 wire _05766_;
 wire _05767_;
 wire _05768_;
 wire _05769_;
 wire _05770_;
 wire _05771_;
 wire _05772_;
 wire _05773_;
 wire _05774_;
 wire _05775_;
 wire _05776_;
 wire _05777_;
 wire _05778_;
 wire _05779_;
 wire _05780_;
 wire _05781_;
 wire _05782_;
 wire _05783_;
 wire _05784_;
 wire _05785_;
 wire _05786_;
 wire _05787_;
 wire _05788_;
 wire _05789_;
 wire _05790_;
 wire _05791_;
 wire _05792_;
 wire _05793_;
 wire _05794_;
 wire _05795_;
 wire _05796_;
 wire _05797_;
 wire _05798_;
 wire _05799_;
 wire _05800_;
 wire _05801_;
 wire _05802_;
 wire _05803_;
 wire _05804_;
 wire _05805_;
 wire _05806_;
 wire _05807_;
 wire _05808_;
 wire _05809_;
 wire _05810_;
 wire _05811_;
 wire _05812_;
 wire _05813_;
 wire _05814_;
 wire _05815_;
 wire _05816_;
 wire _05817_;
 wire _05818_;
 wire _05819_;
 wire _05820_;
 wire _05821_;
 wire _05822_;
 wire _05823_;
 wire _05824_;
 wire _05825_;
 wire _05826_;
 wire _05827_;
 wire _05828_;
 wire _05829_;
 wire _05830_;
 wire _05831_;
 wire _05832_;
 wire _05833_;
 wire _05834_;
 wire _05835_;
 wire _05836_;
 wire _05837_;
 wire _05838_;
 wire _05839_;
 wire _05840_;
 wire _05841_;
 wire _05842_;
 wire _05843_;
 wire _05844_;
 wire _05845_;
 wire _05846_;
 wire _05847_;
 wire _05848_;
 wire _05849_;
 wire _05850_;
 wire _05851_;
 wire _05852_;
 wire _05853_;
 wire _05854_;
 wire _05855_;
 wire _05856_;
 wire _05857_;
 wire _05858_;
 wire _05859_;
 wire _05860_;
 wire _05861_;
 wire _05862_;
 wire _05863_;
 wire _05864_;
 wire _05865_;
 wire _05866_;
 wire _05867_;
 wire _05868_;
 wire _05869_;
 wire _05870_;
 wire _05871_;
 wire _05872_;
 wire _05873_;
 wire _05874_;
 wire _05875_;
 wire _05876_;
 wire _05877_;
 wire _05878_;
 wire _05879_;
 wire _05880_;
 wire _05881_;
 wire _05882_;
 wire _05883_;
 wire _05884_;
 wire _05885_;
 wire _05886_;
 wire _05887_;
 wire _05888_;
 wire _05889_;
 wire _05890_;
 wire _05891_;
 wire _05892_;
 wire _05893_;
 wire _05894_;
 wire _05895_;
 wire _05896_;
 wire _05897_;
 wire _05898_;
 wire _05899_;
 wire _05900_;
 wire _05901_;
 wire _05902_;
 wire _05903_;
 wire _05904_;
 wire _05905_;
 wire _05906_;
 wire _05907_;
 wire _05908_;
 wire _05909_;
 wire _05910_;
 wire _05911_;
 wire _05912_;
 wire _05913_;
 wire _05914_;
 wire _05915_;
 wire _05916_;
 wire _05917_;
 wire _05918_;
 wire _05919_;
 wire _05920_;
 wire _05921_;
 wire _05922_;
 wire _05923_;
 wire _05924_;
 wire _05925_;
 wire _05926_;
 wire _05927_;
 wire _05928_;
 wire _05929_;
 wire _05930_;
 wire _05931_;
 wire _05932_;
 wire _05933_;
 wire _05934_;
 wire _05935_;
 wire _05936_;
 wire _05937_;
 wire _05938_;
 wire _05939_;
 wire _05940_;
 wire _05941_;
 wire _05942_;
 wire _05943_;
 wire _05944_;
 wire _05945_;
 wire _05946_;
 wire _05947_;
 wire _05948_;
 wire _05949_;
 wire _05950_;
 wire _05951_;
 wire _05952_;
 wire _05953_;
 wire _05954_;
 wire _05955_;
 wire _05956_;
 wire _05957_;
 wire _05958_;
 wire _05959_;
 wire _05960_;
 wire _05961_;
 wire _05962_;
 wire _05963_;
 wire _05964_;
 wire _05965_;
 wire _05966_;
 wire _05967_;
 wire _05968_;
 wire _05969_;
 wire _05970_;
 wire _05971_;
 wire _05972_;
 wire _05973_;
 wire _05974_;
 wire _05975_;
 wire _05976_;
 wire _05977_;
 wire _05978_;
 wire _05979_;
 wire _05980_;
 wire _05981_;
 wire _05982_;
 wire _05983_;
 wire _05984_;
 wire _05985_;
 wire _05986_;
 wire _05987_;
 wire _05988_;
 wire _05989_;
 wire _05990_;
 wire _05991_;
 wire _05992_;
 wire _05993_;
 wire _05994_;
 wire _05995_;
 wire _05996_;
 wire _05997_;
 wire _05998_;
 wire _05999_;
 wire _06000_;
 wire _06001_;
 wire _06002_;
 wire _06003_;
 wire _06004_;
 wire _06005_;
 wire _06006_;
 wire _06007_;
 wire _06008_;
 wire _06009_;
 wire _06010_;
 wire _06011_;
 wire _06012_;
 wire _06013_;
 wire _06014_;
 wire _06015_;
 wire _06016_;
 wire _06017_;
 wire _06018_;
 wire _06019_;
 wire _06020_;
 wire _06021_;
 wire _06022_;
 wire _06023_;
 wire _06024_;
 wire _06025_;
 wire _06026_;
 wire _06027_;
 wire _06028_;
 wire _06029_;
 wire _06030_;
 wire _06031_;
 wire _06032_;
 wire _06033_;
 wire _06034_;
 wire _06035_;
 wire _06036_;
 wire _06037_;
 wire _06038_;
 wire _06039_;
 wire _06040_;
 wire _06041_;
 wire _06042_;
 wire _06043_;
 wire _06044_;
 wire _06045_;
 wire _06046_;
 wire _06047_;
 wire _06048_;
 wire _06049_;
 wire _06050_;
 wire _06051_;
 wire _06052_;
 wire _06053_;
 wire _06054_;
 wire _06055_;
 wire _06056_;
 wire _06057_;
 wire _06058_;
 wire _06059_;
 wire _06060_;
 wire _06061_;
 wire _06062_;
 wire _06063_;
 wire _06064_;
 wire _06065_;
 wire _06066_;
 wire _06067_;
 wire _06068_;
 wire _06069_;
 wire _06070_;
 wire _06071_;
 wire _06072_;
 wire _06073_;
 wire _06074_;
 wire _06075_;
 wire _06076_;
 wire _06077_;
 wire _06078_;
 wire _06079_;
 wire _06080_;
 wire _06081_;
 wire _06082_;
 wire _06083_;
 wire _06084_;
 wire _06085_;
 wire _06086_;
 wire _06087_;
 wire _06088_;
 wire _06089_;
 wire _06090_;
 wire _06091_;
 wire _06092_;
 wire _06093_;
 wire _06094_;
 wire _06095_;
 wire _06096_;
 wire _06097_;
 wire _06098_;
 wire _06099_;
 wire _06100_;
 wire _06101_;
 wire _06102_;
 wire _06103_;
 wire _06104_;
 wire _06105_;
 wire _06106_;
 wire _06107_;
 wire _06108_;
 wire _06109_;
 wire _06110_;
 wire _06111_;
 wire _06112_;
 wire _06113_;
 wire _06114_;
 wire _06115_;
 wire _06116_;
 wire _06117_;
 wire _06118_;
 wire _06119_;
 wire _06120_;
 wire _06121_;
 wire _06122_;
 wire _06123_;
 wire _06124_;
 wire _06125_;
 wire _06126_;
 wire _06127_;
 wire _06128_;
 wire _06129_;
 wire _06130_;
 wire _06131_;
 wire _06132_;
 wire _06133_;
 wire _06134_;
 wire _06135_;
 wire _06136_;
 wire _06137_;
 wire _06138_;
 wire _06139_;
 wire _06140_;
 wire _06141_;
 wire _06142_;
 wire _06143_;
 wire _06144_;
 wire _06145_;
 wire _06146_;
 wire _06147_;
 wire _06148_;
 wire _06149_;
 wire _06150_;
 wire _06151_;
 wire _06152_;
 wire _06153_;
 wire _06154_;
 wire _06155_;
 wire _06156_;
 wire _06157_;
 wire _06158_;
 wire _06159_;
 wire _06160_;
 wire _06161_;
 wire _06162_;
 wire _06163_;
 wire _06164_;
 wire _06165_;
 wire _06166_;
 wire _06167_;
 wire _06168_;
 wire _06169_;
 wire _06170_;
 wire _06171_;
 wire _06172_;
 wire _06173_;
 wire _06174_;
 wire _06175_;
 wire _06176_;
 wire _06177_;
 wire _06178_;
 wire _06179_;
 wire _06180_;
 wire _06181_;
 wire _06182_;
 wire _06183_;
 wire _06184_;
 wire _06185_;
 wire _06186_;
 wire _06187_;
 wire _06188_;
 wire _06189_;
 wire _06190_;
 wire _06191_;
 wire _06192_;
 wire _06193_;
 wire _06194_;
 wire _06195_;
 wire _06196_;
 wire _06197_;
 wire _06198_;
 wire _06199_;
 wire _06200_;
 wire _06201_;
 wire _06202_;
 wire _06203_;
 wire _06204_;
 wire _06205_;
 wire _06206_;
 wire _06207_;
 wire _06208_;
 wire _06209_;
 wire _06210_;
 wire _06211_;
 wire _06212_;
 wire _06213_;
 wire _06214_;
 wire _06215_;
 wire _06216_;
 wire _06217_;
 wire _06218_;
 wire _06219_;
 wire _06220_;
 wire _06221_;
 wire _06222_;
 wire _06223_;
 wire _06224_;
 wire _06225_;
 wire _06226_;
 wire _06227_;
 wire _06228_;
 wire _06229_;
 wire _06230_;
 wire _06231_;
 wire _06232_;
 wire _06233_;
 wire _06234_;
 wire _06235_;
 wire _06236_;
 wire _06237_;
 wire _06238_;
 wire _06239_;
 wire _06240_;
 wire _06241_;
 wire _06242_;
 wire _06243_;
 wire _06244_;
 wire _06245_;
 wire _06246_;
 wire _06247_;
 wire _06248_;
 wire _06249_;
 wire _06250_;
 wire _06251_;
 wire _06252_;
 wire _06253_;
 wire _06254_;
 wire _06255_;
 wire _06256_;
 wire _06257_;
 wire _06258_;
 wire _06259_;
 wire _06260_;
 wire _06261_;
 wire _06262_;
 wire _06263_;
 wire _06264_;
 wire _06265_;
 wire _06266_;
 wire _06267_;
 wire _06268_;
 wire _06269_;
 wire _06270_;
 wire _06271_;
 wire _06272_;
 wire _06273_;
 wire _06274_;
 wire _06275_;
 wire _06276_;
 wire _06277_;
 wire _06278_;
 wire _06279_;
 wire _06280_;
 wire _06281_;
 wire _06282_;
 wire _06283_;
 wire _06284_;
 wire _06285_;
 wire _06286_;
 wire _06287_;
 wire _06288_;
 wire _06289_;
 wire _06290_;
 wire _06291_;
 wire _06292_;
 wire _06293_;
 wire _06294_;
 wire _06295_;
 wire _06296_;
 wire _06297_;
 wire _06298_;
 wire _06299_;
 wire _06300_;
 wire _06301_;
 wire _06302_;
 wire _06303_;
 wire _06304_;
 wire _06305_;
 wire _06306_;
 wire _06307_;
 wire _06308_;
 wire _06309_;
 wire _06310_;
 wire _06311_;
 wire _06312_;
 wire _06313_;
 wire _06314_;
 wire _06315_;
 wire _06316_;
 wire _06317_;
 wire _06318_;
 wire _06319_;
 wire _06320_;
 wire _06321_;
 wire _06322_;
 wire _06323_;
 wire _06324_;
 wire _06325_;
 wire _06326_;
 wire _06327_;
 wire _06328_;
 wire _06329_;
 wire _06330_;
 wire _06331_;
 wire _06332_;
 wire _06333_;
 wire _06334_;
 wire _06335_;
 wire _06336_;
 wire _06337_;
 wire _06338_;
 wire _06339_;
 wire _06340_;
 wire _06341_;
 wire _06342_;
 wire _06343_;
 wire _06344_;
 wire _06345_;
 wire _06346_;
 wire _06347_;
 wire _06348_;
 wire _06349_;
 wire _06350_;
 wire _06351_;
 wire _06352_;
 wire _06353_;
 wire _06354_;
 wire _06355_;
 wire _06356_;
 wire _06357_;
 wire _06358_;
 wire _06359_;
 wire _06360_;
 wire _06361_;
 wire _06362_;
 wire _06363_;
 wire _06364_;
 wire _06365_;
 wire _06366_;
 wire _06367_;
 wire _06368_;
 wire _06369_;
 wire _06370_;
 wire _06371_;
 wire _06372_;
 wire _06373_;
 wire _06374_;
 wire _06375_;
 wire _06376_;
 wire _06377_;
 wire _06378_;
 wire _06379_;
 wire _06380_;
 wire _06381_;
 wire _06382_;
 wire _06383_;
 wire _06384_;
 wire _06385_;
 wire _06386_;
 wire _06387_;
 wire _06388_;
 wire _06389_;
 wire _06390_;
 wire _06391_;
 wire _06392_;
 wire _06393_;
 wire _06394_;
 wire _06395_;
 wire _06396_;
 wire _06397_;
 wire _06398_;
 wire _06399_;
 wire _06400_;
 wire _06401_;
 wire _06402_;
 wire _06403_;
 wire _06404_;
 wire _06405_;
 wire _06406_;
 wire _06407_;
 wire _06408_;
 wire _06409_;
 wire _06410_;
 wire _06411_;
 wire _06412_;
 wire _06413_;
 wire _06414_;
 wire _06415_;
 wire _06416_;
 wire _06417_;
 wire _06418_;
 wire _06419_;
 wire _06420_;
 wire _06421_;
 wire _06422_;
 wire _06423_;
 wire _06424_;
 wire _06425_;
 wire _06426_;
 wire _06427_;
 wire _06428_;
 wire _06429_;
 wire _06430_;
 wire _06431_;
 wire _06432_;
 wire _06433_;
 wire _06434_;
 wire _06435_;
 wire _06436_;
 wire _06437_;
 wire _06438_;
 wire _06439_;
 wire _06440_;
 wire _06441_;
 wire _06442_;
 wire _06443_;
 wire _06444_;
 wire _06445_;
 wire _06446_;
 wire _06447_;
 wire _06448_;
 wire _06449_;
 wire _06450_;
 wire _06451_;
 wire _06452_;
 wire _06453_;
 wire _06454_;
 wire _06455_;
 wire _06456_;
 wire _06457_;
 wire _06458_;
 wire _06459_;
 wire _06460_;
 wire _06461_;
 wire _06462_;
 wire _06463_;
 wire _06464_;
 wire _06465_;
 wire _06466_;
 wire _06467_;
 wire _06468_;
 wire _06469_;
 wire _06470_;
 wire _06471_;
 wire _06472_;
 wire _06473_;
 wire _06474_;
 wire _06475_;
 wire _06476_;
 wire _06477_;
 wire _06478_;
 wire _06479_;
 wire _06480_;
 wire _06481_;
 wire _06482_;
 wire _06483_;
 wire _06484_;
 wire _06485_;
 wire _06486_;
 wire _06487_;
 wire _06488_;
 wire _06489_;
 wire _06490_;
 wire _06491_;
 wire _06492_;
 wire _06493_;
 wire _06494_;
 wire _06495_;
 wire _06496_;
 wire _06497_;
 wire _06498_;
 wire _06499_;
 wire _06500_;
 wire _06501_;
 wire _06502_;
 wire _06503_;
 wire _06504_;
 wire _06505_;
 wire _06506_;
 wire _06507_;
 wire _06508_;
 wire _06509_;
 wire _06510_;
 wire _06511_;
 wire _06512_;
 wire _06513_;
 wire _06514_;
 wire _06515_;
 wire _06516_;
 wire _06517_;
 wire _06518_;
 wire _06519_;
 wire _06520_;
 wire _06521_;
 wire _06522_;
 wire _06523_;
 wire _06524_;
 wire _06525_;
 wire _06526_;
 wire _06527_;
 wire _06528_;
 wire _06529_;
 wire _06530_;
 wire _06531_;
 wire _06532_;
 wire _06533_;
 wire _06534_;
 wire _06535_;
 wire _06536_;
 wire _06537_;
 wire _06538_;
 wire _06539_;
 wire _06540_;
 wire _06541_;
 wire _06542_;
 wire _06543_;
 wire _06544_;
 wire _06545_;
 wire _06546_;
 wire _06547_;
 wire _06548_;
 wire _06549_;
 wire _06550_;
 wire _06551_;
 wire _06552_;
 wire _06553_;
 wire _06554_;
 wire _06555_;
 wire _06556_;
 wire _06557_;
 wire _06558_;
 wire _06559_;
 wire _06560_;
 wire _06561_;
 wire _06562_;
 wire _06563_;
 wire _06564_;
 wire _06565_;
 wire _06566_;
 wire _06567_;
 wire _06568_;
 wire _06569_;
 wire _06570_;
 wire _06571_;
 wire _06572_;
 wire _06573_;
 wire _06574_;
 wire _06575_;
 wire _06576_;
 wire _06577_;
 wire _06578_;
 wire _06579_;
 wire _06580_;
 wire _06581_;
 wire _06582_;
 wire _06583_;
 wire _06584_;
 wire _06585_;
 wire _06586_;
 wire _06587_;
 wire _06588_;
 wire _06589_;
 wire _06590_;
 wire _06591_;
 wire _06592_;
 wire _06593_;
 wire _06594_;
 wire _06595_;
 wire _06596_;
 wire _06597_;
 wire _06598_;
 wire _06599_;
 wire _06600_;
 wire _06601_;
 wire _06602_;
 wire _06603_;
 wire _06604_;
 wire _06605_;
 wire _06606_;
 wire _06607_;
 wire _06608_;
 wire _06609_;
 wire _06610_;
 wire _06611_;
 wire _06612_;
 wire _06613_;
 wire _06614_;
 wire _06615_;
 wire _06616_;
 wire _06617_;
 wire _06618_;
 wire _06619_;
 wire _06620_;
 wire _06621_;
 wire _06622_;
 wire _06623_;
 wire _06624_;
 wire _06625_;
 wire _06626_;
 wire _06627_;
 wire _06628_;
 wire _06629_;
 wire _06630_;
 wire _06631_;
 wire _06632_;
 wire _06633_;
 wire _06634_;
 wire _06635_;
 wire _06636_;
 wire _06637_;
 wire _06638_;
 wire _06639_;
 wire _06640_;
 wire _06641_;
 wire _06642_;
 wire _06643_;
 wire _06644_;
 wire _06645_;
 wire _06646_;
 wire _06647_;
 wire _06648_;
 wire _06649_;
 wire _06650_;
 wire _06651_;
 wire _06652_;
 wire _06653_;
 wire _06654_;
 wire _06655_;
 wire _06656_;
 wire _06657_;
 wire _06658_;
 wire _06659_;
 wire _06660_;
 wire _06661_;
 wire _06662_;
 wire _06663_;
 wire _06664_;
 wire _06665_;
 wire _06666_;
 wire _06667_;
 wire _06668_;
 wire _06669_;
 wire _06670_;
 wire _06671_;
 wire _06672_;
 wire _06673_;
 wire _06674_;
 wire _06675_;
 wire _06676_;
 wire _06677_;
 wire _06678_;
 wire _06679_;
 wire _06680_;
 wire _06681_;
 wire _06682_;
 wire _06683_;
 wire _06684_;
 wire _06685_;
 wire _06686_;
 wire _06687_;
 wire _06688_;
 wire _06689_;
 wire _06690_;
 wire _06691_;
 wire _06692_;
 wire _06693_;
 wire _06694_;
 wire _06695_;
 wire _06696_;
 wire _06697_;
 wire _06698_;
 wire _06699_;
 wire _06700_;
 wire _06701_;
 wire _06702_;
 wire _06703_;
 wire _06704_;
 wire _06705_;
 wire _06706_;
 wire _06707_;
 wire _06708_;
 wire _06709_;
 wire _06710_;
 wire _06711_;
 wire _06712_;
 wire _06713_;
 wire _06714_;
 wire _06715_;
 wire _06716_;
 wire _06717_;
 wire _06718_;
 wire _06719_;
 wire _06720_;
 wire _06721_;
 wire _06722_;
 wire _06723_;
 wire _06724_;
 wire _06725_;
 wire _06726_;
 wire _06727_;
 wire _06728_;
 wire _06729_;
 wire _06730_;
 wire _06731_;
 wire _06732_;
 wire _06733_;
 wire _06734_;
 wire _06735_;
 wire _06736_;
 wire _06737_;
 wire _06738_;
 wire _06739_;
 wire _06740_;
 wire _06741_;
 wire _06742_;
 wire _06743_;
 wire _06744_;
 wire _06745_;
 wire _06746_;
 wire _06747_;
 wire _06748_;
 wire _06749_;
 wire _06750_;
 wire _06751_;
 wire _06752_;
 wire _06753_;
 wire _06754_;
 wire _06755_;
 wire _06756_;
 wire _06757_;
 wire _06758_;
 wire _06759_;
 wire _06760_;
 wire _06761_;
 wire _06762_;
 wire _06763_;
 wire _06764_;
 wire _06765_;
 wire _06766_;
 wire _06767_;
 wire _06768_;
 wire _06769_;
 wire _06770_;
 wire _06771_;
 wire _06772_;
 wire _06773_;
 wire _06774_;
 wire _06775_;
 wire _06776_;
 wire _06777_;
 wire _06778_;
 wire _06779_;
 wire _06780_;
 wire _06781_;
 wire _06782_;
 wire _06783_;
 wire _06784_;
 wire _06785_;
 wire _06786_;
 wire _06787_;
 wire _06788_;
 wire _06789_;
 wire _06790_;
 wire _06791_;
 wire _06792_;
 wire _06793_;
 wire _06794_;
 wire _06795_;
 wire _06796_;
 wire _06797_;
 wire _06798_;
 wire _06799_;
 wire _06800_;
 wire _06801_;
 wire _06802_;
 wire _06803_;
 wire _06804_;
 wire _06805_;
 wire _06806_;
 wire _06807_;
 wire _06808_;
 wire _06809_;
 wire _06810_;
 wire _06811_;
 wire _06812_;
 wire _06813_;
 wire _06814_;
 wire _06815_;
 wire _06816_;
 wire _06817_;
 wire _06818_;
 wire _06819_;
 wire _06820_;
 wire _06821_;
 wire _06822_;
 wire _06823_;
 wire _06824_;
 wire _06825_;
 wire _06826_;
 wire _06827_;
 wire _06828_;
 wire _06829_;
 wire _06830_;
 wire _06831_;
 wire _06832_;
 wire _06833_;
 wire _06834_;
 wire _06835_;
 wire _06836_;
 wire _06837_;
 wire _06838_;
 wire _06839_;
 wire _06840_;
 wire _06841_;
 wire _06842_;
 wire _06843_;
 wire _06844_;
 wire _06845_;
 wire _06846_;
 wire _06847_;
 wire _06848_;
 wire _06849_;
 wire _06850_;
 wire _06851_;
 wire _06852_;
 wire _06853_;
 wire _06854_;
 wire _06855_;
 wire _06856_;
 wire _06857_;
 wire _06858_;
 wire _06859_;
 wire _06860_;
 wire _06861_;
 wire _06862_;
 wire _06863_;
 wire _06864_;
 wire _06865_;
 wire _06866_;
 wire _06867_;
 wire _06868_;
 wire _06869_;
 wire _06870_;
 wire _06871_;
 wire _06872_;
 wire _06873_;
 wire _06874_;
 wire _06875_;
 wire _06876_;
 wire _06877_;
 wire _06878_;
 wire _06879_;
 wire _06880_;
 wire _06881_;
 wire _06882_;
 wire _06883_;
 wire _06884_;
 wire _06885_;
 wire _06886_;
 wire _06887_;
 wire _06888_;
 wire _06889_;
 wire _06890_;
 wire _06891_;
 wire _06892_;
 wire _06893_;
 wire _06894_;
 wire _06895_;
 wire _06896_;
 wire _06897_;
 wire _06898_;
 wire _06899_;
 wire _06900_;
 wire _06901_;
 wire _06902_;
 wire _06903_;
 wire _06904_;
 wire _06905_;
 wire _06906_;
 wire _06907_;
 wire _06908_;
 wire _06909_;
 wire _06910_;
 wire _06911_;
 wire _06912_;
 wire _06913_;
 wire _06914_;
 wire _06915_;
 wire _06916_;
 wire _06917_;
 wire _06918_;
 wire _06919_;
 wire _06920_;
 wire _06921_;
 wire _06922_;
 wire _06923_;
 wire _06924_;
 wire _06925_;
 wire _06926_;
 wire _06927_;
 wire _06928_;
 wire _06929_;
 wire _06930_;
 wire _06931_;
 wire _06932_;
 wire _06933_;
 wire _06934_;
 wire _06935_;
 wire _06936_;
 wire _06937_;
 wire _06938_;
 wire _06939_;
 wire _06940_;
 wire _06941_;
 wire _06942_;
 wire _06943_;
 wire _06944_;
 wire _06945_;
 wire _06946_;
 wire _06947_;
 wire _06948_;
 wire _06949_;
 wire _06950_;
 wire _06951_;
 wire _06952_;
 wire _06953_;
 wire _06954_;
 wire _06955_;
 wire _06956_;
 wire _06957_;
 wire _06958_;
 wire _06959_;
 wire _06960_;
 wire _06961_;
 wire _06962_;
 wire _06963_;
 wire _06964_;
 wire _06965_;
 wire _06966_;
 wire _06967_;
 wire _06968_;
 wire _06969_;
 wire _06970_;
 wire _06971_;
 wire _06972_;
 wire _06973_;
 wire _06974_;
 wire _06975_;
 wire _06976_;
 wire _06977_;
 wire _06978_;
 wire _06979_;
 wire _06980_;
 wire _06981_;
 wire _06982_;
 wire _06983_;
 wire _06984_;
 wire _06985_;
 wire _06986_;
 wire _06987_;
 wire _06988_;
 wire _06989_;
 wire _06990_;
 wire _06991_;
 wire _06992_;
 wire _06993_;
 wire _06994_;
 wire _06995_;
 wire _06996_;
 wire _06997_;
 wire _06998_;
 wire _06999_;
 wire _07000_;
 wire _07001_;
 wire _07002_;
 wire _07003_;
 wire _07004_;
 wire _07005_;
 wire _07006_;
 wire _07007_;
 wire _07008_;
 wire _07009_;
 wire _07010_;
 wire _07011_;
 wire _07012_;
 wire _07013_;
 wire _07014_;
 wire _07015_;
 wire _07016_;
 wire _07017_;
 wire _07018_;
 wire _07019_;
 wire _07020_;
 wire _07021_;
 wire _07022_;
 wire _07023_;
 wire _07024_;
 wire _07025_;
 wire _07026_;
 wire _07027_;
 wire _07028_;
 wire _07029_;
 wire _07030_;
 wire _07031_;
 wire _07032_;
 wire _07033_;
 wire _07034_;
 wire _07035_;
 wire _07036_;
 wire _07037_;
 wire _07038_;
 wire _07039_;
 wire _07040_;
 wire _07041_;
 wire _07042_;
 wire _07043_;
 wire _07044_;
 wire _07045_;
 wire _07046_;
 wire _07047_;
 wire _07048_;
 wire _07049_;
 wire _07050_;
 wire _07051_;
 wire _07052_;
 wire _07053_;
 wire _07054_;
 wire _07055_;
 wire _07056_;
 wire _07057_;
 wire _07058_;
 wire _07059_;
 wire _07060_;
 wire _07061_;
 wire _07062_;
 wire _07063_;
 wire _07064_;
 wire _07065_;
 wire _07066_;
 wire _07067_;
 wire _07068_;
 wire _07069_;
 wire _07070_;
 wire _07071_;
 wire _07072_;
 wire _07073_;
 wire _07074_;
 wire _07075_;
 wire _07076_;
 wire _07077_;
 wire _07078_;
 wire _07079_;
 wire _07080_;
 wire _07081_;
 wire _07082_;
 wire _07083_;
 wire _07084_;
 wire _07085_;
 wire _07086_;
 wire _07087_;
 wire _07088_;
 wire _07089_;
 wire _07090_;
 wire _07091_;
 wire _07092_;
 wire _07093_;
 wire _07094_;
 wire _07095_;
 wire _07096_;
 wire _07097_;
 wire _07098_;
 wire _07099_;
 wire _07100_;
 wire _07101_;
 wire _07102_;
 wire _07103_;
 wire _07104_;
 wire _07105_;
 wire _07106_;
 wire _07107_;
 wire _07108_;
 wire _07109_;
 wire _07110_;
 wire _07111_;
 wire _07112_;
 wire _07113_;
 wire _07114_;
 wire _07115_;
 wire _07116_;
 wire _07117_;
 wire _07118_;
 wire _07119_;
 wire _07120_;
 wire _07121_;
 wire _07122_;
 wire _07123_;
 wire _07124_;
 wire _07125_;
 wire _07126_;
 wire _07127_;
 wire _07128_;
 wire _07129_;
 wire _07130_;
 wire _07131_;
 wire _07132_;
 wire _07133_;
 wire _07134_;
 wire _07135_;
 wire _07136_;
 wire _07137_;
 wire _07138_;
 wire _07139_;
 wire _07140_;
 wire _07141_;
 wire _07142_;
 wire _07143_;
 wire _07144_;
 wire _07145_;
 wire _07146_;
 wire _07147_;
 wire _07148_;
 wire _07149_;
 wire _07150_;
 wire _07151_;
 wire _07152_;
 wire _07153_;
 wire _07154_;
 wire _07155_;
 wire _07156_;
 wire _07157_;
 wire _07158_;
 wire _07159_;
 wire _07160_;
 wire _07161_;
 wire _07162_;
 wire _07163_;
 wire _07164_;
 wire _07165_;
 wire _07166_;
 wire _07167_;
 wire _07168_;
 wire _07169_;
 wire _07170_;
 wire _07171_;
 wire _07172_;
 wire _07173_;
 wire _07174_;
 wire _07175_;
 wire _07176_;
 wire _07177_;
 wire _07178_;
 wire _07179_;
 wire _07180_;
 wire _07181_;
 wire _07182_;
 wire _07183_;
 wire _07184_;
 wire _07185_;
 wire _07186_;
 wire _07187_;
 wire _07188_;
 wire _07189_;
 wire _07190_;
 wire _07191_;
 wire _07192_;
 wire _07193_;
 wire _07194_;
 wire _07195_;
 wire _07196_;
 wire _07197_;
 wire _07198_;
 wire _07199_;
 wire _07200_;
 wire _07201_;
 wire _07202_;
 wire _07203_;
 wire _07204_;
 wire _07205_;
 wire _07206_;
 wire _07207_;
 wire _07208_;
 wire _07209_;
 wire _07210_;
 wire _07211_;
 wire _07212_;
 wire _07213_;
 wire _07214_;
 wire _07215_;
 wire _07216_;
 wire _07217_;
 wire _07218_;
 wire _07219_;
 wire _07220_;
 wire _07221_;
 wire _07222_;
 wire _07223_;
 wire _07224_;
 wire _07225_;
 wire _07226_;
 wire _07227_;
 wire _07228_;
 wire _07229_;
 wire _07230_;
 wire _07231_;
 wire _07232_;
 wire _07233_;
 wire _07234_;
 wire _07235_;
 wire _07236_;
 wire _07237_;
 wire _07238_;
 wire _07239_;
 wire _07240_;
 wire _07241_;
 wire _07242_;
 wire _07243_;
 wire _07244_;
 wire _07245_;
 wire _07246_;
 wire _07247_;
 wire _07248_;
 wire _07249_;
 wire _07250_;
 wire _07251_;
 wire _07252_;
 wire _07253_;
 wire _07254_;
 wire _07255_;
 wire _07256_;
 wire _07257_;
 wire _07258_;
 wire _07259_;
 wire _07260_;
 wire _07261_;
 wire _07262_;
 wire _07263_;
 wire _07264_;
 wire _07265_;
 wire _07266_;
 wire _07267_;
 wire _07268_;
 wire _07269_;
 wire _07270_;
 wire _07271_;
 wire _07272_;
 wire _07273_;
 wire _07274_;
 wire _07275_;
 wire _07276_;
 wire _07277_;
 wire _07278_;
 wire _07279_;
 wire _07280_;
 wire _07281_;
 wire _07282_;
 wire _07283_;
 wire _07284_;
 wire _07285_;
 wire _07286_;
 wire _07287_;
 wire _07288_;
 wire _07289_;
 wire _07290_;
 wire _07291_;
 wire _07292_;
 wire _07293_;
 wire _07294_;
 wire _07295_;
 wire _07296_;
 wire _07297_;
 wire _07298_;
 wire _07299_;
 wire _07300_;
 wire _07301_;
 wire _07302_;
 wire _07303_;
 wire _07304_;
 wire _07305_;
 wire _07306_;
 wire _07307_;
 wire _07308_;
 wire _07309_;
 wire _07310_;
 wire _07311_;
 wire _07312_;
 wire _07313_;
 wire _07314_;
 wire _07315_;
 wire _07316_;
 wire _07317_;
 wire _07318_;
 wire _07319_;
 wire _07320_;
 wire _07321_;
 wire _07322_;
 wire _07323_;
 wire _07324_;
 wire _07325_;
 wire _07326_;
 wire _07327_;
 wire _07328_;
 wire _07329_;
 wire _07330_;
 wire _07331_;
 wire _07332_;
 wire _07333_;
 wire _07334_;
 wire _07335_;
 wire _07336_;
 wire _07337_;
 wire _07338_;
 wire _07339_;
 wire _07340_;
 wire _07341_;
 wire _07342_;
 wire _07343_;
 wire _07344_;
 wire _07345_;
 wire _07346_;
 wire _07347_;
 wire _07348_;
 wire _07349_;
 wire _07350_;
 wire _07351_;
 wire _07352_;
 wire _07353_;
 wire _07354_;
 wire _07355_;
 wire _07356_;
 wire _07357_;
 wire _07358_;
 wire _07359_;
 wire _07360_;
 wire _07361_;
 wire _07362_;
 wire _07363_;
 wire _07364_;
 wire _07365_;
 wire _07366_;
 wire _07367_;
 wire _07368_;
 wire _07369_;
 wire _07370_;
 wire _07371_;
 wire _07372_;
 wire _07373_;
 wire _07374_;
 wire _07375_;
 wire _07376_;
 wire _07377_;
 wire _07378_;
 wire _07379_;
 wire _07380_;
 wire _07381_;
 wire _07382_;
 wire _07383_;
 wire _07384_;
 wire _07385_;
 wire _07386_;
 wire _07387_;
 wire _07388_;
 wire _07389_;
 wire _07390_;
 wire _07391_;
 wire _07392_;
 wire _07393_;
 wire _07394_;
 wire _07395_;
 wire _07396_;
 wire _07397_;
 wire _07398_;
 wire _07399_;
 wire _07400_;
 wire _07401_;
 wire _07402_;
 wire _07403_;
 wire _07404_;
 wire _07405_;
 wire _07406_;
 wire _07407_;
 wire _07408_;
 wire _07409_;
 wire _07410_;
 wire _07411_;
 wire _07412_;
 wire _07413_;
 wire _07414_;
 wire _07415_;
 wire _07416_;
 wire _07417_;
 wire _07418_;
 wire _07419_;
 wire _07420_;
 wire _07421_;
 wire _07422_;
 wire _07423_;
 wire _07424_;
 wire _07425_;
 wire _07426_;
 wire _07427_;
 wire _07428_;
 wire _07429_;
 wire _07430_;
 wire _07431_;
 wire _07432_;
 wire _07433_;
 wire _07434_;
 wire _07435_;
 wire _07436_;
 wire _07437_;
 wire _07438_;
 wire _07439_;
 wire _07440_;
 wire _07441_;
 wire _07442_;
 wire _07443_;
 wire _07444_;
 wire _07445_;
 wire _07446_;
 wire _07447_;
 wire _07448_;
 wire _07449_;
 wire _07450_;
 wire _07451_;
 wire _07452_;
 wire _07453_;
 wire _07454_;
 wire _07455_;
 wire _07456_;
 wire _07457_;
 wire _07458_;
 wire _07459_;
 wire _07460_;
 wire _07461_;
 wire _07462_;
 wire _07463_;
 wire _07464_;
 wire _07465_;
 wire _07466_;
 wire _07467_;
 wire _07468_;
 wire _07469_;
 wire _07470_;
 wire _07471_;
 wire _07472_;
 wire _07473_;
 wire _07474_;
 wire _07475_;
 wire _07476_;
 wire _07477_;
 wire _07478_;
 wire _07479_;
 wire _07480_;
 wire _07481_;
 wire _07482_;
 wire _07483_;
 wire _07484_;
 wire _07485_;
 wire _07486_;
 wire _07487_;
 wire _07488_;
 wire _07489_;
 wire _07490_;
 wire _07491_;
 wire _07492_;
 wire _07493_;
 wire _07494_;
 wire _07495_;
 wire _07496_;
 wire _07497_;
 wire _07498_;
 wire _07499_;
 wire _07500_;
 wire _07501_;
 wire _07502_;
 wire _07503_;
 wire _07504_;
 wire _07505_;
 wire _07506_;
 wire _07507_;
 wire _07508_;
 wire _07509_;
 wire _07510_;
 wire _07511_;
 wire _07512_;
 wire _07513_;
 wire _07514_;
 wire _07515_;
 wire _07516_;
 wire _07517_;
 wire _07518_;
 wire _07519_;
 wire _07520_;
 wire _07521_;
 wire _07522_;
 wire _07523_;
 wire _07524_;
 wire _07525_;
 wire _07526_;
 wire _07527_;
 wire _07528_;
 wire _07529_;
 wire _07530_;
 wire _07531_;
 wire _07532_;
 wire _07533_;
 wire _07534_;
 wire _07535_;
 wire _07536_;
 wire _07537_;
 wire _07538_;
 wire _07539_;
 wire _07540_;
 wire _07541_;
 wire _07542_;
 wire _07543_;
 wire _07544_;
 wire _07545_;
 wire _07546_;
 wire _07547_;
 wire _07548_;
 wire _07549_;
 wire _07550_;
 wire _07551_;
 wire _07552_;
 wire _07553_;
 wire _07554_;
 wire _07555_;
 wire _07556_;
 wire _07557_;
 wire _07558_;
 wire _07559_;
 wire _07560_;
 wire _07561_;
 wire _07562_;
 wire _07563_;
 wire _07564_;
 wire _07565_;
 wire _07566_;
 wire _07567_;
 wire _07568_;
 wire _07569_;
 wire _07570_;
 wire _07571_;
 wire _07572_;
 wire _07573_;
 wire _07574_;
 wire _07575_;
 wire _07576_;
 wire _07577_;
 wire _07578_;
 wire _07579_;
 wire _07580_;
 wire _07581_;
 wire _07582_;
 wire _07583_;
 wire _07584_;
 wire _07585_;
 wire _07586_;
 wire _07587_;
 wire _07588_;
 wire _07589_;
 wire _07590_;
 wire _07591_;
 wire _07592_;
 wire _07593_;
 wire _07594_;
 wire _07595_;
 wire _07596_;
 wire _07597_;
 wire _07598_;
 wire _07599_;
 wire _07600_;
 wire _07601_;
 wire _07602_;
 wire _07603_;
 wire _07604_;
 wire _07605_;
 wire _07606_;
 wire _07607_;
 wire _07608_;
 wire _07609_;
 wire _07610_;
 wire _07611_;
 wire _07612_;
 wire _07613_;
 wire _07614_;
 wire _07615_;
 wire _07616_;
 wire _07617_;
 wire _07618_;
 wire _07619_;
 wire _07620_;
 wire _07621_;
 wire _07622_;
 wire _07623_;
 wire _07624_;
 wire _07625_;
 wire _07626_;
 wire _07627_;
 wire _07628_;
 wire _07629_;
 wire _07630_;
 wire _07631_;
 wire _07632_;
 wire _07633_;
 wire _07634_;
 wire _07635_;
 wire _07636_;
 wire _07637_;
 wire _07638_;
 wire _07639_;
 wire _07640_;
 wire _07641_;
 wire _07642_;
 wire _07643_;
 wire _07644_;
 wire _07645_;
 wire _07646_;
 wire _07647_;
 wire _07648_;
 wire _07649_;
 wire _07650_;
 wire _07651_;
 wire _07652_;
 wire _07653_;
 wire _07654_;
 wire _07655_;
 wire _07656_;
 wire _07657_;
 wire _07658_;
 wire _07659_;
 wire _07660_;
 wire _07661_;
 wire _07662_;
 wire _07663_;
 wire _07664_;
 wire _07665_;
 wire _07666_;
 wire _07667_;
 wire _07668_;
 wire _07669_;
 wire _07670_;
 wire _07671_;
 wire _07672_;
 wire _07673_;
 wire _07674_;
 wire _07675_;
 wire _07676_;
 wire _07677_;
 wire _07678_;
 wire _07679_;
 wire _07680_;
 wire _07681_;
 wire _07682_;
 wire _07683_;
 wire _07684_;
 wire _07685_;
 wire _07686_;
 wire _07687_;
 wire _07688_;
 wire _07689_;
 wire _07690_;
 wire _07691_;
 wire _07692_;
 wire _07693_;
 wire _07694_;
 wire _07695_;
 wire _07696_;
 wire _07697_;
 wire _07698_;
 wire _07699_;
 wire _07700_;
 wire _07701_;
 wire _07702_;
 wire _07703_;
 wire _07704_;
 wire _07705_;
 wire _07706_;
 wire _07707_;
 wire _07708_;
 wire _07709_;
 wire _07710_;
 wire _07711_;
 wire _07712_;
 wire _07713_;
 wire _07714_;
 wire _07715_;
 wire _07716_;
 wire _07717_;
 wire _07718_;
 wire _07719_;
 wire _07720_;
 wire _07721_;
 wire _07722_;
 wire _07723_;
 wire _07724_;
 wire _07725_;
 wire _07726_;
 wire _07727_;
 wire _07728_;
 wire _07729_;
 wire _07730_;
 wire _07731_;
 wire _07732_;
 wire _07733_;
 wire _07734_;
 wire _07735_;
 wire _07736_;
 wire _07737_;
 wire _07738_;
 wire _07739_;
 wire _07740_;
 wire _07741_;
 wire _07742_;
 wire _07743_;
 wire _07744_;
 wire _07745_;
 wire _07746_;
 wire _07747_;
 wire _07748_;
 wire _07749_;
 wire _07750_;
 wire _07751_;
 wire _07752_;
 wire _07753_;
 wire _07754_;
 wire _07755_;
 wire _07756_;
 wire _07757_;
 wire _07758_;
 wire _07759_;
 wire _07760_;
 wire _07761_;
 wire _07762_;
 wire _07763_;
 wire _07764_;
 wire _07765_;
 wire _07766_;
 wire _07767_;
 wire _07768_;
 wire _07769_;
 wire _07770_;
 wire _07771_;
 wire _07772_;
 wire _07773_;
 wire _07774_;
 wire _07775_;
 wire _07776_;
 wire _07777_;
 wire _07778_;
 wire _07779_;
 wire _07780_;
 wire _07781_;
 wire _07782_;
 wire _07783_;
 wire _07784_;
 wire _07785_;
 wire _07786_;
 wire _07787_;
 wire _07788_;
 wire _07789_;
 wire _07790_;
 wire _07791_;
 wire _07792_;
 wire _07793_;
 wire _07794_;
 wire _07795_;
 wire _07796_;
 wire _07797_;
 wire _07798_;
 wire _07799_;
 wire _07800_;
 wire _07801_;
 wire _07802_;
 wire _07803_;
 wire _07804_;
 wire _07805_;
 wire _07806_;
 wire _07807_;
 wire _07808_;
 wire _07809_;
 wire _07810_;
 wire _07811_;
 wire _07812_;
 wire _07813_;
 wire _07814_;
 wire _07815_;
 wire _07816_;
 wire _07817_;
 wire _07818_;
 wire _07819_;
 wire _07820_;
 wire _07821_;
 wire _07822_;
 wire _07823_;
 wire _07824_;
 wire _07825_;
 wire _07826_;
 wire _07827_;
 wire _07828_;
 wire _07829_;
 wire _07830_;
 wire _07831_;
 wire _07832_;
 wire _07833_;
 wire _07834_;
 wire _07835_;
 wire _07836_;
 wire _07837_;
 wire _07838_;
 wire _07839_;
 wire _07840_;
 wire _07841_;
 wire _07842_;
 wire _07843_;
 wire _07844_;
 wire _07845_;
 wire _07846_;
 wire _07847_;
 wire _07848_;
 wire _07849_;
 wire _07850_;
 wire _07851_;
 wire _07852_;
 wire _07853_;
 wire _07854_;
 wire _07855_;
 wire _07856_;
 wire _07857_;
 wire _07858_;
 wire _07859_;
 wire _07860_;
 wire _07861_;
 wire _07862_;
 wire _07863_;
 wire _07864_;
 wire _07865_;
 wire _07866_;
 wire _07867_;
 wire _07868_;
 wire _07869_;
 wire _07870_;
 wire _07871_;
 wire _07872_;
 wire _07873_;
 wire _07874_;
 wire _07875_;
 wire _07876_;
 wire _07877_;
 wire _07878_;
 wire _07879_;
 wire _07880_;
 wire _07881_;
 wire _07882_;
 wire _07883_;
 wire _07884_;
 wire _07885_;
 wire _07886_;
 wire _07887_;
 wire _07888_;
 wire _07889_;
 wire _07890_;
 wire _07891_;
 wire _07892_;
 wire _07893_;
 wire _07894_;
 wire _07895_;
 wire _07896_;
 wire _07897_;
 wire _07898_;
 wire _07899_;
 wire _07900_;
 wire _07901_;
 wire _07902_;
 wire _07903_;
 wire _07904_;
 wire _07905_;
 wire _07906_;
 wire _07907_;
 wire _07908_;
 wire _07909_;
 wire _07910_;
 wire _07911_;
 wire _07912_;
 wire _07913_;
 wire _07914_;
 wire _07915_;
 wire _07916_;
 wire _07917_;
 wire _07918_;
 wire _07919_;
 wire _07920_;
 wire _07921_;
 wire _07922_;
 wire _07923_;
 wire _07924_;
 wire _07925_;
 wire _07926_;
 wire _07927_;
 wire _07928_;
 wire _07929_;
 wire _07930_;
 wire _07931_;
 wire _07932_;
 wire _07933_;
 wire _07934_;
 wire _07935_;
 wire _07936_;
 wire _07937_;
 wire _07938_;
 wire _07939_;
 wire _07940_;
 wire _07941_;
 wire _07942_;
 wire _07943_;
 wire _07944_;
 wire _07945_;
 wire _07946_;
 wire _07947_;
 wire _07948_;
 wire _07949_;
 wire _07950_;
 wire _07951_;
 wire _07952_;
 wire _07953_;
 wire _07954_;
 wire _07955_;
 wire _07956_;
 wire _07957_;
 wire _07958_;
 wire _07959_;
 wire _07960_;
 wire _07961_;
 wire _07962_;
 wire _07963_;
 wire _07964_;
 wire _07965_;
 wire _07966_;
 wire _07967_;
 wire _07968_;
 wire _07969_;
 wire _07970_;
 wire _07971_;
 wire _07972_;
 wire _07973_;
 wire _07974_;
 wire _07975_;
 wire _07976_;
 wire _07977_;
 wire _07978_;
 wire _07979_;
 wire _07980_;
 wire _07981_;
 wire _07982_;
 wire _07983_;
 wire _07984_;
 wire _07985_;
 wire _07986_;
 wire _07987_;
 wire _07988_;
 wire _07989_;
 wire _07990_;
 wire _07991_;
 wire _07992_;
 wire _07993_;
 wire _07994_;
 wire _07995_;
 wire _07996_;
 wire _07997_;
 wire _07998_;
 wire _07999_;
 wire _08000_;
 wire _08001_;
 wire _08002_;
 wire _08003_;
 wire _08004_;
 wire _08005_;
 wire _08006_;
 wire _08007_;
 wire _08008_;
 wire _08009_;
 wire _08010_;
 wire _08011_;
 wire _08012_;
 wire _08013_;
 wire _08014_;
 wire _08015_;
 wire _08016_;
 wire _08017_;
 wire _08018_;
 wire _08019_;
 wire _08020_;
 wire _08021_;
 wire _08022_;
 wire _08023_;
 wire _08024_;
 wire _08025_;
 wire _08026_;
 wire _08027_;
 wire _08028_;
 wire _08029_;
 wire _08030_;
 wire _08031_;
 wire _08032_;
 wire _08033_;
 wire _08034_;
 wire _08035_;
 wire _08036_;
 wire _08037_;
 wire _08038_;
 wire _08039_;
 wire _08040_;
 wire _08041_;
 wire _08042_;
 wire _08043_;
 wire _08044_;
 wire _08045_;
 wire _08046_;
 wire _08047_;
 wire _08048_;
 wire _08049_;
 wire _08050_;
 wire _08051_;
 wire _08052_;
 wire _08053_;
 wire _08054_;
 wire _08055_;
 wire _08056_;
 wire _08057_;
 wire _08058_;
 wire _08059_;
 wire _08060_;
 wire _08061_;
 wire _08062_;
 wire _08063_;
 wire _08064_;
 wire _08065_;
 wire _08066_;
 wire _08067_;
 wire _08068_;
 wire _08069_;
 wire _08070_;
 wire _08071_;
 wire _08072_;
 wire _08073_;
 wire _08074_;
 wire _08075_;
 wire _08076_;
 wire _08077_;
 wire _08078_;
 wire _08079_;
 wire _08080_;
 wire _08081_;
 wire _08082_;
 wire _08083_;
 wire _08084_;
 wire _08085_;
 wire _08086_;
 wire _08087_;
 wire _08088_;
 wire _08089_;
 wire _08090_;
 wire _08091_;
 wire _08092_;
 wire _08093_;
 wire _08094_;
 wire _08095_;
 wire _08096_;
 wire _08097_;
 wire _08098_;
 wire _08099_;
 wire _08100_;
 wire _08101_;
 wire _08102_;
 wire _08103_;
 wire _08104_;
 wire _08105_;
 wire _08106_;
 wire _08107_;
 wire _08108_;
 wire _08109_;
 wire _08110_;
 wire _08111_;
 wire _08112_;
 wire _08113_;
 wire _08114_;
 wire _08115_;
 wire _08116_;
 wire _08117_;
 wire _08118_;
 wire _08119_;
 wire _08120_;
 wire _08121_;
 wire _08122_;
 wire _08123_;
 wire _08124_;
 wire _08125_;
 wire _08126_;
 wire _08127_;
 wire _08128_;
 wire _08129_;
 wire _08130_;
 wire _08131_;
 wire _08132_;
 wire _08133_;
 wire _08134_;
 wire _08135_;
 wire _08136_;
 wire _08137_;
 wire _08138_;
 wire _08139_;
 wire _08140_;
 wire _08141_;
 wire _08142_;
 wire _08143_;
 wire _08144_;
 wire _08145_;
 wire _08146_;
 wire _08147_;
 wire _08148_;
 wire _08149_;
 wire _08150_;
 wire _08151_;
 wire _08152_;
 wire _08153_;
 wire _08154_;
 wire _08155_;
 wire _08156_;
 wire _08157_;
 wire _08158_;
 wire _08159_;
 wire _08160_;
 wire _08161_;
 wire _08162_;
 wire _08163_;
 wire _08164_;
 wire _08165_;
 wire _08166_;
 wire _08167_;
 wire _08168_;
 wire _08169_;
 wire _08170_;
 wire _08171_;
 wire _08172_;
 wire _08173_;
 wire _08174_;
 wire _08175_;
 wire _08176_;
 wire _08177_;
 wire _08178_;
 wire _08179_;
 wire _08180_;
 wire _08181_;
 wire _08182_;
 wire _08183_;
 wire _08184_;
 wire _08185_;
 wire _08186_;
 wire _08187_;
 wire _08188_;
 wire _08189_;
 wire _08190_;
 wire _08191_;
 wire _08192_;
 wire _08193_;
 wire _08194_;
 wire _08195_;
 wire _08196_;
 wire _08197_;
 wire _08198_;
 wire _08199_;
 wire _08200_;
 wire _08201_;
 wire _08202_;
 wire _08203_;
 wire _08204_;
 wire _08205_;
 wire _08206_;
 wire _08207_;
 wire _08208_;
 wire _08209_;
 wire _08210_;
 wire _08211_;
 wire _08212_;
 wire _08213_;
 wire _08214_;
 wire _08215_;
 wire _08216_;
 wire _08217_;
 wire _08218_;
 wire _08219_;
 wire _08220_;
 wire _08221_;
 wire _08222_;
 wire _08223_;
 wire _08224_;
 wire _08225_;
 wire _08226_;
 wire _08227_;
 wire _08228_;
 wire _08229_;
 wire _08230_;
 wire _08231_;
 wire _08232_;
 wire _08233_;
 wire _08234_;
 wire _08235_;
 wire _08236_;
 wire _08237_;
 wire _08238_;
 wire _08239_;
 wire _08240_;
 wire _08241_;
 wire _08242_;
 wire _08243_;
 wire _08244_;
 wire _08245_;
 wire _08246_;
 wire _08247_;
 wire _08248_;
 wire _08249_;
 wire _08250_;
 wire _08251_;
 wire _08252_;
 wire _08253_;
 wire _08254_;
 wire _08255_;
 wire _08256_;
 wire _08257_;
 wire _08258_;
 wire _08259_;
 wire _08260_;
 wire _08261_;
 wire _08262_;
 wire _08263_;
 wire _08264_;
 wire _08265_;
 wire _08266_;
 wire _08267_;
 wire _08268_;
 wire _08269_;
 wire _08270_;
 wire _08271_;
 wire _08272_;
 wire _08273_;
 wire _08274_;
 wire _08275_;
 wire _08276_;
 wire _08277_;
 wire _08278_;
 wire _08279_;
 wire _08280_;
 wire _08281_;
 wire _08282_;
 wire _08283_;
 wire _08284_;
 wire _08285_;
 wire _08286_;
 wire _08287_;
 wire _08288_;
 wire _08289_;
 wire _08290_;
 wire _08291_;
 wire _08292_;
 wire _08293_;
 wire _08294_;
 wire _08295_;
 wire _08296_;
 wire _08297_;
 wire _08298_;
 wire _08299_;
 wire _08300_;
 wire _08301_;
 wire _08302_;
 wire _08303_;
 wire _08304_;
 wire _08305_;
 wire _08306_;
 wire _08307_;
 wire _08308_;
 wire _08309_;
 wire _08310_;
 wire _08311_;
 wire _08312_;
 wire _08313_;
 wire _08314_;
 wire _08315_;
 wire _08316_;
 wire _08317_;
 wire _08318_;
 wire _08319_;
 wire _08320_;
 wire _08321_;
 wire _08322_;
 wire _08323_;
 wire _08324_;
 wire _08325_;
 wire _08326_;
 wire _08327_;
 wire _08328_;
 wire _08329_;
 wire _08330_;
 wire _08331_;
 wire _08332_;
 wire _08333_;
 wire _08334_;
 wire _08335_;
 wire _08336_;
 wire _08337_;
 wire _08338_;
 wire _08339_;
 wire _08340_;
 wire _08341_;
 wire _08342_;
 wire _08343_;
 wire _08344_;
 wire _08345_;
 wire _08346_;
 wire _08347_;
 wire _08348_;
 wire _08349_;
 wire _08350_;
 wire _08351_;
 wire _08352_;
 wire _08353_;
 wire _08354_;
 wire _08355_;
 wire _08356_;
 wire _08357_;
 wire _08358_;
 wire _08359_;
 wire _08360_;
 wire _08361_;
 wire _08362_;
 wire _08363_;
 wire _08364_;
 wire _08365_;
 wire _08366_;
 wire _08367_;
 wire _08368_;
 wire _08369_;
 wire _08370_;
 wire _08371_;
 wire _08372_;
 wire _08373_;
 wire _08374_;
 wire _08375_;
 wire _08376_;
 wire _08377_;
 wire _08378_;
 wire _08379_;
 wire _08380_;
 wire _08381_;
 wire _08382_;
 wire _08383_;
 wire _08384_;
 wire _08385_;
 wire _08386_;
 wire _08387_;
 wire _08388_;
 wire _08389_;
 wire _08390_;
 wire _08391_;
 wire _08392_;
 wire _08393_;
 wire _08394_;
 wire _08395_;
 wire _08396_;
 wire _08397_;
 wire _08398_;
 wire _08399_;
 wire _08400_;
 wire _08401_;
 wire _08402_;
 wire _08403_;
 wire _08404_;
 wire _08405_;
 wire _08406_;
 wire _08407_;
 wire _08408_;
 wire _08409_;
 wire _08410_;
 wire _08411_;
 wire _08412_;
 wire _08413_;
 wire _08414_;
 wire _08415_;
 wire _08416_;
 wire _08417_;
 wire _08418_;
 wire _08419_;
 wire _08420_;
 wire _08421_;
 wire _08422_;
 wire _08423_;
 wire _08424_;
 wire _08425_;
 wire _08426_;
 wire _08427_;
 wire _08428_;
 wire _08429_;
 wire _08430_;
 wire _08431_;
 wire _08432_;
 wire _08433_;
 wire _08434_;
 wire _08435_;
 wire _08436_;
 wire _08437_;
 wire _08438_;
 wire _08439_;
 wire _08440_;
 wire _08441_;
 wire _08442_;
 wire _08443_;
 wire _08444_;
 wire _08445_;
 wire _08446_;
 wire _08447_;
 wire _08448_;
 wire _08449_;
 wire _08450_;
 wire _08451_;
 wire _08452_;
 wire _08453_;
 wire _08454_;
 wire _08455_;
 wire _08456_;
 wire _08457_;
 wire _08458_;
 wire _08459_;
 wire _08460_;
 wire _08461_;
 wire _08462_;
 wire _08463_;
 wire _08464_;
 wire _08465_;
 wire _08466_;
 wire _08467_;
 wire _08468_;
 wire _08469_;
 wire _08470_;
 wire _08471_;
 wire _08472_;
 wire _08473_;
 wire _08474_;
 wire _08475_;
 wire _08476_;
 wire _08477_;
 wire _08478_;
 wire _08479_;
 wire _08480_;
 wire _08481_;
 wire _08482_;
 wire _08483_;
 wire _08484_;
 wire _08485_;
 wire _08486_;
 wire _08487_;
 wire _08488_;
 wire _08489_;
 wire _08490_;
 wire _08491_;
 wire _08492_;
 wire _08493_;
 wire _08494_;
 wire _08495_;
 wire _08496_;
 wire _08497_;
 wire _08498_;
 wire _08499_;
 wire _08500_;
 wire _08501_;
 wire _08502_;
 wire _08503_;
 wire _08504_;
 wire _08505_;
 wire _08506_;
 wire _08507_;
 wire _08508_;
 wire _08509_;
 wire _08510_;
 wire _08511_;
 wire _08512_;
 wire _08513_;
 wire _08514_;
 wire _08515_;
 wire _08516_;
 wire _08517_;
 wire _08518_;
 wire _08519_;
 wire _08520_;
 wire _08521_;
 wire _08522_;
 wire _08523_;
 wire _08524_;
 wire _08525_;
 wire _08526_;
 wire _08527_;
 wire _08528_;
 wire _08529_;
 wire _08530_;
 wire _08531_;
 wire _08532_;
 wire _08533_;
 wire _08534_;
 wire _08535_;
 wire _08536_;
 wire _08537_;
 wire _08538_;
 wire _08539_;
 wire _08540_;
 wire _08541_;
 wire _08542_;
 wire _08543_;
 wire _08544_;
 wire _08545_;
 wire _08546_;
 wire _08547_;
 wire _08548_;
 wire _08549_;
 wire _08550_;
 wire _08551_;
 wire _08552_;
 wire _08553_;
 wire _08554_;
 wire _08555_;
 wire _08556_;
 wire _08557_;
 wire _08558_;
 wire _08559_;
 wire _08560_;
 wire _08561_;
 wire _08562_;
 wire _08563_;
 wire _08564_;
 wire _08565_;
 wire _08566_;
 wire _08567_;
 wire _08568_;
 wire _08569_;
 wire _08570_;
 wire _08571_;
 wire _08572_;
 wire _08573_;
 wire _08574_;
 wire _08575_;
 wire _08576_;
 wire _08577_;
 wire _08578_;
 wire _08579_;
 wire _08580_;
 wire _08581_;
 wire _08582_;
 wire _08583_;
 wire _08584_;
 wire _08585_;
 wire _08586_;
 wire _08587_;
 wire _08588_;
 wire _08589_;
 wire _08590_;
 wire _08591_;
 wire _08592_;
 wire _08593_;
 wire _08594_;
 wire _08595_;
 wire _08596_;
 wire _08597_;
 wire _08598_;
 wire _08599_;
 wire _08600_;
 wire _08601_;
 wire _08602_;
 wire _08603_;
 wire _08604_;
 wire _08605_;
 wire _08606_;
 wire _08607_;
 wire _08608_;
 wire _08609_;
 wire _08610_;
 wire _08611_;
 wire _08612_;
 wire _08613_;
 wire _08614_;
 wire _08615_;
 wire _08616_;
 wire _08617_;
 wire _08618_;
 wire _08619_;
 wire _08620_;
 wire _08621_;
 wire _08622_;
 wire _08623_;
 wire _08624_;
 wire _08625_;
 wire _08626_;
 wire _08627_;
 wire _08628_;
 wire _08629_;
 wire _08630_;
 wire _08631_;
 wire _08632_;
 wire _08633_;
 wire _08634_;
 wire _08635_;
 wire _08636_;
 wire _08637_;
 wire _08638_;
 wire _08639_;
 wire _08640_;
 wire _08641_;
 wire _08642_;
 wire _08643_;
 wire _08644_;
 wire _08645_;
 wire _08646_;
 wire _08647_;
 wire _08648_;
 wire _08649_;
 wire _08650_;
 wire _08651_;
 wire _08652_;
 wire _08653_;
 wire _08654_;
 wire _08655_;
 wire _08656_;
 wire _08657_;
 wire _08658_;
 wire _08659_;
 wire _08660_;
 wire _08661_;
 wire _08662_;
 wire _08663_;
 wire _08664_;
 wire _08665_;
 wire _08666_;
 wire _08667_;
 wire _08668_;
 wire _08669_;
 wire _08670_;
 wire _08671_;
 wire _08672_;
 wire _08673_;
 wire _08674_;
 wire _08675_;
 wire _08676_;
 wire _08677_;
 wire _08678_;
 wire _08679_;
 wire _08680_;
 wire _08681_;
 wire _08682_;
 wire _08683_;
 wire _08684_;
 wire _08685_;
 wire _08686_;
 wire _08687_;
 wire _08688_;
 wire _08689_;
 wire _08690_;
 wire _08691_;
 wire _08692_;
 wire _08693_;
 wire _08694_;
 wire _08695_;
 wire _08696_;
 wire _08697_;
 wire _08698_;
 wire _08699_;
 wire _08700_;
 wire _08701_;
 wire _08702_;
 wire _08703_;
 wire _08704_;
 wire _08705_;
 wire _08706_;
 wire _08707_;
 wire _08708_;
 wire _08709_;
 wire _08710_;
 wire _08711_;
 wire _08712_;
 wire _08713_;
 wire _08714_;
 wire _08715_;
 wire _08716_;
 wire _08717_;
 wire _08718_;
 wire _08719_;
 wire _08720_;
 wire _08721_;
 wire _08722_;
 wire _08723_;
 wire _08724_;
 wire _08725_;
 wire _08726_;
 wire _08727_;
 wire _08728_;
 wire _08729_;
 wire _08730_;
 wire _08731_;
 wire _08732_;
 wire _08733_;
 wire _08734_;
 wire _08735_;
 wire _08736_;
 wire _08737_;
 wire _08738_;
 wire _08739_;
 wire _08740_;
 wire _08741_;
 wire _08742_;
 wire _08743_;
 wire _08744_;
 wire _08745_;
 wire _08746_;
 wire _08747_;
 wire _08748_;
 wire _08749_;
 wire _08750_;
 wire _08751_;
 wire _08752_;
 wire _08753_;
 wire _08754_;
 wire _08755_;
 wire _08756_;
 wire _08757_;
 wire _08758_;
 wire _08759_;
 wire _08760_;
 wire _08761_;
 wire _08762_;
 wire _08763_;
 wire _08764_;
 wire _08765_;
 wire _08766_;
 wire _08767_;
 wire _08768_;
 wire _08769_;
 wire _08770_;
 wire _08771_;
 wire _08772_;
 wire _08773_;
 wire _08774_;
 wire _08775_;
 wire _08776_;
 wire _08777_;
 wire _08778_;
 wire _08779_;
 wire _08780_;
 wire _08781_;
 wire _08782_;
 wire _08783_;
 wire _08784_;
 wire _08785_;
 wire _08786_;
 wire _08787_;
 wire _08788_;
 wire _08789_;
 wire _08790_;
 wire _08791_;
 wire _08792_;
 wire _08793_;
 wire _08794_;
 wire _08795_;
 wire _08796_;
 wire _08797_;
 wire _08798_;
 wire _08799_;
 wire _08800_;
 wire _08801_;
 wire _08802_;
 wire _08803_;
 wire _08804_;
 wire _08805_;
 wire _08806_;
 wire _08807_;
 wire _08808_;
 wire _08809_;
 wire _08810_;
 wire _08811_;
 wire _08812_;
 wire _08813_;
 wire _08814_;
 wire _08815_;
 wire _08816_;
 wire _08817_;
 wire _08818_;
 wire _08819_;
 wire _08820_;
 wire _08821_;
 wire _08822_;
 wire _08823_;
 wire _08824_;
 wire _08825_;
 wire _08826_;
 wire _08827_;
 wire _08828_;
 wire _08829_;
 wire _08830_;
 wire _08831_;
 wire _08832_;
 wire _08833_;
 wire _08834_;
 wire _08835_;
 wire _08836_;
 wire _08837_;
 wire _08838_;
 wire _08839_;
 wire _08840_;
 wire _08841_;
 wire _08842_;
 wire _08843_;
 wire _08844_;
 wire _08845_;
 wire _08846_;
 wire _08847_;
 wire _08848_;
 wire _08849_;
 wire _08850_;
 wire _08851_;
 wire _08852_;
 wire _08853_;
 wire _08854_;
 wire _08855_;
 wire _08856_;
 wire _08857_;
 wire _08858_;
 wire _08859_;
 wire _08860_;
 wire _08861_;
 wire _08862_;
 wire _08863_;
 wire _08864_;
 wire _08865_;
 wire _08866_;
 wire _08867_;
 wire _08868_;
 wire _08869_;
 wire _08870_;
 wire _08871_;
 wire _08872_;
 wire _08873_;
 wire _08874_;
 wire _08875_;
 wire _08876_;
 wire _08877_;
 wire _08878_;
 wire _08879_;
 wire _08880_;
 wire _08881_;
 wire _08882_;
 wire _08883_;
 wire _08884_;
 wire _08885_;
 wire _08886_;
 wire _08887_;
 wire _08888_;
 wire _08889_;
 wire _08890_;
 wire _08891_;
 wire _08892_;
 wire _08893_;
 wire _08894_;
 wire _08895_;
 wire _08896_;
 wire _08897_;
 wire _08898_;
 wire _08899_;
 wire _08900_;
 wire _08901_;
 wire _08902_;
 wire _08903_;
 wire _08904_;
 wire _08905_;
 wire _08906_;
 wire _08907_;
 wire _08908_;
 wire _08909_;
 wire _08910_;
 wire _08911_;
 wire _08912_;
 wire _08913_;
 wire _08914_;
 wire _08915_;
 wire _08916_;
 wire _08917_;
 wire _08918_;
 wire _08919_;
 wire _08920_;
 wire _08921_;
 wire _08922_;
 wire _08923_;
 wire _08924_;
 wire _08925_;
 wire _08926_;
 wire _08927_;
 wire _08928_;
 wire _08929_;
 wire _08930_;
 wire _08931_;
 wire _08932_;
 wire _08933_;
 wire _08934_;
 wire _08935_;
 wire _08936_;
 wire _08937_;
 wire _08938_;
 wire _08939_;
 wire _08940_;
 wire _08941_;
 wire _08942_;
 wire _08943_;
 wire _08944_;
 wire _08945_;
 wire _08946_;
 wire _08947_;
 wire _08948_;
 wire _08949_;
 wire _08950_;
 wire _08951_;
 wire _08952_;
 wire _08953_;
 wire _08954_;
 wire _08955_;
 wire _08956_;
 wire _08957_;
 wire _08958_;
 wire _08959_;
 wire _08960_;
 wire _08961_;
 wire _08962_;
 wire _08963_;
 wire _08964_;
 wire _08965_;
 wire _08966_;
 wire _08967_;
 wire _08968_;
 wire _08969_;
 wire _08970_;
 wire _08971_;
 wire _08972_;
 wire _08973_;
 wire _08974_;
 wire _08975_;
 wire _08976_;
 wire _08977_;
 wire _08978_;
 wire _08979_;
 wire _08980_;
 wire _08981_;
 wire _08982_;
 wire _08983_;
 wire _08984_;
 wire _08985_;
 wire _08986_;
 wire _08987_;
 wire _08988_;
 wire _08989_;
 wire _08990_;
 wire _08991_;
 wire _08992_;
 wire _08993_;
 wire _08994_;
 wire _08995_;
 wire _08996_;
 wire _08997_;
 wire _08998_;
 wire _08999_;
 wire _09000_;
 wire _09001_;
 wire _09002_;
 wire _09003_;
 wire _09004_;
 wire _09005_;
 wire _09006_;
 wire _09007_;
 wire _09008_;
 wire _09009_;
 wire _09010_;
 wire _09011_;
 wire _09012_;
 wire _09013_;
 wire _09014_;
 wire _09015_;
 wire _09016_;
 wire _09017_;
 wire _09018_;
 wire _09019_;
 wire _09020_;
 wire _09021_;
 wire _09022_;
 wire _09023_;
 wire _09024_;
 wire _09025_;
 wire _09026_;
 wire _09027_;
 wire _09028_;
 wire _09029_;
 wire _09030_;
 wire _09031_;
 wire _09032_;
 wire _09033_;
 wire _09034_;
 wire _09035_;
 wire _09036_;
 wire _09037_;
 wire _09038_;
 wire _09039_;
 wire _09040_;
 wire _09041_;
 wire _09042_;
 wire _09043_;
 wire _09044_;
 wire _09045_;
 wire _09046_;
 wire _09047_;
 wire _09048_;
 wire _09049_;
 wire _09050_;
 wire _09051_;
 wire _09052_;
 wire _09053_;
 wire _09054_;
 wire _09055_;
 wire _09056_;
 wire _09057_;
 wire _09058_;
 wire _09059_;
 wire _09060_;
 wire _09061_;
 wire _09062_;
 wire _09063_;
 wire _09064_;
 wire _09065_;
 wire _09066_;
 wire _09067_;
 wire _09068_;
 wire _09069_;
 wire _09070_;
 wire _09071_;
 wire _09072_;
 wire _09073_;
 wire _09074_;
 wire _09075_;
 wire _09076_;
 wire _09077_;
 wire _09078_;
 wire _09079_;
 wire _09080_;
 wire _09081_;
 wire _09082_;
 wire _09083_;
 wire _09084_;
 wire _09085_;
 wire _09086_;
 wire _09087_;
 wire _09088_;
 wire _09089_;
 wire _09090_;
 wire _09091_;
 wire _09092_;
 wire _09093_;
 wire _09094_;
 wire _09095_;
 wire _09096_;
 wire _09097_;
 wire _09098_;
 wire _09099_;
 wire _09100_;
 wire _09101_;
 wire _09102_;
 wire _09103_;
 wire _09104_;
 wire _09105_;
 wire _09106_;
 wire _09107_;
 wire _09108_;
 wire _09109_;
 wire _09110_;
 wire _09111_;
 wire _09112_;
 wire _09113_;
 wire _09114_;
 wire _09115_;
 wire _09116_;
 wire _09117_;
 wire _09118_;
 wire _09119_;
 wire _09120_;
 wire _09121_;
 wire _09122_;
 wire _09123_;
 wire _09124_;
 wire _09125_;
 wire _09126_;
 wire _09127_;
 wire _09128_;
 wire _09129_;
 wire _09130_;
 wire _09131_;
 wire _09132_;
 wire _09133_;
 wire _09134_;
 wire _09135_;
 wire _09136_;
 wire _09137_;
 wire _09138_;
 wire _09139_;
 wire _09140_;
 wire _09141_;
 wire _09142_;
 wire _09143_;
 wire _09144_;
 wire _09145_;
 wire _09146_;
 wire _09147_;
 wire _09148_;
 wire _09149_;
 wire _09150_;
 wire _09151_;
 wire _09152_;
 wire _09153_;
 wire _09154_;
 wire _09155_;
 wire _09156_;
 wire _09157_;
 wire _09158_;
 wire _09159_;
 wire _09160_;
 wire _09161_;
 wire _09162_;
 wire _09163_;
 wire _09164_;
 wire _09165_;
 wire _09166_;
 wire _09167_;
 wire _09168_;
 wire _09169_;
 wire _09170_;
 wire _09171_;
 wire _09172_;
 wire _09173_;
 wire _09174_;
 wire _09175_;
 wire _09176_;
 wire _09177_;
 wire _09178_;
 wire _09179_;
 wire _09180_;
 wire _09181_;
 wire _09182_;
 wire _09183_;
 wire _09184_;
 wire _09185_;
 wire _09186_;
 wire _09187_;
 wire _09188_;
 wire _09189_;
 wire _09190_;
 wire _09191_;
 wire _09192_;
 wire _09193_;
 wire _09194_;
 wire _09195_;
 wire _09196_;
 wire _09197_;
 wire _09198_;
 wire _09199_;
 wire _09200_;
 wire _09201_;
 wire _09202_;
 wire _09203_;
 wire _09204_;
 wire _09205_;
 wire _09206_;
 wire _09207_;
 wire _09208_;
 wire _09209_;
 wire _09210_;
 wire _09211_;
 wire _09212_;
 wire _09213_;
 wire _09214_;
 wire _09215_;
 wire _09216_;
 wire _09217_;
 wire _09218_;
 wire _09219_;
 wire _09220_;
 wire _09221_;
 wire _09222_;
 wire _09223_;
 wire _09224_;
 wire _09225_;
 wire _09226_;
 wire _09227_;
 wire _09228_;
 wire _09229_;
 wire _09230_;
 wire _09231_;
 wire _09232_;
 wire _09233_;
 wire _09234_;
 wire _09235_;
 wire _09236_;
 wire _09237_;
 wire _09238_;
 wire _09239_;
 wire _09240_;
 wire _09241_;
 wire _09242_;
 wire _09243_;
 wire _09244_;
 wire _09245_;
 wire _09246_;
 wire _09247_;
 wire _09248_;
 wire _09249_;
 wire _09250_;
 wire _09251_;
 wire _09252_;
 wire _09253_;
 wire _09254_;
 wire _09255_;
 wire _09256_;
 wire _09257_;
 wire _09258_;
 wire _09259_;
 wire _09260_;
 wire _09261_;
 wire _09262_;
 wire _09263_;
 wire _09264_;
 wire _09265_;
 wire _09266_;
 wire _09267_;
 wire _09268_;
 wire _09269_;
 wire _09270_;
 wire _09271_;
 wire _09272_;
 wire _09273_;
 wire _09274_;
 wire _09275_;
 wire _09276_;
 wire _09277_;
 wire _09278_;
 wire _09279_;
 wire _09280_;
 wire _09281_;
 wire _09282_;
 wire _09283_;
 wire _09284_;
 wire _09285_;
 wire _09286_;
 wire _09287_;
 wire _09288_;
 wire _09289_;
 wire _09290_;
 wire _09291_;
 wire _09292_;
 wire _09293_;
 wire _09294_;
 wire _09295_;
 wire _09296_;
 wire _09297_;
 wire _09298_;
 wire _09299_;
 wire _09300_;
 wire _09301_;
 wire _09302_;
 wire _09303_;
 wire _09304_;
 wire _09305_;
 wire _09306_;
 wire _09307_;
 wire _09308_;
 wire _09309_;
 wire _09310_;
 wire _09311_;
 wire _09312_;
 wire _09313_;
 wire _09314_;
 wire _09315_;
 wire _09316_;
 wire _09317_;
 wire _09318_;
 wire _09319_;
 wire _09320_;
 wire _09321_;
 wire _09322_;
 wire _09323_;
 wire _09324_;
 wire _09325_;
 wire _09326_;
 wire _09327_;
 wire _09328_;
 wire _09329_;
 wire _09330_;
 wire _09331_;
 wire _09332_;
 wire _09333_;
 wire _09334_;
 wire _09335_;
 wire _09336_;
 wire _09337_;
 wire _09338_;
 wire _09339_;
 wire _09340_;
 wire _09341_;
 wire _09342_;
 wire _09343_;
 wire _09344_;
 wire _09345_;
 wire _09346_;
 wire _09347_;
 wire _09348_;
 wire _09349_;
 wire _09350_;
 wire _09351_;
 wire _09352_;
 wire _09353_;
 wire _09354_;
 wire _09355_;
 wire _09356_;
 wire _09357_;
 wire _09358_;
 wire _09359_;
 wire _09360_;
 wire _09361_;
 wire _09362_;
 wire _09363_;
 wire _09364_;
 wire _09365_;
 wire _09366_;
 wire _09367_;
 wire _09368_;
 wire _09369_;
 wire _09370_;
 wire _09371_;
 wire _09372_;
 wire _09373_;
 wire _09374_;
 wire _09375_;
 wire _09376_;
 wire _09377_;
 wire _09378_;
 wire _09379_;
 wire _09380_;
 wire _09381_;
 wire _09382_;
 wire _09383_;
 wire _09384_;
 wire _09385_;
 wire _09386_;
 wire _09387_;
 wire _09388_;
 wire _09389_;
 wire _09390_;
 wire _09391_;
 wire _09392_;
 wire _09393_;
 wire _09394_;
 wire _09395_;
 wire _09396_;
 wire _09397_;
 wire _09398_;
 wire _09399_;
 wire _09400_;
 wire _09401_;
 wire _09402_;
 wire _09403_;
 wire _09404_;
 wire _09405_;
 wire _09406_;
 wire _09407_;
 wire _09408_;
 wire _09409_;
 wire _09410_;
 wire _09411_;
 wire _09412_;
 wire _09413_;
 wire _09414_;
 wire _09415_;
 wire _09416_;
 wire _09417_;
 wire _09418_;
 wire _09419_;
 wire _09420_;
 wire _09421_;
 wire _09422_;
 wire _09423_;
 wire _09424_;
 wire _09425_;
 wire _09426_;
 wire _09427_;
 wire _09428_;
 wire _09429_;
 wire _09430_;
 wire _09431_;
 wire _09432_;
 wire _09433_;
 wire _09434_;
 wire _09435_;
 wire _09436_;
 wire _09437_;
 wire _09438_;
 wire _09439_;
 wire _09440_;
 wire _09441_;
 wire _09442_;
 wire _09443_;
 wire _09444_;
 wire _09445_;
 wire _09446_;
 wire _09447_;
 wire _09448_;
 wire _09449_;
 wire _09450_;
 wire _09451_;
 wire _09452_;
 wire _09453_;
 wire _09454_;
 wire _09455_;
 wire _09456_;
 wire _09457_;
 wire _09458_;
 wire _09459_;
 wire _09460_;
 wire _09461_;
 wire _09462_;
 wire _09463_;
 wire _09464_;
 wire _09465_;
 wire _09466_;
 wire _09467_;
 wire _09468_;
 wire _09469_;
 wire _09470_;
 wire _09471_;
 wire _09472_;
 wire _09473_;
 wire _09474_;
 wire _09475_;
 wire _09476_;
 wire _09477_;
 wire _09478_;
 wire _09479_;
 wire _09480_;
 wire _09481_;
 wire _09482_;
 wire _09483_;
 wire _09484_;
 wire _09485_;
 wire _09486_;
 wire _09487_;
 wire _09488_;
 wire _09489_;
 wire _09490_;
 wire _09491_;
 wire _09492_;
 wire _09493_;
 wire _09494_;
 wire _09495_;
 wire _09496_;
 wire _09497_;
 wire _09498_;
 wire _09499_;
 wire _09500_;
 wire _09501_;
 wire _09502_;
 wire _09503_;
 wire _09504_;
 wire _09505_;
 wire _09506_;
 wire _09507_;
 wire _09508_;
 wire _09509_;
 wire _09510_;
 wire _09511_;
 wire _09512_;
 wire _09513_;
 wire _09514_;
 wire _09515_;
 wire _09516_;
 wire _09517_;
 wire _09518_;
 wire _09519_;
 wire _09520_;
 wire _09521_;
 wire _09522_;
 wire _09523_;
 wire _09524_;
 wire _09525_;
 wire _09526_;
 wire _09527_;
 wire _09528_;
 wire _09529_;
 wire _09530_;
 wire _09531_;
 wire _09532_;
 wire _09533_;
 wire _09534_;
 wire _09535_;
 wire _09536_;
 wire _09537_;
 wire _09538_;
 wire _09539_;
 wire _09540_;
 wire _09541_;
 wire _09542_;
 wire _09543_;
 wire _09544_;
 wire _09545_;
 wire _09546_;
 wire _09547_;
 wire _09548_;
 wire _09549_;
 wire _09550_;
 wire _09551_;
 wire _09552_;
 wire _09553_;
 wire _09554_;
 wire _09555_;
 wire _09556_;
 wire _09557_;
 wire _09558_;
 wire _09559_;
 wire _09560_;
 wire _09561_;
 wire _09562_;
 wire _09563_;
 wire _09564_;
 wire _09565_;
 wire _09566_;
 wire _09567_;
 wire _09568_;
 wire _09569_;
 wire _09570_;
 wire _09571_;
 wire _09572_;
 wire _09573_;
 wire _09574_;
 wire _09575_;
 wire _09576_;
 wire _09577_;
 wire _09578_;
 wire _09579_;
 wire _09580_;
 wire _09581_;
 wire _09582_;
 wire _09583_;
 wire _09584_;
 wire _09585_;
 wire _09586_;
 wire _09587_;
 wire _09588_;
 wire _09589_;
 wire _09590_;
 wire _09591_;
 wire _09592_;
 wire _09593_;
 wire _09594_;
 wire _09595_;
 wire _09596_;
 wire _09597_;
 wire _09598_;
 wire _09599_;
 wire _09600_;
 wire _09601_;
 wire _09602_;
 wire _09603_;
 wire _09604_;
 wire _09605_;
 wire _09606_;
 wire _09607_;
 wire _09608_;
 wire _09609_;
 wire _09610_;
 wire _09611_;
 wire _09612_;
 wire _09613_;
 wire _09614_;
 wire _09615_;
 wire _09616_;
 wire _09617_;
 wire _09618_;
 wire _09619_;
 wire _09620_;
 wire _09621_;
 wire _09622_;
 wire _09623_;
 wire _09624_;
 wire _09625_;
 wire _09626_;
 wire _09627_;
 wire _09628_;
 wire _09629_;
 wire _09630_;
 wire _09631_;
 wire _09632_;
 wire _09633_;
 wire _09634_;
 wire _09635_;
 wire _09636_;
 wire _09637_;
 wire _09638_;
 wire _09639_;
 wire _09640_;
 wire _09641_;
 wire _09642_;
 wire _09643_;
 wire _09644_;
 wire _09645_;
 wire _09646_;
 wire _09647_;
 wire _09648_;
 wire _09649_;
 wire _09650_;
 wire _09651_;
 wire _09652_;
 wire _09653_;
 wire _09654_;
 wire _09655_;
 wire _09656_;
 wire _09657_;
 wire _09658_;
 wire _09659_;
 wire _09660_;
 wire _09661_;
 wire _09662_;
 wire _09663_;
 wire _09664_;
 wire _09665_;
 wire _09666_;
 wire _09667_;
 wire _09668_;
 wire _09669_;
 wire _09670_;
 wire _09671_;
 wire _09672_;
 wire _09673_;
 wire _09674_;
 wire _09675_;
 wire _09676_;
 wire _09677_;
 wire _09678_;
 wire _09679_;
 wire _09680_;
 wire _09681_;
 wire _09682_;
 wire _09683_;
 wire _09684_;
 wire _09685_;
 wire _09686_;
 wire _09687_;
 wire _09688_;
 wire _09689_;
 wire _09690_;
 wire _09691_;
 wire _09692_;
 wire _09693_;
 wire _09694_;
 wire _09695_;
 wire _09696_;
 wire _09697_;
 wire _09698_;
 wire _09699_;
 wire _09700_;
 wire _09701_;
 wire _09702_;
 wire _09703_;
 wire _09704_;
 wire _09705_;
 wire _09706_;
 wire _09707_;
 wire _09708_;
 wire _09709_;
 wire _09710_;
 wire _09711_;
 wire _09712_;
 wire _09713_;
 wire _09714_;
 wire _09715_;
 wire _09716_;
 wire _09717_;
 wire _09718_;
 wire _09719_;
 wire _09720_;
 wire _09721_;
 wire _09722_;
 wire _09723_;
 wire _09724_;
 wire _09725_;
 wire _09726_;
 wire _09727_;
 wire _09728_;
 wire _09729_;
 wire _09730_;
 wire _09731_;
 wire _09732_;
 wire _09733_;
 wire _09734_;
 wire _09735_;
 wire _09736_;
 wire _09737_;
 wire _09738_;
 wire _09739_;
 wire _09740_;
 wire _09741_;
 wire _09742_;
 wire _09743_;
 wire _09744_;
 wire _09745_;
 wire _09746_;
 wire _09747_;
 wire _09748_;
 wire _09749_;
 wire _09750_;
 wire _09751_;
 wire _09752_;
 wire _09753_;
 wire _09754_;
 wire _09755_;
 wire _09756_;
 wire _09757_;
 wire _09758_;
 wire _09759_;
 wire _09760_;
 wire _09761_;
 wire _09762_;
 wire _09763_;
 wire _09764_;
 wire _09765_;
 wire _09766_;
 wire _09767_;
 wire _09768_;
 wire _09769_;
 wire _09770_;
 wire _09771_;
 wire _09772_;
 wire _09773_;
 wire _09774_;
 wire _09775_;
 wire _09776_;
 wire _09777_;
 wire _09778_;
 wire _09779_;
 wire _09780_;
 wire _09781_;
 wire _09782_;
 wire _09783_;
 wire _09784_;
 wire _09785_;
 wire _09786_;
 wire _09787_;
 wire _09788_;
 wire _09789_;
 wire _09790_;
 wire _09791_;
 wire _09792_;
 wire _09793_;
 wire _09794_;
 wire _09795_;
 wire _09796_;
 wire _09797_;
 wire _09798_;
 wire _09799_;
 wire _09800_;
 wire _09801_;
 wire _09802_;
 wire _09803_;
 wire _09804_;
 wire _09805_;
 wire _09806_;
 wire _09807_;
 wire _09808_;
 wire _09809_;
 wire _09810_;
 wire _09811_;
 wire _09812_;
 wire _09813_;
 wire _09814_;
 wire _09815_;
 wire _09816_;
 wire _09817_;
 wire _09818_;
 wire _09819_;
 wire _09820_;
 wire _09821_;
 wire _09822_;
 wire _09823_;
 wire _09824_;
 wire _09825_;
 wire _09826_;
 wire _09827_;
 wire _09828_;
 wire _09829_;
 wire _09830_;
 wire _09831_;
 wire _09832_;
 wire _09833_;
 wire _09834_;
 wire _09835_;
 wire _09836_;
 wire _09837_;
 wire _09838_;
 wire _09839_;
 wire _09840_;
 wire _09841_;
 wire _09842_;
 wire _09843_;
 wire _09844_;
 wire _09845_;
 wire _09846_;
 wire _09847_;
 wire _09848_;
 wire _09849_;
 wire _09850_;
 wire _09851_;
 wire _09852_;
 wire _09853_;
 wire _09854_;
 wire _09855_;
 wire _09856_;
 wire _09857_;
 wire _09858_;
 wire _09859_;
 wire _09860_;
 wire _09861_;
 wire _09862_;
 wire _09863_;
 wire _09864_;
 wire _09865_;
 wire _09866_;
 wire _09867_;
 wire _09868_;
 wire _09869_;
 wire _09870_;
 wire _09871_;
 wire _09872_;
 wire _09873_;
 wire _09874_;
 wire _09875_;
 wire _09876_;
 wire _09877_;
 wire _09878_;
 wire _09879_;
 wire _09880_;
 wire _09881_;
 wire _09882_;
 wire _09883_;
 wire _09884_;
 wire _09885_;
 wire _09886_;
 wire _09887_;
 wire _09888_;
 wire _09889_;
 wire _09890_;
 wire _09891_;
 wire _09892_;
 wire _09893_;
 wire _09894_;
 wire _09895_;
 wire _09896_;
 wire _09897_;
 wire _09898_;
 wire _09899_;
 wire _09900_;
 wire _09901_;
 wire _09902_;
 wire _09903_;
 wire _09904_;
 wire _09905_;
 wire _09906_;
 wire _09907_;
 wire _09908_;
 wire _09909_;
 wire _09910_;
 wire _09911_;
 wire _09912_;
 wire _09913_;
 wire _09914_;
 wire _09915_;
 wire _09916_;
 wire _09917_;
 wire _09918_;
 wire _09919_;
 wire _09920_;
 wire _09921_;
 wire _09922_;
 wire _09923_;
 wire _09924_;
 wire _09925_;
 wire _09926_;
 wire _09927_;
 wire _09928_;
 wire _09929_;
 wire _09930_;
 wire _09931_;
 wire _09932_;
 wire _09933_;
 wire _09934_;
 wire _09935_;
 wire _09936_;
 wire _09937_;
 wire _09938_;
 wire _09939_;
 wire _09940_;
 wire _09941_;
 wire _09942_;
 wire _09943_;
 wire _09944_;
 wire _09945_;
 wire _09946_;
 wire _09947_;
 wire _09948_;
 wire _09949_;
 wire _09950_;
 wire _09951_;
 wire _09952_;
 wire _09953_;
 wire _09954_;
 wire _09955_;
 wire _09956_;
 wire _09957_;
 wire _09958_;
 wire _09959_;
 wire _09960_;
 wire _09961_;
 wire _09962_;
 wire _09963_;
 wire _09964_;
 wire _09965_;
 wire _09966_;
 wire _09967_;
 wire _09968_;
 wire _09969_;
 wire _09970_;
 wire _09971_;
 wire _09972_;
 wire _09973_;
 wire _09974_;
 wire _09975_;
 wire _09976_;
 wire _09977_;
 wire _09978_;
 wire _09979_;
 wire _09980_;
 wire _09981_;
 wire _09982_;
 wire _09983_;
 wire _09984_;
 wire _09985_;
 wire _09986_;
 wire _09987_;
 wire _09988_;
 wire _09989_;
 wire _09990_;
 wire _09991_;
 wire _09992_;
 wire _09993_;
 wire _09994_;
 wire _09995_;
 wire _09996_;
 wire _09997_;
 wire _09998_;
 wire _09999_;
 wire _10000_;
 wire _10001_;
 wire _10002_;
 wire _10003_;
 wire _10004_;
 wire _10005_;
 wire _10006_;
 wire _10007_;
 wire _10008_;
 wire _10009_;
 wire _10010_;
 wire _10011_;
 wire _10012_;
 wire _10013_;
 wire _10014_;
 wire _10015_;
 wire _10016_;
 wire _10017_;
 wire _10018_;
 wire _10019_;
 wire _10020_;
 wire _10021_;
 wire _10022_;
 wire _10023_;
 wire _10024_;
 wire _10025_;
 wire _10026_;
 wire _10027_;
 wire _10028_;
 wire _10029_;
 wire _10030_;
 wire _10031_;
 wire _10032_;
 wire _10033_;
 wire _10034_;
 wire _10035_;
 wire _10036_;
 wire _10037_;
 wire _10038_;
 wire _10039_;
 wire _10040_;
 wire _10041_;
 wire _10042_;
 wire _10043_;
 wire _10044_;
 wire _10045_;
 wire _10046_;
 wire _10047_;
 wire _10048_;
 wire _10049_;
 wire _10050_;
 wire _10051_;
 wire _10052_;
 wire _10053_;
 wire _10054_;
 wire _10055_;
 wire _10056_;
 wire _10057_;
 wire _10058_;
 wire _10059_;
 wire _10060_;
 wire _10061_;
 wire _10062_;
 wire _10063_;
 wire _10064_;
 wire _10065_;
 wire _10066_;
 wire _10067_;
 wire _10068_;
 wire _10069_;
 wire _10070_;
 wire _10071_;
 wire _10072_;
 wire _10073_;
 wire _10074_;
 wire _10075_;
 wire _10076_;
 wire _10077_;
 wire _10078_;
 wire _10079_;
 wire _10080_;
 wire _10081_;
 wire _10082_;
 wire _10083_;
 wire _10084_;
 wire _10085_;
 wire _10086_;
 wire _10087_;
 wire _10088_;
 wire _10089_;
 wire _10090_;
 wire _10091_;
 wire _10092_;
 wire _10093_;
 wire _10094_;
 wire _10095_;
 wire _10096_;
 wire _10097_;
 wire _10098_;
 wire _10099_;
 wire _10100_;
 wire _10101_;
 wire _10102_;
 wire _10103_;
 wire _10104_;
 wire _10105_;
 wire _10106_;
 wire _10107_;
 wire _10108_;
 wire _10109_;
 wire _10110_;
 wire _10111_;
 wire _10112_;
 wire _10113_;
 wire _10114_;
 wire _10115_;
 wire _10116_;
 wire _10117_;
 wire _10118_;
 wire _10119_;
 wire _10120_;
 wire _10121_;
 wire _10122_;
 wire _10123_;
 wire _10124_;
 wire _10125_;
 wire _10126_;
 wire _10127_;
 wire _10128_;
 wire _10129_;
 wire _10130_;
 wire _10131_;
 wire _10132_;
 wire _10133_;
 wire _10134_;
 wire _10135_;
 wire _10136_;
 wire _10137_;
 wire _10138_;
 wire _10139_;
 wire _10140_;
 wire _10141_;
 wire _10142_;
 wire _10143_;
 wire _10144_;
 wire _10145_;
 wire _10146_;
 wire _10147_;
 wire _10148_;
 wire _10149_;
 wire _10150_;
 wire _10151_;
 wire _10152_;
 wire _10153_;
 wire _10154_;
 wire _10155_;
 wire _10156_;
 wire _10157_;
 wire _10158_;
 wire _10159_;
 wire _10160_;
 wire _10161_;
 wire _10162_;
 wire _10163_;
 wire _10164_;
 wire _10165_;
 wire _10166_;
 wire _10167_;
 wire _10168_;
 wire _10169_;
 wire _10170_;
 wire _10171_;
 wire _10172_;
 wire _10173_;
 wire _10174_;
 wire _10175_;
 wire _10176_;
 wire _10177_;
 wire _10178_;
 wire _10179_;
 wire _10180_;
 wire _10181_;
 wire _10182_;
 wire _10183_;
 wire _10184_;
 wire _10185_;
 wire _10186_;
 wire _10187_;
 wire _10188_;
 wire _10189_;
 wire _10190_;
 wire _10191_;
 wire _10192_;
 wire _10193_;
 wire _10194_;
 wire _10195_;
 wire _10196_;
 wire _10197_;
 wire _10198_;
 wire _10199_;
 wire _10200_;
 wire _10201_;
 wire _10202_;
 wire _10203_;
 wire _10204_;
 wire _10205_;
 wire _10206_;
 wire _10207_;
 wire _10208_;
 wire _10209_;
 wire _10210_;
 wire _10211_;
 wire _10212_;
 wire _10213_;
 wire _10214_;
 wire _10215_;
 wire _10216_;
 wire _10217_;
 wire _10218_;
 wire _10219_;
 wire _10220_;
 wire _10221_;
 wire _10222_;
 wire _10223_;
 wire _10224_;
 wire _10225_;
 wire _10226_;
 wire _10227_;
 wire _10228_;
 wire _10229_;
 wire _10230_;
 wire _10231_;
 wire _10232_;
 wire _10233_;
 wire _10234_;
 wire _10235_;
 wire _10236_;
 wire _10237_;
 wire _10238_;
 wire _10239_;
 wire _10240_;
 wire _10241_;
 wire _10242_;
 wire _10243_;
 wire _10244_;
 wire _10245_;
 wire _10246_;
 wire _10247_;
 wire _10248_;
 wire _10249_;
 wire _10250_;
 wire _10251_;
 wire _10252_;
 wire _10253_;
 wire _10254_;
 wire _10255_;
 wire _10256_;
 wire _10257_;
 wire _10258_;
 wire _10259_;
 wire _10260_;
 wire _10261_;
 wire _10262_;
 wire _10263_;
 wire _10264_;
 wire _10265_;
 wire _10266_;
 wire _10267_;
 wire _10268_;
 wire _10269_;
 wire _10270_;
 wire _10271_;
 wire _10272_;
 wire _10273_;
 wire _10274_;
 wire _10275_;
 wire _10276_;
 wire _10277_;
 wire _10278_;
 wire _10279_;
 wire _10280_;
 wire _10281_;
 wire _10282_;
 wire _10283_;
 wire _10284_;
 wire _10285_;
 wire _10286_;
 wire _10287_;
 wire _10288_;
 wire _10289_;
 wire _10290_;
 wire _10291_;
 wire _10292_;
 wire _10293_;
 wire _10294_;
 wire _10295_;
 wire _10296_;
 wire _10297_;
 wire _10298_;
 wire _10299_;
 wire _10300_;
 wire _10301_;
 wire _10302_;
 wire _10303_;
 wire _10304_;
 wire _10305_;
 wire _10306_;
 wire _10307_;
 wire _10308_;
 wire _10309_;
 wire _10310_;
 wire _10311_;
 wire _10312_;
 wire _10313_;
 wire _10314_;
 wire _10315_;
 wire _10316_;
 wire _10317_;
 wire _10318_;
 wire _10319_;
 wire _10320_;
 wire _10321_;
 wire _10322_;
 wire _10323_;
 wire _10324_;
 wire _10325_;
 wire _10326_;
 wire _10327_;
 wire _10328_;
 wire _10329_;
 wire _10330_;
 wire _10331_;
 wire _10332_;
 wire _10333_;
 wire _10334_;
 wire _10335_;
 wire _10336_;
 wire _10337_;
 wire _10338_;
 wire _10339_;
 wire _10340_;
 wire _10341_;
 wire _10342_;
 wire _10343_;
 wire _10344_;
 wire _10345_;
 wire _10346_;
 wire _10347_;
 wire _10348_;
 wire _10349_;
 wire _10350_;
 wire _10351_;
 wire _10352_;
 wire _10353_;
 wire _10354_;
 wire _10355_;
 wire _10356_;
 wire _10357_;
 wire _10358_;
 wire _10359_;
 wire _10360_;
 wire _10361_;
 wire _10362_;
 wire _10363_;
 wire _10364_;
 wire _10365_;
 wire _10366_;
 wire _10367_;
 wire _10368_;
 wire _10369_;
 wire _10370_;
 wire _10371_;
 wire _10372_;
 wire _10373_;
 wire _10374_;
 wire _10375_;
 wire _10376_;
 wire _10377_;
 wire _10378_;
 wire _10379_;
 wire _10380_;
 wire _10381_;
 wire _10382_;
 wire _10383_;
 wire _10384_;
 wire _10385_;
 wire _10386_;
 wire _10387_;
 wire _10388_;
 wire _10389_;
 wire _10390_;
 wire _10391_;
 wire _10392_;
 wire _10393_;
 wire _10394_;
 wire _10395_;
 wire _10396_;
 wire _10397_;
 wire _10398_;
 wire _10399_;
 wire _10400_;
 wire _10401_;
 wire _10402_;
 wire _10403_;
 wire _10404_;
 wire _10405_;
 wire _10406_;
 wire _10407_;
 wire _10408_;
 wire _10409_;
 wire _10410_;
 wire _10411_;
 wire _10412_;
 wire _10413_;
 wire _10414_;
 wire _10415_;
 wire _10416_;
 wire _10417_;
 wire _10418_;
 wire _10419_;
 wire _10420_;
 wire _10421_;
 wire _10422_;
 wire _10423_;
 wire _10424_;
 wire _10425_;
 wire _10426_;
 wire _10427_;
 wire _10428_;
 wire _10429_;
 wire _10430_;
 wire _10431_;
 wire _10432_;
 wire _10433_;
 wire _10434_;
 wire _10435_;
 wire _10436_;
 wire _10437_;
 wire _10438_;
 wire _10439_;
 wire _10440_;
 wire _10441_;
 wire _10442_;
 wire _10443_;
 wire _10444_;
 wire _10445_;
 wire _10446_;
 wire _10447_;
 wire _10448_;
 wire _10449_;
 wire _10450_;
 wire _10451_;
 wire _10452_;
 wire _10453_;
 wire _10454_;
 wire _10455_;
 wire _10456_;
 wire _10457_;
 wire _10458_;
 wire _10459_;
 wire _10460_;
 wire _10461_;
 wire _10462_;
 wire _10463_;
 wire _10464_;
 wire _10465_;
 wire _10466_;
 wire _10467_;
 wire _10468_;
 wire _10469_;
 wire _10470_;
 wire _10471_;
 wire _10472_;
 wire _10473_;
 wire _10474_;
 wire _10475_;
 wire _10476_;
 wire _10477_;
 wire _10478_;
 wire _10479_;
 wire _10480_;
 wire _10481_;
 wire _10482_;
 wire _10483_;
 wire _10484_;
 wire _10485_;
 wire _10486_;
 wire _10487_;
 wire _10488_;
 wire _10489_;
 wire _10490_;
 wire _10491_;
 wire _10492_;
 wire _10493_;
 wire _10494_;
 wire _10495_;
 wire _10496_;
 wire _10497_;
 wire _10498_;
 wire _10499_;
 wire _10500_;
 wire _10501_;
 wire _10502_;
 wire _10503_;
 wire _10504_;
 wire _10505_;
 wire _10506_;
 wire _10507_;
 wire _10508_;
 wire _10509_;
 wire _10510_;
 wire _10511_;
 wire _10512_;
 wire _10513_;
 wire _10514_;
 wire _10515_;
 wire _10516_;
 wire _10517_;
 wire _10518_;
 wire _10519_;
 wire _10520_;
 wire _10521_;
 wire _10522_;
 wire _10523_;
 wire _10524_;
 wire _10525_;
 wire _10526_;
 wire _10527_;
 wire _10528_;
 wire _10529_;
 wire _10530_;
 wire _10531_;
 wire _10532_;
 wire _10533_;
 wire _10534_;
 wire _10535_;
 wire _10536_;
 wire _10537_;
 wire _10538_;
 wire _10539_;
 wire _10540_;
 wire _10541_;
 wire _10542_;
 wire _10543_;
 wire _10544_;
 wire _10545_;
 wire _10546_;
 wire _10547_;
 wire _10548_;
 wire _10549_;
 wire _10550_;
 wire _10551_;
 wire _10552_;
 wire _10553_;
 wire _10554_;
 wire _10555_;
 wire _10556_;
 wire _10557_;
 wire _10558_;
 wire _10559_;
 wire _10560_;
 wire _10561_;
 wire _10562_;
 wire _10563_;
 wire _10564_;
 wire _10565_;
 wire _10566_;
 wire _10567_;
 wire _10568_;
 wire _10569_;
 wire _10570_;
 wire _10571_;
 wire _10572_;
 wire _10573_;
 wire _10574_;
 wire _10575_;
 wire _10576_;
 wire _10577_;
 wire _10578_;
 wire _10579_;
 wire _10580_;
 wire _10581_;
 wire _10582_;
 wire _10583_;
 wire _10584_;
 wire _10585_;
 wire _10586_;
 wire _10587_;
 wire _10588_;
 wire _10589_;
 wire _10590_;
 wire _10591_;
 wire _10592_;
 wire _10593_;
 wire _10594_;
 wire _10595_;
 wire _10596_;
 wire _10597_;
 wire _10598_;
 wire _10599_;
 wire _10600_;
 wire _10601_;
 wire _10602_;
 wire _10603_;
 wire _10604_;
 wire _10605_;
 wire _10606_;
 wire _10607_;
 wire _10608_;
 wire _10609_;
 wire _10610_;
 wire _10611_;
 wire _10612_;
 wire _10613_;
 wire _10614_;
 wire _10615_;
 wire _10616_;
 wire _10617_;
 wire _10618_;
 wire _10619_;
 wire _10620_;
 wire _10621_;
 wire _10622_;
 wire _10623_;
 wire _10624_;
 wire _10625_;
 wire _10626_;
 wire _10627_;
 wire _10628_;
 wire _10629_;
 wire _10630_;
 wire _10631_;
 wire _10632_;
 wire _10633_;
 wire _10634_;
 wire _10635_;
 wire _10636_;
 wire _10637_;
 wire _10638_;
 wire _10639_;
 wire _10640_;
 wire _10641_;
 wire _10642_;
 wire _10643_;
 wire _10644_;
 wire _10645_;
 wire _10646_;
 wire _10647_;
 wire _10648_;
 wire _10649_;
 wire _10650_;
 wire _10651_;
 wire _10652_;
 wire _10653_;
 wire _10654_;
 wire _10655_;
 wire _10656_;
 wire _10657_;
 wire _10658_;
 wire _10659_;
 wire _10660_;
 wire _10661_;
 wire _10662_;
 wire _10663_;
 wire _10664_;
 wire _10665_;
 wire _10666_;
 wire _10667_;
 wire _10668_;
 wire _10669_;
 wire _10670_;
 wire _10671_;
 wire _10672_;
 wire _10673_;
 wire _10674_;
 wire _10675_;
 wire _10676_;
 wire _10677_;
 wire _10678_;
 wire _10679_;
 wire _10680_;
 wire _10681_;
 wire _10682_;
 wire _10683_;
 wire _10684_;
 wire _10685_;
 wire _10686_;
 wire _10687_;
 wire _10688_;
 wire _10689_;
 wire _10690_;
 wire _10691_;
 wire _10692_;
 wire _10693_;
 wire _10694_;
 wire _10695_;
 wire _10696_;
 wire _10697_;
 wire _10698_;
 wire _10699_;
 wire _10700_;
 wire _10701_;
 wire _10702_;
 wire _10703_;
 wire _10704_;
 wire _10705_;
 wire _10706_;
 wire _10707_;
 wire _10708_;
 wire _10709_;
 wire _10710_;
 wire _10711_;
 wire _10712_;
 wire _10713_;
 wire _10714_;
 wire _10715_;
 wire _10716_;
 wire _10717_;
 wire _10718_;
 wire _10719_;
 wire _10720_;
 wire _10721_;
 wire _10722_;
 wire _10723_;
 wire _10724_;
 wire _10725_;
 wire _10726_;
 wire _10727_;
 wire _10728_;
 wire _10729_;
 wire _10730_;
 wire _10731_;
 wire _10732_;
 wire _10733_;
 wire _10734_;
 wire _10735_;
 wire _10736_;
 wire _10737_;
 wire _10738_;
 wire _10739_;
 wire _10740_;
 wire _10741_;
 wire _10742_;
 wire _10743_;
 wire _10744_;
 wire _10745_;
 wire _10746_;
 wire _10747_;
 wire _10748_;
 wire _10749_;
 wire _10750_;
 wire _10751_;
 wire _10752_;
 wire _10753_;
 wire _10754_;
 wire _10755_;
 wire _10756_;
 wire _10757_;
 wire _10758_;
 wire _10759_;
 wire _10760_;
 wire _10761_;
 wire _10762_;
 wire _10763_;
 wire _10764_;
 wire _10765_;
 wire _10766_;
 wire _10767_;
 wire _10768_;
 wire _10769_;
 wire _10770_;
 wire _10771_;
 wire _10772_;
 wire _10773_;
 wire _10774_;
 wire _10775_;
 wire _10776_;
 wire _10777_;
 wire _10778_;
 wire _10779_;
 wire _10780_;
 wire _10781_;
 wire _10782_;
 wire _10783_;
 wire _10784_;
 wire _10785_;
 wire _10786_;
 wire _10787_;
 wire _10788_;
 wire _10789_;
 wire \add0.a_i[0] ;
 wire \add0.a_i[10] ;
 wire \add0.a_i[11] ;
 wire \add0.a_i[12] ;
 wire \add0.a_i[13] ;
 wire \add0.a_i[14] ;
 wire \add0.a_i[15] ;
 wire \add0.a_i[16] ;
 wire \add0.a_i[17] ;
 wire \add0.a_i[18] ;
 wire \add0.a_i[19] ;
 wire \add0.a_i[1] ;
 wire \add0.a_i[20] ;
 wire \add0.a_i[21] ;
 wire \add0.a_i[22] ;
 wire \add0.a_i[23] ;
 wire \add0.a_i[24] ;
 wire \add0.a_i[25] ;
 wire \add0.a_i[26] ;
 wire \add0.a_i[27] ;
 wire \add0.a_i[28] ;
 wire \add0.a_i[29] ;
 wire \add0.a_i[2] ;
 wire \add0.a_i[30] ;
 wire \add0.a_i[31] ;
 wire \add0.a_i[3] ;
 wire \add0.a_i[4] ;
 wire \add0.a_i[5] ;
 wire \add0.a_i[6] ;
 wire \add0.a_i[7] ;
 wire \add0.a_i[8] ;
 wire \add0.a_i[9] ;
 wire \add0.b_i[0] ;
 wire \add0.b_i[10] ;
 wire \add0.b_i[11] ;
 wire \add0.b_i[12] ;
 wire \add0.b_i[13] ;
 wire \add0.b_i[14] ;
 wire \add0.b_i[15] ;
 wire \add0.b_i[16] ;
 wire \add0.b_i[17] ;
 wire \add0.b_i[18] ;
 wire \add0.b_i[19] ;
 wire \add0.b_i[1] ;
 wire \add0.b_i[20] ;
 wire \add0.b_i[21] ;
 wire \add0.b_i[22] ;
 wire \add0.b_i[23] ;
 wire \add0.b_i[24] ;
 wire \add0.b_i[25] ;
 wire \add0.b_i[26] ;
 wire \add0.b_i[27] ;
 wire \add0.b_i[28] ;
 wire \add0.b_i[29] ;
 wire \add0.b_i[2] ;
 wire \add0.b_i[30] ;
 wire \add0.b_i[31] ;
 wire \add0.b_i[3] ;
 wire \add0.b_i[4] ;
 wire \add0.b_i[5] ;
 wire \add0.b_i[6] ;
 wire \add0.b_i[7] ;
 wire \add0.b_i[8] ;
 wire \add0.b_i[9] ;
 wire clknet_0_clk_i;
 wire clknet_2_0__leaf_clk_i;
 wire clknet_2_1__leaf_clk_i;
 wire clknet_2_2__leaf_clk_i;
 wire clknet_2_3__leaf_clk_i;
 wire clknet_leaf_0_clk_i;
 wire clknet_leaf_10_clk_i;
 wire clknet_leaf_11_clk_i;
 wire clknet_leaf_12_clk_i;
 wire clknet_leaf_13_clk_i;
 wire clknet_leaf_14_clk_i;
 wire clknet_leaf_15_clk_i;
 wire clknet_leaf_16_clk_i;
 wire clknet_leaf_17_clk_i;
 wire clknet_leaf_18_clk_i;
 wire clknet_leaf_19_clk_i;
 wire clknet_leaf_1_clk_i;
 wire clknet_leaf_20_clk_i;
 wire clknet_leaf_21_clk_i;
 wire clknet_leaf_22_clk_i;
 wire clknet_leaf_23_clk_i;
 wire clknet_leaf_24_clk_i;
 wire clknet_leaf_25_clk_i;
 wire clknet_leaf_26_clk_i;
 wire clknet_leaf_27_clk_i;
 wire clknet_leaf_28_clk_i;
 wire clknet_leaf_29_clk_i;
 wire clknet_leaf_2_clk_i;
 wire clknet_leaf_30_clk_i;
 wire clknet_leaf_31_clk_i;
 wire clknet_leaf_32_clk_i;
 wire clknet_leaf_33_clk_i;
 wire clknet_leaf_34_clk_i;
 wire clknet_leaf_35_clk_i;
 wire clknet_leaf_36_clk_i;
 wire clknet_leaf_37_clk_i;
 wire clknet_leaf_38_clk_i;
 wire clknet_leaf_3_clk_i;
 wire clknet_leaf_40_clk_i;
 wire clknet_leaf_41_clk_i;
 wire clknet_leaf_43_clk_i;
 wire clknet_leaf_44_clk_i;
 wire clknet_leaf_4_clk_i;
 wire clknet_leaf_5_clk_i;
 wire clknet_leaf_6_clk_i;
 wire clknet_leaf_7_clk_i;
 wire clknet_leaf_9_clk_i;
 wire \depth[0] ;
 wire \depth[10] ;
 wire \depth[11] ;
 wire \depth[12] ;
 wire \depth[13] ;
 wire \depth[14] ;
 wire \depth[15] ;
 wire \depth[16] ;
 wire \depth[17] ;
 wire \depth[18] ;
 wire \depth[19] ;
 wire \depth[1] ;
 wire \depth[20] ;
 wire \depth[21] ;
 wire \depth[22] ;
 wire \depth[23] ;
 wire \depth[24] ;
 wire \depth[25] ;
 wire \depth[26] ;
 wire \depth[27] ;
 wire \depth[28] ;
 wire \depth[29] ;
 wire \depth[2] ;
 wire \depth[30] ;
 wire \depth[31] ;
 wire \depth[3] ;
 wire \depth[4] ;
 wire \depth[5] ;
 wire \depth[6] ;
 wire \depth[7] ;
 wire \depth[8] ;
 wire \depth[9] ;
 wire \in_data[0] ;
 wire \in_data[100] ;
 wire \in_data[101] ;
 wire \in_data[102] ;
 wire \in_data[103] ;
 wire \in_data[104] ;
 wire \in_data[105] ;
 wire \in_data[106] ;
 wire \in_data[107] ;
 wire \in_data[108] ;
 wire \in_data[109] ;
 wire \in_data[10] ;
 wire \in_data[110] ;
 wire \in_data[111] ;
 wire \in_data[112] ;
 wire \in_data[113] ;
 wire \in_data[11] ;
 wire \in_data[12] ;
 wire \in_data[13] ;
 wire \in_data[14] ;
 wire \in_data[15] ;
 wire \in_data[16] ;
 wire \in_data[17] ;
 wire \in_data[18] ;
 wire \in_data[19] ;
 wire \in_data[1] ;
 wire \in_data[20] ;
 wire \in_data[21] ;
 wire \in_data[22] ;
 wire \in_data[23] ;
 wire \in_data[24] ;
 wire \in_data[25] ;
 wire \in_data[26] ;
 wire \in_data[27] ;
 wire \in_data[28] ;
 wire \in_data[29] ;
 wire \in_data[2] ;
 wire \in_data[30] ;
 wire \in_data[31] ;
 wire \in_data[32] ;
 wire \in_data[33] ;
 wire \in_data[34] ;
 wire \in_data[35] ;
 wire \in_data[36] ;
 wire \in_data[37] ;
 wire \in_data[38] ;
 wire \in_data[39] ;
 wire \in_data[3] ;
 wire \in_data[40] ;
 wire \in_data[41] ;
 wire \in_data[42] ;
 wire \in_data[43] ;
 wire \in_data[44] ;
 wire \in_data[45] ;
 wire \in_data[46] ;
 wire \in_data[47] ;
 wire \in_data[48] ;
 wire \in_data[49] ;
 wire \in_data[4] ;
 wire \in_data[50] ;
 wire \in_data[51] ;
 wire \in_data[52] ;
 wire \in_data[53] ;
 wire \in_data[54] ;
 wire \in_data[55] ;
 wire \in_data[56] ;
 wire \in_data[57] ;
 wire \in_data[58] ;
 wire \in_data[59] ;
 wire \in_data[5] ;
 wire \in_data[60] ;
 wire \in_data[61] ;
 wire \in_data[62] ;
 wire \in_data[63] ;
 wire \in_data[64] ;
 wire \in_data[65] ;
 wire \in_data[66] ;
 wire \in_data[67] ;
 wire \in_data[68] ;
 wire \in_data[69] ;
 wire \in_data[6] ;
 wire \in_data[70] ;
 wire \in_data[71] ;
 wire \in_data[72] ;
 wire \in_data[73] ;
 wire \in_data[74] ;
 wire \in_data[75] ;
 wire \in_data[76] ;
 wire \in_data[77] ;
 wire \in_data[78] ;
 wire \in_data[79] ;
 wire \in_data[7] ;
 wire \in_data[80] ;
 wire \in_data[81] ;
 wire \in_data[82] ;
 wire \in_data[83] ;
 wire \in_data[84] ;
 wire \in_data[85] ;
 wire \in_data[86] ;
 wire \in_data[87] ;
 wire \in_data[88] ;
 wire \in_data[89] ;
 wire \in_data[8] ;
 wire \in_data[90] ;
 wire \in_data[91] ;
 wire \in_data[92] ;
 wire \in_data[93] ;
 wire \in_data[94] ;
 wire \in_data[95] ;
 wire \in_data[96] ;
 wire \in_data[97] ;
 wire \in_data[98] ;
 wire \in_data[99] ;
 wire \in_data[9] ;
 wire \mul0.a[0] ;
 wire \mul0.a[10] ;
 wire \mul0.a[11] ;
 wire \mul0.a[12] ;
 wire \mul0.a[13] ;
 wire \mul0.a[14] ;
 wire \mul0.a[15] ;
 wire \mul0.a[16] ;
 wire \mul0.a[17] ;
 wire \mul0.a[18] ;
 wire \mul0.a[19] ;
 wire \mul0.a[1] ;
 wire \mul0.a[20] ;
 wire \mul0.a[21] ;
 wire \mul0.a[22] ;
 wire \mul0.a[23] ;
 wire \mul0.a[24] ;
 wire \mul0.a[25] ;
 wire \mul0.a[26] ;
 wire \mul0.a[27] ;
 wire \mul0.a[28] ;
 wire \mul0.a[29] ;
 wire \mul0.a[2] ;
 wire \mul0.a[30] ;
 wire \mul0.a[31] ;
 wire \mul0.a[3] ;
 wire \mul0.a[4] ;
 wire \mul0.a[5] ;
 wire \mul0.a[6] ;
 wire \mul0.a[7] ;
 wire \mul0.a[8] ;
 wire \mul0.a[9] ;
 wire \mul0.b[0] ;
 wire \mul0.b[10] ;
 wire \mul0.b[11] ;
 wire \mul0.b[12] ;
 wire \mul0.b[13] ;
 wire \mul0.b[14] ;
 wire \mul0.b[15] ;
 wire \mul0.b[16] ;
 wire \mul0.b[17] ;
 wire \mul0.b[18] ;
 wire \mul0.b[19] ;
 wire \mul0.b[1] ;
 wire \mul0.b[20] ;
 wire \mul0.b[21] ;
 wire \mul0.b[22] ;
 wire \mul0.b[23] ;
 wire \mul0.b[24] ;
 wire \mul0.b[25] ;
 wire \mul0.b[26] ;
 wire \mul0.b[27] ;
 wire \mul0.b[28] ;
 wire \mul0.b[29] ;
 wire \mul0.b[2] ;
 wire \mul0.b[30] ;
 wire \mul0.b[31] ;
 wire \mul0.b[3] ;
 wire \mul0.b[4] ;
 wire \mul0.b[5] ;
 wire \mul0.b[6] ;
 wire \mul0.b[7] ;
 wire \mul0.b[8] ;
 wire \mul0.b[9] ;
 wire \mul1.a[0] ;
 wire \mul1.a[10] ;
 wire \mul1.a[11] ;
 wire \mul1.a[12] ;
 wire \mul1.a[13] ;
 wire \mul1.a[14] ;
 wire \mul1.a[15] ;
 wire \mul1.a[16] ;
 wire \mul1.a[17] ;
 wire \mul1.a[18] ;
 wire \mul1.a[19] ;
 wire \mul1.a[1] ;
 wire \mul1.a[20] ;
 wire \mul1.a[21] ;
 wire \mul1.a[22] ;
 wire \mul1.a[23] ;
 wire \mul1.a[24] ;
 wire \mul1.a[25] ;
 wire \mul1.a[26] ;
 wire \mul1.a[27] ;
 wire \mul1.a[28] ;
 wire \mul1.a[29] ;
 wire \mul1.a[2] ;
 wire \mul1.a[30] ;
 wire \mul1.a[31] ;
 wire \mul1.a[3] ;
 wire \mul1.a[4] ;
 wire \mul1.a[5] ;
 wire \mul1.a[6] ;
 wire \mul1.a[7] ;
 wire \mul1.a[8] ;
 wire \mul1.a[9] ;
 wire \mul1.b[0] ;
 wire \mul1.b[10] ;
 wire \mul1.b[11] ;
 wire \mul1.b[12] ;
 wire \mul1.b[13] ;
 wire \mul1.b[14] ;
 wire \mul1.b[15] ;
 wire \mul1.b[16] ;
 wire \mul1.b[17] ;
 wire \mul1.b[18] ;
 wire \mul1.b[19] ;
 wire \mul1.b[1] ;
 wire \mul1.b[20] ;
 wire \mul1.b[21] ;
 wire \mul1.b[22] ;
 wire \mul1.b[23] ;
 wire \mul1.b[24] ;
 wire \mul1.b[25] ;
 wire \mul1.b[26] ;
 wire \mul1.b[27] ;
 wire \mul1.b[28] ;
 wire \mul1.b[29] ;
 wire \mul1.b[2] ;
 wire \mul1.b[30] ;
 wire \mul1.b[31] ;
 wire \mul1.b[3] ;
 wire \mul1.b[4] ;
 wire \mul1.b[5] ;
 wire \mul1.b[6] ;
 wire \mul1.b[7] ;
 wire \mul1.b[8] ;
 wire \mul1.b[9] ;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net15;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net16;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net17;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net18;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net19;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net2;
 wire net20;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net21;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net22;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net23;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net24;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net25;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net26;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net27;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net28;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net29;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net3;
 wire net30;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net31;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net32;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net33;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net34;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net35;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net36;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net37;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net38;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net39;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net4;
 wire net40;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net41;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net42;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net43;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net44;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net45;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net46;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net47;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net48;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net49;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net5;
 wire net50;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net51;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net52;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net53;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net54;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net55;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net56;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net57;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net58;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net59;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net6;
 wire net60;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net61;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net62;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net63;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net64;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net65;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net66;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net67;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net68;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net69;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net7;
 wire net70;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net71;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net72;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net73;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net74;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net75;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net76;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net77;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net78;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net79;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net8;
 wire net80;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net81;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net82;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net83;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net84;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net85;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net86;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net87;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net88;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net89;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net9;
 wire net90;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net91;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net92;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net93;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net94;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net95;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net96;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net97;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net98;
 wire net99;
 wire \state[1] ;
 wire \state[2] ;
 wire \state[3] ;
 wire \state[4] ;
 wire \state[5] ;
 wire \state[7] ;
 wire \state[8] ;
 wire \state[9] ;
 wire \temp[0] ;
 wire \temp[10] ;
 wire \temp[11] ;
 wire \temp[12] ;
 wire \temp[13] ;
 wire \temp[14] ;
 wire \temp[15] ;
 wire \temp[16] ;
 wire \temp[17] ;
 wire \temp[18] ;
 wire \temp[19] ;
 wire \temp[1] ;
 wire \temp[20] ;
 wire \temp[21] ;
 wire \temp[22] ;
 wire \temp[23] ;
 wire \temp[24] ;
 wire \temp[25] ;
 wire \temp[26] ;
 wire \temp[27] ;
 wire \temp[28] ;
 wire \temp[29] ;
 wire \temp[2] ;
 wire \temp[30] ;
 wire \temp[31] ;
 wire \temp[3] ;
 wire \temp[4] ;
 wire \temp[5] ;
 wire \temp[6] ;
 wire \temp[7] ;
 wire \temp[8] ;
 wire \temp[9] ;
 wire \tx[0] ;
 wire \tx[10] ;
 wire \tx[11] ;
 wire \tx[12] ;
 wire \tx[13] ;
 wire \tx[14] ;
 wire \tx[15] ;
 wire \tx[16] ;
 wire \tx[17] ;
 wire \tx[18] ;
 wire \tx[19] ;
 wire \tx[1] ;
 wire \tx[20] ;
 wire \tx[21] ;
 wire \tx[22] ;
 wire \tx[23] ;
 wire \tx[24] ;
 wire \tx[25] ;
 wire \tx[26] ;
 wire \tx[27] ;
 wire \tx[28] ;
 wire \tx[29] ;
 wire \tx[2] ;
 wire \tx[30] ;
 wire \tx[31] ;
 wire \tx[3] ;
 wire \tx[4] ;
 wire \tx[5] ;
 wire \tx[6] ;
 wire \tx[7] ;
 wire \tx[8] ;
 wire \tx[9] ;

 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(_00000_));
 sky130_fd_sc_hd__diode_2 ANTENNA_10 (.DIODE(_02904_));
 sky130_fd_sc_hd__diode_2 ANTENNA_100 (.DIODE(mstream_o[115]));
 sky130_fd_sc_hd__diode_2 ANTENNA_101 (.DIODE(mstream_o[115]));
 sky130_fd_sc_hd__diode_2 ANTENNA_102 (.DIODE(mstream_o[115]));
 sky130_fd_sc_hd__diode_2 ANTENNA_103 (.DIODE(mstream_o[115]));
 sky130_fd_sc_hd__diode_2 ANTENNA_104 (.DIODE(mstream_o[115]));
 sky130_fd_sc_hd__diode_2 ANTENNA_105 (.DIODE(\mul1.a[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_106 (.DIODE(sstream_i[26]));
 sky130_fd_sc_hd__diode_2 ANTENNA_107 (.DIODE(sstream_i[28]));
 sky130_fd_sc_hd__diode_2 ANTENNA_108 (.DIODE(sstream_i[29]));
 sky130_fd_sc_hd__diode_2 ANTENNA_109 (.DIODE(sstream_i[30]));
 sky130_fd_sc_hd__diode_2 ANTENNA_11 (.DIODE(_02904_));
 sky130_fd_sc_hd__diode_2 ANTENNA_110 (.DIODE(sstream_i[31]));
 sky130_fd_sc_hd__diode_2 ANTENNA_111 (.DIODE(sstream_i[64]));
 sky130_fd_sc_hd__diode_2 ANTENNA_112 (.DIODE(sstream_i[65]));
 sky130_fd_sc_hd__diode_2 ANTENNA_113 (.DIODE(sstream_i[66]));
 sky130_fd_sc_hd__diode_2 ANTENNA_114 (.DIODE(sstream_i[67]));
 sky130_fd_sc_hd__diode_2 ANTENNA_115 (.DIODE(sstream_i[68]));
 sky130_fd_sc_hd__diode_2 ANTENNA_116 (.DIODE(sstream_i[69]));
 sky130_fd_sc_hd__diode_2 ANTENNA_117 (.DIODE(sstream_i[70]));
 sky130_fd_sc_hd__diode_2 ANTENNA_118 (.DIODE(sstream_i[71]));
 sky130_fd_sc_hd__diode_2 ANTENNA_119 (.DIODE(v0z[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_12 (.DIODE(_02904_));
 sky130_fd_sc_hd__diode_2 ANTENNA_120 (.DIODE(v0z[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA_121 (.DIODE(v0z[14]));
 sky130_fd_sc_hd__diode_2 ANTENNA_122 (.DIODE(v0z[15]));
 sky130_fd_sc_hd__diode_2 ANTENNA_123 (.DIODE(v0z[18]));
 sky130_fd_sc_hd__diode_2 ANTENNA_124 (.DIODE(v0z[23]));
 sky130_fd_sc_hd__diode_2 ANTENNA_125 (.DIODE(v0z[27]));
 sky130_fd_sc_hd__diode_2 ANTENNA_126 (.DIODE(v0z[28]));
 sky130_fd_sc_hd__diode_2 ANTENNA_127 (.DIODE(v0z[30]));
 sky130_fd_sc_hd__diode_2 ANTENNA_128 (.DIODE(v1z[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_129 (.DIODE(v1z[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA_13 (.DIODE(_02904_));
 sky130_fd_sc_hd__diode_2 ANTENNA_130 (.DIODE(v1z[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA_131 (.DIODE(v1z[14]));
 sky130_fd_sc_hd__diode_2 ANTENNA_132 (.DIODE(v1z[15]));
 sky130_fd_sc_hd__diode_2 ANTENNA_133 (.DIODE(v1z[17]));
 sky130_fd_sc_hd__diode_2 ANTENNA_134 (.DIODE(v1z[17]));
 sky130_fd_sc_hd__diode_2 ANTENNA_135 (.DIODE(v1z[18]));
 sky130_fd_sc_hd__diode_2 ANTENNA_136 (.DIODE(v1z[19]));
 sky130_fd_sc_hd__diode_2 ANTENNA_137 (.DIODE(v1z[20]));
 sky130_fd_sc_hd__diode_2 ANTENNA_138 (.DIODE(v1z[21]));
 sky130_fd_sc_hd__diode_2 ANTENNA_139 (.DIODE(v1z[22]));
 sky130_fd_sc_hd__diode_2 ANTENNA_14 (.DIODE(_02907_));
 sky130_fd_sc_hd__diode_2 ANTENNA_140 (.DIODE(v1z[23]));
 sky130_fd_sc_hd__diode_2 ANTENNA_141 (.DIODE(v1z[24]));
 sky130_fd_sc_hd__diode_2 ANTENNA_142 (.DIODE(v1z[25]));
 sky130_fd_sc_hd__diode_2 ANTENNA_143 (.DIODE(v1z[26]));
 sky130_fd_sc_hd__diode_2 ANTENNA_144 (.DIODE(v1z[27]));
 sky130_fd_sc_hd__diode_2 ANTENNA_145 (.DIODE(v1z[28]));
 sky130_fd_sc_hd__diode_2 ANTENNA_146 (.DIODE(v1z[29]));
 sky130_fd_sc_hd__diode_2 ANTENNA_147 (.DIODE(v1z[30]));
 sky130_fd_sc_hd__diode_2 ANTENNA_148 (.DIODE(v1z[31]));
 sky130_fd_sc_hd__diode_2 ANTENNA_149 (.DIODE(v1z[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_15 (.DIODE(_02907_));
 sky130_fd_sc_hd__diode_2 ANTENNA_150 (.DIODE(v1z[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_151 (.DIODE(v1z[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_152 (.DIODE(v1z[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_153 (.DIODE(v1z[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_154 (.DIODE(v2z[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_155 (.DIODE(v2z[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA_156 (.DIODE(v2z[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA_157 (.DIODE(v2z[14]));
 sky130_fd_sc_hd__diode_2 ANTENNA_158 (.DIODE(v2z[14]));
 sky130_fd_sc_hd__diode_2 ANTENNA_159 (.DIODE(v2z[15]));
 sky130_fd_sc_hd__diode_2 ANTENNA_16 (.DIODE(_02907_));
 sky130_fd_sc_hd__diode_2 ANTENNA_160 (.DIODE(v2z[16]));
 sky130_fd_sc_hd__diode_2 ANTENNA_161 (.DIODE(v2z[17]));
 sky130_fd_sc_hd__diode_2 ANTENNA_162 (.DIODE(v2z[18]));
 sky130_fd_sc_hd__diode_2 ANTENNA_163 (.DIODE(v2z[18]));
 sky130_fd_sc_hd__diode_2 ANTENNA_164 (.DIODE(v2z[19]));
 sky130_fd_sc_hd__diode_2 ANTENNA_165 (.DIODE(v2z[20]));
 sky130_fd_sc_hd__diode_2 ANTENNA_166 (.DIODE(v2z[21]));
 sky130_fd_sc_hd__diode_2 ANTENNA_167 (.DIODE(v2z[21]));
 sky130_fd_sc_hd__diode_2 ANTENNA_168 (.DIODE(v2z[22]));
 sky130_fd_sc_hd__diode_2 ANTENNA_169 (.DIODE(v2z[23]));
 sky130_fd_sc_hd__diode_2 ANTENNA_17 (.DIODE(_02907_));
 sky130_fd_sc_hd__diode_2 ANTENNA_170 (.DIODE(v2z[24]));
 sky130_fd_sc_hd__diode_2 ANTENNA_171 (.DIODE(v2z[25]));
 sky130_fd_sc_hd__diode_2 ANTENNA_172 (.DIODE(v2z[26]));
 sky130_fd_sc_hd__diode_2 ANTENNA_173 (.DIODE(v2z[27]));
 sky130_fd_sc_hd__diode_2 ANTENNA_174 (.DIODE(v2z[28]));
 sky130_fd_sc_hd__diode_2 ANTENNA_175 (.DIODE(v2z[28]));
 sky130_fd_sc_hd__diode_2 ANTENNA_176 (.DIODE(v2z[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_177 (.DIODE(v2z[30]));
 sky130_fd_sc_hd__diode_2 ANTENNA_178 (.DIODE(v2z[31]));
 sky130_fd_sc_hd__diode_2 ANTENNA_179 (.DIODE(v2z[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_18 (.DIODE(_02907_));
 sky130_fd_sc_hd__diode_2 ANTENNA_180 (.DIODE(v2z[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_181 (.DIODE(v2z[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_182 (.DIODE(v2z[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_183 (.DIODE(net547));
 sky130_fd_sc_hd__diode_2 ANTENNA_184 (.DIODE(net885));
 sky130_fd_sc_hd__diode_2 ANTENNA_185 (.DIODE(net885));
 sky130_fd_sc_hd__diode_2 ANTENNA_186 (.DIODE(net885));
 sky130_fd_sc_hd__diode_2 ANTENNA_187 (.DIODE(net885));
 sky130_fd_sc_hd__diode_2 ANTENNA_188 (.DIODE(net885));
 sky130_fd_sc_hd__diode_2 ANTENNA_189 (.DIODE(net893));
 sky130_fd_sc_hd__diode_2 ANTENNA_19 (.DIODE(_02907_));
 sky130_fd_sc_hd__diode_2 ANTENNA_190 (.DIODE(net893));
 sky130_fd_sc_hd__diode_2 ANTENNA_191 (.DIODE(net893));
 sky130_fd_sc_hd__diode_2 ANTENNA_192 (.DIODE(net893));
 sky130_fd_sc_hd__diode_2 ANTENNA_193 (.DIODE(net893));
 sky130_fd_sc_hd__diode_2 ANTENNA_194 (.DIODE(net902));
 sky130_fd_sc_hd__diode_2 ANTENNA_195 (.DIODE(net902));
 sky130_fd_sc_hd__diode_2 ANTENNA_196 (.DIODE(net902));
 sky130_fd_sc_hd__diode_2 ANTENNA_197 (.DIODE(net902));
 sky130_fd_sc_hd__diode_2 ANTENNA_198 (.DIODE(net902));
 sky130_fd_sc_hd__diode_2 ANTENNA_199 (.DIODE(net914));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(_02562_));
 sky130_fd_sc_hd__diode_2 ANTENNA_20 (.DIODE(_02910_));
 sky130_fd_sc_hd__diode_2 ANTENNA_200 (.DIODE(net914));
 sky130_fd_sc_hd__diode_2 ANTENNA_201 (.DIODE(net914));
 sky130_fd_sc_hd__diode_2 ANTENNA_202 (.DIODE(net914));
 sky130_fd_sc_hd__diode_2 ANTENNA_203 (.DIODE(net914));
 sky130_fd_sc_hd__diode_2 ANTENNA_204 (.DIODE(net916));
 sky130_fd_sc_hd__diode_2 ANTENNA_205 (.DIODE(net916));
 sky130_fd_sc_hd__diode_2 ANTENNA_206 (.DIODE(net916));
 sky130_fd_sc_hd__diode_2 ANTENNA_207 (.DIODE(net916));
 sky130_fd_sc_hd__diode_2 ANTENNA_208 (.DIODE(net916));
 sky130_fd_sc_hd__diode_2 ANTENNA_209 (.DIODE(net921));
 sky130_fd_sc_hd__diode_2 ANTENNA_21 (.DIODE(_02910_));
 sky130_fd_sc_hd__diode_2 ANTENNA_210 (.DIODE(net921));
 sky130_fd_sc_hd__diode_2 ANTENNA_211 (.DIODE(net921));
 sky130_fd_sc_hd__diode_2 ANTENNA_212 (.DIODE(net921));
 sky130_fd_sc_hd__diode_2 ANTENNA_213 (.DIODE(net921));
 sky130_fd_sc_hd__diode_2 ANTENNA_214 (.DIODE(net921));
 sky130_fd_sc_hd__diode_2 ANTENNA_215 (.DIODE(net921));
 sky130_fd_sc_hd__diode_2 ANTENNA_216 (.DIODE(net921));
 sky130_fd_sc_hd__diode_2 ANTENNA_217 (.DIODE(net923));
 sky130_fd_sc_hd__diode_2 ANTENNA_218 (.DIODE(net923));
 sky130_fd_sc_hd__diode_2 ANTENNA_219 (.DIODE(net923));
 sky130_fd_sc_hd__diode_2 ANTENNA_22 (.DIODE(_02910_));
 sky130_fd_sc_hd__diode_2 ANTENNA_220 (.DIODE(net923));
 sky130_fd_sc_hd__diode_2 ANTENNA_221 (.DIODE(net923));
 sky130_fd_sc_hd__diode_2 ANTENNA_222 (.DIODE(net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_223 (.DIODE(net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_224 (.DIODE(net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_225 (.DIODE(net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_226 (.DIODE(net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_227 (.DIODE(net936));
 sky130_fd_sc_hd__diode_2 ANTENNA_228 (.DIODE(net936));
 sky130_fd_sc_hd__diode_2 ANTENNA_229 (.DIODE(net936));
 sky130_fd_sc_hd__diode_2 ANTENNA_23 (.DIODE(_02910_));
 sky130_fd_sc_hd__diode_2 ANTENNA_230 (.DIODE(net936));
 sky130_fd_sc_hd__diode_2 ANTENNA_231 (.DIODE(net936));
 sky130_fd_sc_hd__diode_2 ANTENNA_232 (.DIODE(net945));
 sky130_fd_sc_hd__diode_2 ANTENNA_233 (.DIODE(net945));
 sky130_fd_sc_hd__diode_2 ANTENNA_234 (.DIODE(net945));
 sky130_fd_sc_hd__diode_2 ANTENNA_235 (.DIODE(net945));
 sky130_fd_sc_hd__diode_2 ANTENNA_236 (.DIODE(net945));
 sky130_fd_sc_hd__diode_2 ANTENNA_237 (.DIODE(net955));
 sky130_fd_sc_hd__diode_2 ANTENNA_238 (.DIODE(net955));
 sky130_fd_sc_hd__diode_2 ANTENNA_239 (.DIODE(net955));
 sky130_fd_sc_hd__diode_2 ANTENNA_24 (.DIODE(_02910_));
 sky130_fd_sc_hd__diode_2 ANTENNA_240 (.DIODE(net955));
 sky130_fd_sc_hd__diode_2 ANTENNA_241 (.DIODE(net955));
 sky130_fd_sc_hd__diode_2 ANTENNA_242 (.DIODE(_02916_));
 sky130_fd_sc_hd__diode_2 ANTENNA_243 (.DIODE(_02916_));
 sky130_fd_sc_hd__diode_2 ANTENNA_244 (.DIODE(_02916_));
 sky130_fd_sc_hd__diode_2 ANTENNA_245 (.DIODE(_02916_));
 sky130_fd_sc_hd__diode_2 ANTENNA_246 (.DIODE(_02916_));
 sky130_fd_sc_hd__diode_2 ANTENNA_247 (.DIODE(_02916_));
 sky130_fd_sc_hd__diode_2 ANTENNA_248 (.DIODE(\in_data[109] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_249 (.DIODE(\in_data[109] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_25 (.DIODE(_02910_));
 sky130_fd_sc_hd__diode_2 ANTENNA_250 (.DIODE(\in_data[109] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_251 (.DIODE(\mul1.b[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_252 (.DIODE(v0z[20]));
 sky130_fd_sc_hd__diode_2 ANTENNA_253 (.DIODE(v0z[22]));
 sky130_fd_sc_hd__diode_2 ANTENNA_254 (.DIODE(v2z[29]));
 sky130_fd_sc_hd__diode_2 ANTENNA_255 (.DIODE(v2z[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_256 (.DIODE(v2z[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_257 (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_258 (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_259 (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_26 (.DIODE(_02913_));
 sky130_fd_sc_hd__diode_2 ANTENNA_260 (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_261 (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_262 (.DIODE(net932));
 sky130_fd_sc_hd__diode_2 ANTENNA_263 (.DIODE(net932));
 sky130_fd_sc_hd__diode_2 ANTENNA_264 (.DIODE(net932));
 sky130_fd_sc_hd__diode_2 ANTENNA_265 (.DIODE(net932));
 sky130_fd_sc_hd__diode_2 ANTENNA_266 (.DIODE(net932));
 sky130_fd_sc_hd__diode_2 ANTENNA_267 (.DIODE(net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_268 (.DIODE(net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_269 (.DIODE(net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_27 (.DIODE(_02913_));
 sky130_fd_sc_hd__diode_2 ANTENNA_270 (.DIODE(net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_271 (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_272 (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_273 (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_274 (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_275 (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_276 (.DIODE(v0z[19]));
 sky130_fd_sc_hd__diode_2 ANTENNA_277 (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA_278 (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA_279 (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA_28 (.DIODE(_02913_));
 sky130_fd_sc_hd__diode_2 ANTENNA_280 (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA_281 (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA_282 (.DIODE(net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_283 (.DIODE(net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_284 (.DIODE(net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_285 (.DIODE(net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_286 (.DIODE(net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_287 (.DIODE(net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_288 (.DIODE(net920));
 sky130_fd_sc_hd__diode_2 ANTENNA_289 (.DIODE(net920));
 sky130_fd_sc_hd__diode_2 ANTENNA_29 (.DIODE(_02913_));
 sky130_fd_sc_hd__diode_2 ANTENNA_290 (.DIODE(net920));
 sky130_fd_sc_hd__diode_2 ANTENNA_291 (.DIODE(net920));
 sky130_fd_sc_hd__diode_2 ANTENNA_292 (.DIODE(net920));
 sky130_fd_sc_hd__diode_2 ANTENNA_293 (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_294 (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_295 (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_296 (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_297 (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_298 (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_299 (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(_02562_));
 sky130_fd_sc_hd__diode_2 ANTENNA_30 (.DIODE(_02913_));
 sky130_fd_sc_hd__diode_2 ANTENNA_300 (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_301 (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_302 (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_303 (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_304 (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_305 (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_306 (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_307 (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_308 (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_309 (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_31 (.DIODE(_02913_));
 sky130_fd_sc_hd__diode_2 ANTENNA_310 (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_311 (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_312 (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_313 (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_314 (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_315 (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_316 (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_317 (.DIODE(net920));
 sky130_fd_sc_hd__diode_2 ANTENNA_318 (.DIODE(net920));
 sky130_fd_sc_hd__diode_2 ANTENNA_319 (.DIODE(net920));
 sky130_fd_sc_hd__diode_2 ANTENNA_32 (.DIODE(_02960_));
 sky130_fd_sc_hd__diode_2 ANTENNA_320 (.DIODE(net920));
 sky130_fd_sc_hd__diode_2 ANTENNA_321 (.DIODE(net920));
 sky130_fd_sc_hd__diode_2 ANTENNA_322 (.DIODE(net920));
 sky130_fd_sc_hd__diode_2 ANTENNA_323 (.DIODE(net920));
 sky130_fd_sc_hd__diode_2 ANTENNA_324 (.DIODE(net920));
 sky130_fd_sc_hd__diode_2 ANTENNA_325 (.DIODE(net920));
 sky130_fd_sc_hd__diode_2 ANTENNA_326 (.DIODE(net920));
 sky130_fd_sc_hd__diode_2 ANTENNA_327 (.DIODE(net920));
 sky130_fd_sc_hd__diode_2 ANTENNA_328 (.DIODE(net920));
 sky130_fd_sc_hd__diode_2 ANTENNA_329 (.DIODE(net920));
 sky130_fd_sc_hd__diode_2 ANTENNA_33 (.DIODE(_02960_));
 sky130_fd_sc_hd__diode_2 ANTENNA_330 (.DIODE(net920));
 sky130_fd_sc_hd__diode_2 ANTENNA_331 (.DIODE(net920));
 sky130_fd_sc_hd__diode_2 ANTENNA_332 (.DIODE(net920));
 sky130_fd_sc_hd__diode_2 ANTENNA_333 (.DIODE(net920));
 sky130_fd_sc_hd__diode_2 ANTENNA_334 (.DIODE(net920));
 sky130_fd_sc_hd__diode_2 ANTENNA_335 (.DIODE(net920));
 sky130_fd_sc_hd__diode_2 ANTENNA_336 (.DIODE(net920));
 sky130_fd_sc_hd__diode_2 ANTENNA_337 (.DIODE(net920));
 sky130_fd_sc_hd__diode_2 ANTENNA_338 (.DIODE(net920));
 sky130_fd_sc_hd__diode_2 ANTENNA_339 (.DIODE(net920));
 sky130_fd_sc_hd__diode_2 ANTENNA_34 (.DIODE(_02960_));
 sky130_fd_sc_hd__diode_2 ANTENNA_340 (.DIODE(net920));
 sky130_fd_sc_hd__diode_2 ANTENNA_35 (.DIODE(_02972_));
 sky130_fd_sc_hd__diode_2 ANTENNA_36 (.DIODE(_02972_));
 sky130_fd_sc_hd__diode_2 ANTENNA_37 (.DIODE(_02972_));
 sky130_fd_sc_hd__diode_2 ANTENNA_38 (.DIODE(_02976_));
 sky130_fd_sc_hd__diode_2 ANTENNA_39 (.DIODE(_02976_));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(_02562_));
 sky130_fd_sc_hd__diode_2 ANTENNA_40 (.DIODE(_02976_));
 sky130_fd_sc_hd__diode_2 ANTENNA_41 (.DIODE(_02982_));
 sky130_fd_sc_hd__diode_2 ANTENNA_42 (.DIODE(_02982_));
 sky130_fd_sc_hd__diode_2 ANTENNA_43 (.DIODE(_02982_));
 sky130_fd_sc_hd__diode_2 ANTENNA_44 (.DIODE(\in_data[101] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_45 (.DIODE(\in_data[101] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_46 (.DIODE(\in_data[101] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_47 (.DIODE(\in_data[101] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_48 (.DIODE(\in_data[101] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_49 (.DIODE(\in_data[101] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_5 (.DIODE(_02895_));
 sky130_fd_sc_hd__diode_2 ANTENNA_50 (.DIODE(\in_data[102] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_51 (.DIODE(\in_data[102] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_52 (.DIODE(\in_data[102] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_53 (.DIODE(\in_data[102] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_54 (.DIODE(\in_data[102] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_55 (.DIODE(\in_data[102] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_56 (.DIODE(\in_data[105] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_57 (.DIODE(\in_data[105] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_58 (.DIODE(\in_data[105] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_59 (.DIODE(\in_data[105] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_6 (.DIODE(_02895_));
 sky130_fd_sc_hd__diode_2 ANTENNA_60 (.DIODE(\in_data[105] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_61 (.DIODE(\in_data[105] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_62 (.DIODE(\in_data[108] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_63 (.DIODE(\in_data[108] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_64 (.DIODE(\in_data[108] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_65 (.DIODE(\in_data[108] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_66 (.DIODE(\in_data[108] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_67 (.DIODE(\in_data[108] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_68 (.DIODE(\in_data[111] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_69 (.DIODE(\in_data[111] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_7 (.DIODE(_02895_));
 sky130_fd_sc_hd__diode_2 ANTENNA_70 (.DIODE(\in_data[111] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_71 (.DIODE(\in_data[111] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_72 (.DIODE(\in_data[111] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_73 (.DIODE(\in_data[111] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_74 (.DIODE(\in_data[112] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_75 (.DIODE(\in_data[112] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_76 (.DIODE(\in_data[112] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_77 (.DIODE(\in_data[112] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_78 (.DIODE(\in_data[112] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_79 (.DIODE(\in_data[112] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_8 (.DIODE(_02904_));
 sky130_fd_sc_hd__diode_2 ANTENNA_80 (.DIODE(\in_data[96] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_81 (.DIODE(\in_data[96] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_82 (.DIODE(\in_data[96] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_83 (.DIODE(mstream_o[115]));
 sky130_fd_sc_hd__diode_2 ANTENNA_84 (.DIODE(mstream_o[115]));
 sky130_fd_sc_hd__diode_2 ANTENNA_85 (.DIODE(mstream_o[115]));
 sky130_fd_sc_hd__diode_2 ANTENNA_86 (.DIODE(mstream_o[115]));
 sky130_fd_sc_hd__diode_2 ANTENNA_87 (.DIODE(mstream_o[115]));
 sky130_fd_sc_hd__diode_2 ANTENNA_88 (.DIODE(mstream_o[115]));
 sky130_fd_sc_hd__diode_2 ANTENNA_89 (.DIODE(mstream_o[115]));
 sky130_fd_sc_hd__diode_2 ANTENNA_9 (.DIODE(_02904_));
 sky130_fd_sc_hd__diode_2 ANTENNA_90 (.DIODE(mstream_o[115]));
 sky130_fd_sc_hd__diode_2 ANTENNA_91 (.DIODE(mstream_o[115]));
 sky130_fd_sc_hd__diode_2 ANTENNA_92 (.DIODE(mstream_o[115]));
 sky130_fd_sc_hd__diode_2 ANTENNA_93 (.DIODE(mstream_o[115]));
 sky130_fd_sc_hd__diode_2 ANTENNA_94 (.DIODE(mstream_o[115]));
 sky130_fd_sc_hd__diode_2 ANTENNA_95 (.DIODE(mstream_o[115]));
 sky130_fd_sc_hd__diode_2 ANTENNA_96 (.DIODE(mstream_o[115]));
 sky130_fd_sc_hd__diode_2 ANTENNA_97 (.DIODE(mstream_o[115]));
 sky130_fd_sc_hd__diode_2 ANTENNA_98 (.DIODE(mstream_o[115]));
 sky130_fd_sc_hd__diode_2 ANTENNA_99 (.DIODE(mstream_o[115]));
 sky130_fd_sc_hd__diode_2 ANTENNA__10791__A (.DIODE(net598));
 sky130_fd_sc_hd__diode_2 ANTENNA__10793__A (.DIODE(net510));
 sky130_fd_sc_hd__diode_2 ANTENNA__10794__A (.DIODE(net374));
 sky130_fd_sc_hd__diode_2 ANTENNA__10795__A (.DIODE(net628));
 sky130_fd_sc_hd__diode_2 ANTENNA__10796__A (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__10797__A (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA__10798__A (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__10800__B2 (.DIODE(_02562_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10853__A1 (.DIODE(_02619_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10861__A1 (.DIODE(_02626_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10868__A1 (.DIODE(_02632_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10875__A1 (.DIODE(_02638_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10882__A1 (.DIODE(_02644_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10887__A1 (.DIODE(_02648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10893__A1 (.DIODE(_02653_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10904__A1 (.DIODE(_02663_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10913__A1 (.DIODE(_02671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10920__A1 (.DIODE(_02677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10927__A1 (.DIODE(_02683_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10935__A1 (.DIODE(_02690_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10942__A1 (.DIODE(_02696_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10947__A1 (.DIODE(_02700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10951__A1 (.DIODE(_02703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10960__A1 (.DIODE(_02711_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10966__A1 (.DIODE(_02716_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10973__A1 (.DIODE(_02722_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10979__A1 (.DIODE(_02727_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10985__A1 (.DIODE(_02732_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10989__A1 (.DIODE(_02735_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11022__A1 (.DIODE(net880));
 sky130_fd_sc_hd__diode_2 ANTENNA__11023__A1 (.DIODE(net904));
 sky130_fd_sc_hd__diode_2 ANTENNA__11024__A1 (.DIODE(net885));
 sky130_fd_sc_hd__diode_2 ANTENNA__11025__A1 (.DIODE(net902));
 sky130_fd_sc_hd__diode_2 ANTENNA__11026__A1 (.DIODE(net936));
 sky130_fd_sc_hd__diode_2 ANTENNA__11027__A1 (.DIODE(net893));
 sky130_fd_sc_hd__diode_2 ANTENNA__11028__A1 (.DIODE(net921));
 sky130_fd_sc_hd__diode_2 ANTENNA__11029__A1 (.DIODE(net955));
 sky130_fd_sc_hd__diode_2 ANTENNA__11030__A1 (.DIODE(net932));
 sky130_fd_sc_hd__diode_2 ANTENNA__11031__A1 (.DIODE(net916));
 sky130_fd_sc_hd__diode_2 ANTENNA__11032__A1 (.DIODE(net945));
 sky130_fd_sc_hd__diode_2 ANTENNA__11033__A1 (.DIODE(net934));
 sky130_fd_sc_hd__diode_2 ANTENNA__11034__A1 (.DIODE(net920));
 sky130_fd_sc_hd__diode_2 ANTENNA__11035__A1 (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA__11036__A1 (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA__11037__A1 (.DIODE(net914));
 sky130_fd_sc_hd__diode_2 ANTENNA__11038__A1 (.DIODE(net923));
 sky130_fd_sc_hd__diode_2 ANTENNA__11039__A1 (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA__11040__S (.DIODE(_00000_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11041__B (.DIODE(net599));
 sky130_fd_sc_hd__diode_2 ANTENNA__11044__A0 (.DIODE(_02738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11044__S (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__11046__A0 (.DIODE(_02739_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11046__S (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__11049__A0 (.DIODE(_02741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11049__S (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__11052__A0 (.DIODE(_02743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11052__S (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__11054__A0 (.DIODE(_02744_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11054__S (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__11056__A0 (.DIODE(_02745_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11056__S (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__11058__A0 (.DIODE(_02746_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11058__S (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__11060__A0 (.DIODE(_02747_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11060__S (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__11062__A0 (.DIODE(_02748_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11062__S (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__11064__A0 (.DIODE(_02749_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11064__S (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__11067__A0 (.DIODE(_02751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11067__S (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__11068__A0 (.DIODE(_02619_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11069__A0 (.DIODE(_02626_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11070__A0 (.DIODE(_02632_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11071__A0 (.DIODE(_02638_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11072__A0 (.DIODE(_02644_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11073__A0 (.DIODE(_02648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11074__A0 (.DIODE(_02653_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11075__A0 (.DIODE(_02663_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11076__A0 (.DIODE(_02671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11077__A0 (.DIODE(_02677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11078__A0 (.DIODE(_02683_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11078__S (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__11079__A0 (.DIODE(_02690_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11080__A0 (.DIODE(_02696_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11081__A0 (.DIODE(_02700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11082__A0 (.DIODE(_02703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11083__A0 (.DIODE(_02711_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11084__A0 (.DIODE(_02716_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11085__A0 (.DIODE(_02722_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11085__S (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__11086__A0 (.DIODE(_02727_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11086__S (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__11087__A0 (.DIODE(_02732_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11087__S (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__11088__A0 (.DIODE(_02735_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11089__A (.DIODE(net638));
 sky130_fd_sc_hd__diode_2 ANTENNA__11089__B (.DIODE(net611));
 sky130_fd_sc_hd__diode_2 ANTENNA__11090__A0 (.DIODE(_02738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11091__A0 (.DIODE(_02739_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11092__A0 (.DIODE(_02741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11093__A0 (.DIODE(_02743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11094__A0 (.DIODE(_02744_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11095__A0 (.DIODE(_02745_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11096__A0 (.DIODE(_02746_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11097__A0 (.DIODE(_02747_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11098__A0 (.DIODE(_02748_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11099__A0 (.DIODE(_02749_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11100__A0 (.DIODE(_02751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11101__A0 (.DIODE(_02619_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11102__A0 (.DIODE(_02626_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11103__A0 (.DIODE(_02632_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11104__A0 (.DIODE(_02638_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11105__A0 (.DIODE(_02644_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11106__A0 (.DIODE(_02648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11107__A0 (.DIODE(_02653_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11108__A0 (.DIODE(_02663_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11109__A0 (.DIODE(_02671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11110__A0 (.DIODE(_02677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11111__A0 (.DIODE(_02683_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11112__A0 (.DIODE(_02690_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11113__A0 (.DIODE(_02696_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11114__A0 (.DIODE(_02700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11115__A0 (.DIODE(_02703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11116__A0 (.DIODE(_02711_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11117__A0 (.DIODE(_02716_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11118__A0 (.DIODE(_02722_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11119__A0 (.DIODE(_02727_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11120__A0 (.DIODE(_02732_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11121__A0 (.DIODE(_02735_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11122__A (.DIODE(net598));
 sky130_fd_sc_hd__diode_2 ANTENNA__11122__B (.DIODE(net601));
 sky130_fd_sc_hd__diode_2 ANTENNA__11123__A (.DIODE(net607));
 sky130_fd_sc_hd__diode_2 ANTENNA__11125__B1 (.DIODE(net646));
 sky130_fd_sc_hd__diode_2 ANTENNA__11128__A2 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__11129__A0 (.DIODE(net582));
 sky130_fd_sc_hd__diode_2 ANTENNA__11129__S (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA__11131__A2 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__11132__A0 (.DIODE(net576));
 sky130_fd_sc_hd__diode_2 ANTENNA__11132__S (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA__11134__A2 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__11135__A0 (.DIODE(net571));
 sky130_fd_sc_hd__diode_2 ANTENNA__11135__S (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA__11137__A2 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__11138__A0 (.DIODE(net566));
 sky130_fd_sc_hd__diode_2 ANTENNA__11138__S (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA__11140__A2 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__11141__A0 (.DIODE(net561));
 sky130_fd_sc_hd__diode_2 ANTENNA__11141__S (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA__11143__A2 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__11144__A0 (.DIODE(net557));
 sky130_fd_sc_hd__diode_2 ANTENNA__11144__S (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA__11145__A2 (.DIODE(_02753_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11146__A2 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__11147__A0 (.DIODE(net553));
 sky130_fd_sc_hd__diode_2 ANTENNA__11147__S (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA__11149__A2 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__11150__A0 (.DIODE(net549));
 sky130_fd_sc_hd__diode_2 ANTENNA__11150__S (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA__11152__A2 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__11153__A0 (.DIODE(net544));
 sky130_fd_sc_hd__diode_2 ANTENNA__11153__S (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA__11155__A2 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__11156__A0 (.DIODE(net540));
 sky130_fd_sc_hd__diode_2 ANTENNA__11156__S (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA__11158__A2 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__11159__A0 (.DIODE(net535));
 sky130_fd_sc_hd__diode_2 ANTENNA__11159__S (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA__11161__A2 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__11162__S (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA__11164__A2 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__11165__A0 (.DIODE(net525));
 sky130_fd_sc_hd__diode_2 ANTENNA__11165__S (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA__11167__A2 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__11168__A0 (.DIODE(net520));
 sky130_fd_sc_hd__diode_2 ANTENNA__11168__S (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA__11169__B1 (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__11171__A0 (.DIODE(net515));
 sky130_fd_sc_hd__diode_2 ANTENNA__11171__S (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA__11173__A2 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__11174__A0 (.DIODE(net511));
 sky130_fd_sc_hd__diode_2 ANTENNA__11174__S (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA__11177__A0 (.DIODE(net507));
 sky130_fd_sc_hd__diode_2 ANTENNA__11177__S (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA__11180__A0 (.DIODE(net503));
 sky130_fd_sc_hd__diode_2 ANTENNA__11180__S (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA__11183__A0 (.DIODE(net498));
 sky130_fd_sc_hd__diode_2 ANTENNA__11183__S (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA__11186__A0 (.DIODE(net494));
 sky130_fd_sc_hd__diode_2 ANTENNA__11186__S (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA__11189__A0 (.DIODE(net490));
 sky130_fd_sc_hd__diode_2 ANTENNA__11189__S (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA__11192__A0 (.DIODE(net486));
 sky130_fd_sc_hd__diode_2 ANTENNA__11192__S (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA__11195__A0 (.DIODE(net482));
 sky130_fd_sc_hd__diode_2 ANTENNA__11195__S (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA__11198__A0 (.DIODE(net478));
 sky130_fd_sc_hd__diode_2 ANTENNA__11198__S (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA__11201__A0 (.DIODE(net474));
 sky130_fd_sc_hd__diode_2 ANTENNA__11201__S (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA__11204__A0 (.DIODE(net470));
 sky130_fd_sc_hd__diode_2 ANTENNA__11204__S (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA__11207__A0 (.DIODE(net466));
 sky130_fd_sc_hd__diode_2 ANTENNA__11207__S (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA__11210__A0 (.DIODE(net463));
 sky130_fd_sc_hd__diode_2 ANTENNA__11210__S (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA__11211__A2 (.DIODE(_02753_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11213__A0 (.DIODE(net460));
 sky130_fd_sc_hd__diode_2 ANTENNA__11213__S (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA__11215__A2 (.DIODE(_02757_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11216__A0 (.DIODE(net459));
 sky130_fd_sc_hd__diode_2 ANTENNA__11216__A1 (.DIODE(_02817_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11216__S (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA__11219__S (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA__11222__S (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA__11223__B (.DIODE(net610));
 sky130_fd_sc_hd__diode_2 ANTENNA__11224__A (.DIODE(net591));
 sky130_fd_sc_hd__diode_2 ANTENNA__11224__B (.DIODE(_02822_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11225__A1 (.DIODE(net598));
 sky130_fd_sc_hd__diode_2 ANTENNA__11225__B2 (.DIODE(net607));
 sky130_fd_sc_hd__diode_2 ANTENNA__11226__A1 (.DIODE(net587));
 sky130_fd_sc_hd__diode_2 ANTENNA__11226__B2 (.DIODE(net601));
 sky130_fd_sc_hd__diode_2 ANTENNA__11227__A1 (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__11227__A3 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__11227__B1 (.DIODE(_02825_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11228__A1 (.DIODE(_02826_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11228__S (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA__11229__A1 (.DIODE(net598));
 sky130_fd_sc_hd__diode_2 ANTENNA__11229__B2 (.DIODE(net607));
 sky130_fd_sc_hd__diode_2 ANTENNA__11230__A1 (.DIODE(net587));
 sky130_fd_sc_hd__diode_2 ANTENNA__11230__B2 (.DIODE(net601));
 sky130_fd_sc_hd__diode_2 ANTENNA__11231__A1 (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__11231__A3 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__11231__B1 (.DIODE(_02828_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11232__A1 (.DIODE(_02829_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11232__S (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA__11233__A1 (.DIODE(net598));
 sky130_fd_sc_hd__diode_2 ANTENNA__11233__B2 (.DIODE(net607));
 sky130_fd_sc_hd__diode_2 ANTENNA__11234__A1 (.DIODE(net587));
 sky130_fd_sc_hd__diode_2 ANTENNA__11234__B2 (.DIODE(net601));
 sky130_fd_sc_hd__diode_2 ANTENNA__11235__A1 (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__11235__A3 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__11235__B1 (.DIODE(_02831_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11236__A0 (.DIODE(net440));
 sky130_fd_sc_hd__diode_2 ANTENNA__11236__S (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA__11237__A1 (.DIODE(net598));
 sky130_fd_sc_hd__diode_2 ANTENNA__11237__B2 (.DIODE(net607));
 sky130_fd_sc_hd__diode_2 ANTENNA__11238__A1 (.DIODE(net587));
 sky130_fd_sc_hd__diode_2 ANTENNA__11238__B2 (.DIODE(net606));
 sky130_fd_sc_hd__diode_2 ANTENNA__11239__A1 (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__11239__A3 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__11239__B1 (.DIODE(_02834_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11240__A0 (.DIODE(net436));
 sky130_fd_sc_hd__diode_2 ANTENNA__11240__S (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA__11241__A1 (.DIODE(net598));
 sky130_fd_sc_hd__diode_2 ANTENNA__11241__B2 (.DIODE(net607));
 sky130_fd_sc_hd__diode_2 ANTENNA__11242__A1 (.DIODE(net587));
 sky130_fd_sc_hd__diode_2 ANTENNA__11242__B2 (.DIODE(net601));
 sky130_fd_sc_hd__diode_2 ANTENNA__11243__A1 (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__11243__A3 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__11243__B1 (.DIODE(_02837_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11244__A0 (.DIODE(net431));
 sky130_fd_sc_hd__diode_2 ANTENNA__11244__S (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA__11245__A1 (.DIODE(net598));
 sky130_fd_sc_hd__diode_2 ANTENNA__11245__B2 (.DIODE(net607));
 sky130_fd_sc_hd__diode_2 ANTENNA__11246__A1 (.DIODE(net592));
 sky130_fd_sc_hd__diode_2 ANTENNA__11246__B2 (.DIODE(net601));
 sky130_fd_sc_hd__diode_2 ANTENNA__11247__A1 (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__11247__A3 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__11247__B1 (.DIODE(_02840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11248__A0 (.DIODE(net426));
 sky130_fd_sc_hd__diode_2 ANTENNA__11248__S (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA__11249__A1 (.DIODE(net598));
 sky130_fd_sc_hd__diode_2 ANTENNA__11249__B2 (.DIODE(net607));
 sky130_fd_sc_hd__diode_2 ANTENNA__11250__A1 (.DIODE(net588));
 sky130_fd_sc_hd__diode_2 ANTENNA__11250__B2 (.DIODE(net601));
 sky130_fd_sc_hd__diode_2 ANTENNA__11251__A1 (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__11251__A3 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__11251__B1 (.DIODE(_02843_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11252__A0 (.DIODE(net421));
 sky130_fd_sc_hd__diode_2 ANTENNA__11252__S (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA__11253__A1 (.DIODE(net598));
 sky130_fd_sc_hd__diode_2 ANTENNA__11253__B2 (.DIODE(net607));
 sky130_fd_sc_hd__diode_2 ANTENNA__11254__A1 (.DIODE(net588));
 sky130_fd_sc_hd__diode_2 ANTENNA__11254__B2 (.DIODE(net606));
 sky130_fd_sc_hd__diode_2 ANTENNA__11255__A1 (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__11255__A3 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__11255__B1 (.DIODE(_02846_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11256__A0 (.DIODE(net417));
 sky130_fd_sc_hd__diode_2 ANTENNA__11256__S (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA__11257__A1 (.DIODE(net593));
 sky130_fd_sc_hd__diode_2 ANTENNA__11258__A1 (.DIODE(net588));
 sky130_fd_sc_hd__diode_2 ANTENNA__11258__B2 (.DIODE(net602));
 sky130_fd_sc_hd__diode_2 ANTENNA__11259__A1 (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__11259__A3 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__11259__B1 (.DIODE(_02849_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11260__A0 (.DIODE(net413));
 sky130_fd_sc_hd__diode_2 ANTENNA__11260__S (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA__11261__A1 (.DIODE(net593));
 sky130_fd_sc_hd__diode_2 ANTENNA__11262__A1 (.DIODE(net588));
 sky130_fd_sc_hd__diode_2 ANTENNA__11262__B2 (.DIODE(net602));
 sky130_fd_sc_hd__diode_2 ANTENNA__11263__A1 (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__11263__A3 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__11263__B1 (.DIODE(_02852_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11264__A0 (.DIODE(net408));
 sky130_fd_sc_hd__diode_2 ANTENNA__11264__S (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA__11265__A1 (.DIODE(net593));
 sky130_fd_sc_hd__diode_2 ANTENNA__11266__A1 (.DIODE(net588));
 sky130_fd_sc_hd__diode_2 ANTENNA__11266__B2 (.DIODE(net602));
 sky130_fd_sc_hd__diode_2 ANTENNA__11267__B1 (.DIODE(_02855_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11268__A0 (.DIODE(net404));
 sky130_fd_sc_hd__diode_2 ANTENNA__11268__S (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA__11269__A1 (.DIODE(net593));
 sky130_fd_sc_hd__diode_2 ANTENNA__11270__A1 (.DIODE(net588));
 sky130_fd_sc_hd__diode_2 ANTENNA__11270__B2 (.DIODE(net602));
 sky130_fd_sc_hd__diode_2 ANTENNA__11271__B1 (.DIODE(_02858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11272__A0 (.DIODE(net400));
 sky130_fd_sc_hd__diode_2 ANTENNA__11272__S (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA__11273__A1 (.DIODE(net593));
 sky130_fd_sc_hd__diode_2 ANTENNA__11274__B2 (.DIODE(net602));
 sky130_fd_sc_hd__diode_2 ANTENNA__11275__B1 (.DIODE(_02861_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11276__A0 (.DIODE(net396));
 sky130_fd_sc_hd__diode_2 ANTENNA__11276__S (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA__11277__A1 (.DIODE(net593));
 sky130_fd_sc_hd__diode_2 ANTENNA__11278__B2 (.DIODE(net602));
 sky130_fd_sc_hd__diode_2 ANTENNA__11279__B1 (.DIODE(_02864_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11280__A0 (.DIODE(net390));
 sky130_fd_sc_hd__diode_2 ANTENNA__11280__S (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA__11281__A1 (.DIODE(net593));
 sky130_fd_sc_hd__diode_2 ANTENNA__11282__A1 (.DIODE(net588));
 sky130_fd_sc_hd__diode_2 ANTENNA__11282__B2 (.DIODE(net602));
 sky130_fd_sc_hd__diode_2 ANTENNA__11283__B1 (.DIODE(_02867_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11284__A0 (.DIODE(net386));
 sky130_fd_sc_hd__diode_2 ANTENNA__11284__S (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA__11285__A1 (.DIODE(net593));
 sky130_fd_sc_hd__diode_2 ANTENNA__11287__B1 (.DIODE(_02870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11288__A0 (.DIODE(net381));
 sky130_fd_sc_hd__diode_2 ANTENNA__11288__S (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA__11289__A1 (.DIODE(net593));
 sky130_fd_sc_hd__diode_2 ANTENNA__11291__B1 (.DIODE(_02873_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11292__A0 (.DIODE(net375));
 sky130_fd_sc_hd__diode_2 ANTENNA__11292__S (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA__11293__A1 (.DIODE(net593));
 sky130_fd_sc_hd__diode_2 ANTENNA__11295__B1 (.DIODE(_02876_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11296__A0 (.DIODE(net371));
 sky130_fd_sc_hd__diode_2 ANTENNA__11296__A1 (.DIODE(_02877_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11296__S (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA__11297__A1 (.DIODE(net593));
 sky130_fd_sc_hd__diode_2 ANTENNA__11298__A1 (.DIODE(net591));
 sky130_fd_sc_hd__diode_2 ANTENNA__11299__B1 (.DIODE(_02879_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11300__A0 (.DIODE(net631));
 sky130_fd_sc_hd__diode_2 ANTENNA__11300__A1 (.DIODE(_02880_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11300__S (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA__11301__A1 (.DIODE(net593));
 sky130_fd_sc_hd__diode_2 ANTENNA__11302__A1 (.DIODE(net591));
 sky130_fd_sc_hd__diode_2 ANTENNA__11303__B1 (.DIODE(_02882_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11304__A0 (.DIODE(net365));
 sky130_fd_sc_hd__diode_2 ANTENNA__11304__A1 (.DIODE(_02883_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11304__S (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA__11305__A1 (.DIODE(net593));
 sky130_fd_sc_hd__diode_2 ANTENNA__11305__B2 (.DIODE(net610));
 sky130_fd_sc_hd__diode_2 ANTENNA__11306__A1 (.DIODE(net591));
 sky130_fd_sc_hd__diode_2 ANTENNA__11307__B1 (.DIODE(_02885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11308__A0 (.DIODE(net364));
 sky130_fd_sc_hd__diode_2 ANTENNA__11308__A1 (.DIODE(_02886_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11308__S (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA__11309__B2 (.DIODE(net610));
 sky130_fd_sc_hd__diode_2 ANTENNA__11310__A1 (.DIODE(net591));
 sky130_fd_sc_hd__diode_2 ANTENNA__11311__B1 (.DIODE(_02888_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11312__A0 (.DIODE(net360));
 sky130_fd_sc_hd__diode_2 ANTENNA__11312__S (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA__11313__B2 (.DIODE(net610));
 sky130_fd_sc_hd__diode_2 ANTENNA__11314__A1 (.DIODE(net591));
 sky130_fd_sc_hd__diode_2 ANTENNA__11315__B1 (.DIODE(_02891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11316__A0 (.DIODE(net355));
 sky130_fd_sc_hd__diode_2 ANTENNA__11316__A1 (.DIODE(_02892_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11316__S (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA__11317__A1 (.DIODE(net593));
 sky130_fd_sc_hd__diode_2 ANTENNA__11317__B2 (.DIODE(net610));
 sky130_fd_sc_hd__diode_2 ANTENNA__11318__A1 (.DIODE(net591));
 sky130_fd_sc_hd__diode_2 ANTENNA__11319__A1 (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__11319__B1 (.DIODE(_02894_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11320__A1 (.DIODE(_02895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11320__S (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA__11321__A1 (.DIODE(net593));
 sky130_fd_sc_hd__diode_2 ANTENNA__11321__B2 (.DIODE(net610));
 sky130_fd_sc_hd__diode_2 ANTENNA__11323__A1 (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__11323__B1 (.DIODE(_02897_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11324__A0 (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA__11324__A1 (.DIODE(_02898_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11324__S (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA__11325__A1 (.DIODE(net593));
 sky130_fd_sc_hd__diode_2 ANTENNA__11325__B2 (.DIODE(net611));
 sky130_fd_sc_hd__diode_2 ANTENNA__11327__B1 (.DIODE(_02900_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11328__A0 (.DIODE(net341));
 sky130_fd_sc_hd__diode_2 ANTENNA__11328__A1 (.DIODE(_02901_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11328__S (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA__11329__B2 (.DIODE(net611));
 sky130_fd_sc_hd__diode_2 ANTENNA__11331__B1 (.DIODE(_02903_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11332__A0 (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA__11332__A1 (.DIODE(_02904_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11332__S (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA__11333__B2 (.DIODE(net610));
 sky130_fd_sc_hd__diode_2 ANTENNA__11335__A1 (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__11335__A3 (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__11335__B1 (.DIODE(_02906_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11336__A0 (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA__11336__A1 (.DIODE(_02907_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11336__S (.DIODE(_02756_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11337__B2 (.DIODE(net610));
 sky130_fd_sc_hd__diode_2 ANTENNA__11339__A1 (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__11339__A3 (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__11339__B1 (.DIODE(_02909_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11340__A0 (.DIODE(net331));
 sky130_fd_sc_hd__diode_2 ANTENNA__11340__A1 (.DIODE(_02910_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11340__S (.DIODE(_02756_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11341__B2 (.DIODE(net610));
 sky130_fd_sc_hd__diode_2 ANTENNA__11343__A1 (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__11343__A3 (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__11343__B1 (.DIODE(_02912_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11344__A0 (.DIODE(net329));
 sky130_fd_sc_hd__diode_2 ANTENNA__11344__A1 (.DIODE(_02913_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11344__S (.DIODE(_02756_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11345__B2 (.DIODE(net611));
 sky130_fd_sc_hd__diode_2 ANTENNA__11347__A1 (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__11347__A3 (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__11347__B1 (.DIODE(_02915_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11348__A0 (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA__11348__A1 (.DIODE(_02916_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11348__S (.DIODE(_02756_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11349__B2 (.DIODE(net611));
 sky130_fd_sc_hd__diode_2 ANTENNA__11351__B1 (.DIODE(_02918_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11352__S (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA__11353__A1 (.DIODE(net587));
 sky130_fd_sc_hd__diode_2 ANTENNA__11353__A2 (.DIODE(net601));
 sky130_fd_sc_hd__diode_2 ANTENNA__11353__B1 (.DIODE(net646));
 sky130_fd_sc_hd__diode_2 ANTENNA__11355__A2 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA__11356__A1 (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA__11356__S (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__11358__A2 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA__11359__A1 (.DIODE(net318));
 sky130_fd_sc_hd__diode_2 ANTENNA__11359__S (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__11360__A1 (.DIODE(net587));
 sky130_fd_sc_hd__diode_2 ANTENNA__11361__A2 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA__11362__A1 (.DIODE(net313));
 sky130_fd_sc_hd__diode_2 ANTENNA__11362__S (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__11364__A2 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA__11365__A1 (.DIODE(net309));
 sky130_fd_sc_hd__diode_2 ANTENNA__11365__S (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__11367__A2 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA__11368__A1 (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA__11368__S (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__11370__A2 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA__11371__A1 (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 ANTENNA__11371__S (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__11373__A2 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA__11374__A1 (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA__11374__S (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__11375__A1 (.DIODE(net586));
 sky130_fd_sc_hd__diode_2 ANTENNA__11376__A2 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA__11377__A1 (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA__11377__S (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__11379__A2 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA__11380__A1 (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA__11380__S (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__11382__A2 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA__11383__A1 (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA__11383__S (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__11385__A2 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA__11386__A1 (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__11386__S (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__11388__A2 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA__11389__A1 (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA__11389__S (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__11391__A2 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA__11392__A1 (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA__11392__S (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__11395__A1 (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__11395__S (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__11396__A1 (.DIODE(net587));
 sky130_fd_sc_hd__diode_2 ANTENNA__11396__B1 (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__11398__A1 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__11398__S (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__11401__A1 (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__11401__S (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__11404__A0 (.DIODE(_02954_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11404__A1 (.DIODE(net630));
 sky130_fd_sc_hd__diode_2 ANTENNA__11404__S (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__11405__A1 (.DIODE(net586));
 sky130_fd_sc_hd__diode_2 ANTENNA__11405__B1 (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__11407__A0 (.DIODE(_02956_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11407__A1 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__11407__S (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__11408__A1 (.DIODE(net586));
 sky130_fd_sc_hd__diode_2 ANTENNA__11410__A0 (.DIODE(_02958_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11410__A1 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__11410__S (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__11411__A1 (.DIODE(net586));
 sky130_fd_sc_hd__diode_2 ANTENNA__11413__A0 (.DIODE(_02960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11413__A1 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__11413__S (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__11414__A1 (.DIODE(net586));
 sky130_fd_sc_hd__diode_2 ANTENNA__11416__A0 (.DIODE(_02962_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11416__A1 (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA__11416__S (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__11417__A1 (.DIODE(net586));
 sky130_fd_sc_hd__diode_2 ANTENNA__11419__A0 (.DIODE(_02964_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11419__A1 (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA__11419__S (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__11420__A1 (.DIODE(net586));
 sky130_fd_sc_hd__diode_2 ANTENNA__11420__B1 (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__11422__A0 (.DIODE(_02966_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11422__A1 (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__11422__S (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__11423__A1 (.DIODE(net587));
 sky130_fd_sc_hd__diode_2 ANTENNA__11424__A2 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA__11425__A0 (.DIODE(_02968_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11425__A1 (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA__11425__S (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__11426__A1 (.DIODE(net586));
 sky130_fd_sc_hd__diode_2 ANTENNA__11428__A0 (.DIODE(_02970_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11428__A1 (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA__11428__S (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__11429__A1 (.DIODE(net586));
 sky130_fd_sc_hd__diode_2 ANTENNA__11431__A0 (.DIODE(_02972_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11431__A1 (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__11431__S (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__11432__A1 (.DIODE(net586));
 sky130_fd_sc_hd__diode_2 ANTENNA__11434__A0 (.DIODE(_02974_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11434__A1 (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__11434__S (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__11435__A1 (.DIODE(net586));
 sky130_fd_sc_hd__diode_2 ANTENNA__11437__A0 (.DIODE(_02976_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11437__A1 (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__11437__S (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__11438__A1 (.DIODE(net586));
 sky130_fd_sc_hd__diode_2 ANTENNA__11440__A0 (.DIODE(_02978_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11440__A1 (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__11440__S (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__11441__A1 (.DIODE(net586));
 sky130_fd_sc_hd__diode_2 ANTENNA__11441__B1 (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__11443__A0 (.DIODE(_02980_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11443__S (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__11444__A1 (.DIODE(net586));
 sky130_fd_sc_hd__diode_2 ANTENNA__11445__A2 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA__11446__A0 (.DIODE(_02982_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11446__S (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__11447__A1 (.DIODE(net586));
 sky130_fd_sc_hd__diode_2 ANTENNA__11448__A2 (.DIODE(_02755_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11449__A0 (.DIODE(_02984_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11449__A1 (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__11449__S (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__11450__A1 (.DIODE(net607));
 sky130_fd_sc_hd__diode_2 ANTENNA__11450__B2 (.DIODE(net601));
 sky130_fd_sc_hd__diode_2 ANTENNA__11451__A1 (.DIODE(net592));
 sky130_fd_sc_hd__diode_2 ANTENNA__11452__A1 (.DIODE(net625));
 sky130_fd_sc_hd__diode_2 ANTENNA__11452__S (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__11453__A1 (.DIODE(\state[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11453__B2 (.DIODE(net601));
 sky130_fd_sc_hd__diode_2 ANTENNA__11454__A1 (.DIODE(net587));
 sky130_fd_sc_hd__diode_2 ANTENNA__11455__A1 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__11455__S (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__11456__A1 (.DIODE(net607));
 sky130_fd_sc_hd__diode_2 ANTENNA__11456__B2 (.DIODE(net601));
 sky130_fd_sc_hd__diode_2 ANTENNA__11457__A1 (.DIODE(net587));
 sky130_fd_sc_hd__diode_2 ANTENNA__11458__A1 (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__11458__S (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__11459__A1 (.DIODE(net607));
 sky130_fd_sc_hd__diode_2 ANTENNA__11459__B2 (.DIODE(net606));
 sky130_fd_sc_hd__diode_2 ANTENNA__11460__A1 (.DIODE(net587));
 sky130_fd_sc_hd__diode_2 ANTENNA__11461__A1 (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__11461__S (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__11462__A1 (.DIODE(net607));
 sky130_fd_sc_hd__diode_2 ANTENNA__11462__B2 (.DIODE(net601));
 sky130_fd_sc_hd__diode_2 ANTENNA__11463__A1 (.DIODE(net587));
 sky130_fd_sc_hd__diode_2 ANTENNA__11464__A1 (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__11464__S (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__11465__A1 (.DIODE(net607));
 sky130_fd_sc_hd__diode_2 ANTENNA__11465__B2 (.DIODE(net601));
 sky130_fd_sc_hd__diode_2 ANTENNA__11466__A1 (.DIODE(net587));
 sky130_fd_sc_hd__diode_2 ANTENNA__11467__A1 (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__11467__S (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__11468__A1 (.DIODE(net607));
 sky130_fd_sc_hd__diode_2 ANTENNA__11468__B2 (.DIODE(net601));
 sky130_fd_sc_hd__diode_2 ANTENNA__11469__A1 (.DIODE(net588));
 sky130_fd_sc_hd__diode_2 ANTENNA__11470__A1 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__11470__S (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__11471__A1 (.DIODE(net607));
 sky130_fd_sc_hd__diode_2 ANTENNA__11471__B2 (.DIODE(net601));
 sky130_fd_sc_hd__diode_2 ANTENNA__11472__A1 (.DIODE(net588));
 sky130_fd_sc_hd__diode_2 ANTENNA__11473__A1 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__11473__S (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__11474__B2 (.DIODE(net602));
 sky130_fd_sc_hd__diode_2 ANTENNA__11475__A1 (.DIODE(net588));
 sky130_fd_sc_hd__diode_2 ANTENNA__11475__B2 (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__11476__A1 (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__11476__S (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__11477__B2 (.DIODE(net602));
 sky130_fd_sc_hd__diode_2 ANTENNA__11478__A1 (.DIODE(net588));
 sky130_fd_sc_hd__diode_2 ANTENNA__11478__B2 (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__11479__A1 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__11479__S (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__11480__B2 (.DIODE(net602));
 sky130_fd_sc_hd__diode_2 ANTENNA__11481__A1 (.DIODE(net588));
 sky130_fd_sc_hd__diode_2 ANTENNA__11481__B2 (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__11482__A1 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__11482__S (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__11483__B2 (.DIODE(net602));
 sky130_fd_sc_hd__diode_2 ANTENNA__11484__A1 (.DIODE(net588));
 sky130_fd_sc_hd__diode_2 ANTENNA__11484__B2 (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__11485__A1 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__11485__S (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__11486__B2 (.DIODE(net602));
 sky130_fd_sc_hd__diode_2 ANTENNA__11487__B2 (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__11488__A1 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__11488__S (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__11489__B2 (.DIODE(net602));
 sky130_fd_sc_hd__diode_2 ANTENNA__11490__B2 (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__11491__A1 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__11491__S (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__11492__B2 (.DIODE(net602));
 sky130_fd_sc_hd__diode_2 ANTENNA__11493__B2 (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__11494__A1 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__11494__S (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__11495__B2 (.DIODE(net602));
 sky130_fd_sc_hd__diode_2 ANTENNA__11496__A1 (.DIODE(net588));
 sky130_fd_sc_hd__diode_2 ANTENNA__11496__B2 (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__11497__A1 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__11497__S (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__11499__A1 (.DIODE(net588));
 sky130_fd_sc_hd__diode_2 ANTENNA__11499__B2 (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__11500__A1 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__11500__S (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__11501__B2 (.DIODE(net602));
 sky130_fd_sc_hd__diode_2 ANTENNA__11502__A1 (.DIODE(net588));
 sky130_fd_sc_hd__diode_2 ANTENNA__11502__B2 (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__11503__A1 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__11503__S (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__11505__A1 (.DIODE(net591));
 sky130_fd_sc_hd__diode_2 ANTENNA__11505__B2 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__11506__A1 (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__11506__S (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__11508__A1 (.DIODE(net591));
 sky130_fd_sc_hd__diode_2 ANTENNA__11508__B2 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__11509__A1 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__11509__S (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__11510__A1 (.DIODE(net610));
 sky130_fd_sc_hd__diode_2 ANTENNA__11511__A1 (.DIODE(net591));
 sky130_fd_sc_hd__diode_2 ANTENNA__11511__B2 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__11512__A1 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__11512__S (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__11513__A1 (.DIODE(net610));
 sky130_fd_sc_hd__diode_2 ANTENNA__11514__A1 (.DIODE(net591));
 sky130_fd_sc_hd__diode_2 ANTENNA__11514__B2 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__11515__A1 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__11515__S (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__11516__A1 (.DIODE(net610));
 sky130_fd_sc_hd__diode_2 ANTENNA__11517__A1 (.DIODE(net591));
 sky130_fd_sc_hd__diode_2 ANTENNA__11517__B2 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__11518__A1 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__11518__S (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__11519__A1 (.DIODE(net610));
 sky130_fd_sc_hd__diode_2 ANTENNA__11520__A1 (.DIODE(net591));
 sky130_fd_sc_hd__diode_2 ANTENNA__11520__B2 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__11521__A1 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__11521__S (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__11522__A1 (.DIODE(net610));
 sky130_fd_sc_hd__diode_2 ANTENNA__11523__B2 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__11524__A1 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__11524__S (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__11525__A1 (.DIODE(net611));
 sky130_fd_sc_hd__diode_2 ANTENNA__11526__B2 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__11527__A1 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__11527__S (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__11528__A1 (.DIODE(net610));
 sky130_fd_sc_hd__diode_2 ANTENNA__11529__B2 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__11530__A1 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__11530__S (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__11531__A1 (.DIODE(net611));
 sky130_fd_sc_hd__diode_2 ANTENNA__11532__B2 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__11533__A1 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__11533__S (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__11534__A1 (.DIODE(net611));
 sky130_fd_sc_hd__diode_2 ANTENNA__11535__B2 (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__11536__A1 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__11536__S (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__11537__A1 (.DIODE(net611));
 sky130_fd_sc_hd__diode_2 ANTENNA__11538__B2 (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__11539__A1 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__11539__S (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__11540__A1 (.DIODE(net611));
 sky130_fd_sc_hd__diode_2 ANTENNA__11541__B2 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__11542__A1 (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA__11542__S (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__11543__A1 (.DIODE(net611));
 sky130_fd_sc_hd__diode_2 ANTENNA__11544__B2 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__11545__A1 (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__11545__S (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__11546__A (.DIODE(net599));
 sky130_fd_sc_hd__diode_2 ANTENNA__11546__B (.DIODE(_02822_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11547__A (.DIODE(net599));
 sky130_fd_sc_hd__diode_2 ANTENNA__11547__B (.DIODE(_02822_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11548__A (.DIODE(net592));
 sky130_fd_sc_hd__diode_2 ANTENNA__11549__A (.DIODE(net592));
 sky130_fd_sc_hd__diode_2 ANTENNA__11550__A (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__11550__B (.DIODE(_03052_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11551__A (.DIODE(_03049_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11551__B (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__11552__A1 (.DIODE(net595));
 sky130_fd_sc_hd__diode_2 ANTENNA__11552__B1 (.DIODE(net645));
 sky130_fd_sc_hd__diode_2 ANTENNA__11553__A1 (.DIODE(net595));
 sky130_fd_sc_hd__diode_2 ANTENNA__11553__B1 (.DIODE(net645));
 sky130_fd_sc_hd__diode_2 ANTENNA__11554__B (.DIODE(_02822_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11555__B (.DIODE(_02822_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11556__B (.DIODE(net431));
 sky130_fd_sc_hd__diode_2 ANTENNA__11556__C (.DIODE(net540));
 sky130_fd_sc_hd__diode_2 ANTENNA__11557__C (.DIODE(net535));
 sky130_fd_sc_hd__diode_2 ANTENNA__11557__D (.DIODE(net540));
 sky130_fd_sc_hd__diode_2 ANTENNA__11558__A (.DIODE(net426));
 sky130_fd_sc_hd__diode_2 ANTENNA__11558__B (.DIODE(net544));
 sky130_fd_sc_hd__diode_2 ANTENNA__11559__A2 (.DIODE(net535));
 sky130_fd_sc_hd__diode_2 ANTENNA__11559__B1 (.DIODE(net540));
 sky130_fd_sc_hd__diode_2 ANTENNA__11561__A1 (.DIODE(net426));
 sky130_fd_sc_hd__diode_2 ANTENNA__11561__A2 (.DIODE(net544));
 sky130_fd_sc_hd__diode_2 ANTENNA__11562__A (.DIODE(net413));
 sky130_fd_sc_hd__diode_2 ANTENNA__11562__B (.DIODE(net552));
 sky130_fd_sc_hd__diode_2 ANTENNA__11563__A1 (.DIODE(net421));
 sky130_fd_sc_hd__diode_2 ANTENNA__11563__A2 (.DIODE(net545));
 sky130_fd_sc_hd__diode_2 ANTENNA__11563__B1 (.DIODE(net548));
 sky130_fd_sc_hd__diode_2 ANTENNA__11563__B2 (.DIODE(net417));
 sky130_fd_sc_hd__diode_2 ANTENNA__11564__A (.DIODE(net421));
 sky130_fd_sc_hd__diode_2 ANTENNA__11564__B (.DIODE(net417));
 sky130_fd_sc_hd__diode_2 ANTENNA__11564__C (.DIODE(net548));
 sky130_fd_sc_hd__diode_2 ANTENNA__11565__A1 (.DIODE(net545));
 sky130_fd_sc_hd__diode_2 ANTENNA__11568__A (.DIODE(net421));
 sky130_fd_sc_hd__diode_2 ANTENNA__11568__B (.DIODE(net417));
 sky130_fd_sc_hd__diode_2 ANTENNA__11568__C (.DIODE(net548));
 sky130_fd_sc_hd__diode_2 ANTENNA__11568__D (.DIODE(net552));
 sky130_fd_sc_hd__diode_2 ANTENNA__11569__A (.DIODE(net413));
 sky130_fd_sc_hd__diode_2 ANTENNA__11569__B (.DIODE(net558));
 sky130_fd_sc_hd__diode_2 ANTENNA__11570__A1 (.DIODE(net421));
 sky130_fd_sc_hd__diode_2 ANTENNA__11570__A2 (.DIODE(net548));
 sky130_fd_sc_hd__diode_2 ANTENNA__11570__B1 (.DIODE(net552));
 sky130_fd_sc_hd__diode_2 ANTENNA__11570__B2 (.DIODE(net417));
 sky130_fd_sc_hd__diode_2 ANTENNA__11572__A1 (.DIODE(net413));
 sky130_fd_sc_hd__diode_2 ANTENNA__11572__A2 (.DIODE(net558));
 sky130_fd_sc_hd__diode_2 ANTENNA__11575__A (.DIODE(net400));
 sky130_fd_sc_hd__diode_2 ANTENNA__11575__B (.DIODE(net564));
 sky130_fd_sc_hd__diode_2 ANTENNA__11576__A1 (.DIODE(net412));
 sky130_fd_sc_hd__diode_2 ANTENNA__11576__A2 (.DIODE(net552));
 sky130_fd_sc_hd__diode_2 ANTENNA__11576__B1 (.DIODE(net560));
 sky130_fd_sc_hd__diode_2 ANTENNA__11576__B2 (.DIODE(net405));
 sky130_fd_sc_hd__diode_2 ANTENNA__11577__A (.DIODE(net408));
 sky130_fd_sc_hd__diode_2 ANTENNA__11577__B (.DIODE(net404));
 sky130_fd_sc_hd__diode_2 ANTENNA__11577__C (.DIODE(net560));
 sky130_fd_sc_hd__diode_2 ANTENNA__11578__A1 (.DIODE(net552));
 sky130_fd_sc_hd__diode_2 ANTENNA__11580__A (.DIODE(net408));
 sky130_fd_sc_hd__diode_2 ANTENNA__11580__B (.DIODE(net404));
 sky130_fd_sc_hd__diode_2 ANTENNA__11580__C (.DIODE(net560));
 sky130_fd_sc_hd__diode_2 ANTENNA__11580__D (.DIODE(net564));
 sky130_fd_sc_hd__diode_2 ANTENNA__11581__A (.DIODE(net400));
 sky130_fd_sc_hd__diode_2 ANTENNA__11581__B (.DIODE(net567));
 sky130_fd_sc_hd__diode_2 ANTENNA__11582__A1 (.DIODE(net408));
 sky130_fd_sc_hd__diode_2 ANTENNA__11582__A2 (.DIODE(net560));
 sky130_fd_sc_hd__diode_2 ANTENNA__11582__B1 (.DIODE(net564));
 sky130_fd_sc_hd__diode_2 ANTENNA__11582__B2 (.DIODE(net404));
 sky130_fd_sc_hd__diode_2 ANTENNA__11584__A1 (.DIODE(net400));
 sky130_fd_sc_hd__diode_2 ANTENNA__11584__A2 (.DIODE(net567));
 sky130_fd_sc_hd__diode_2 ANTENNA__11586__A1 (.DIODE(net396));
 sky130_fd_sc_hd__diode_2 ANTENNA__11586__A2 (.DIODE(net567));
 sky130_fd_sc_hd__diode_2 ANTENNA__11586__B1 (.DIODE(net572));
 sky130_fd_sc_hd__diode_2 ANTENNA__11586__B2 (.DIODE(net390));
 sky130_fd_sc_hd__diode_2 ANTENNA__11587__A (.DIODE(net396));
 sky130_fd_sc_hd__diode_2 ANTENNA__11587__B (.DIODE(net390));
 sky130_fd_sc_hd__diode_2 ANTENNA__11587__C (.DIODE(net567));
 sky130_fd_sc_hd__diode_2 ANTENNA__11587__D (.DIODE(net575));
 sky130_fd_sc_hd__diode_2 ANTENNA__11589__A (.DIODE(net386));
 sky130_fd_sc_hd__diode_2 ANTENNA__11589__B (.DIODE(net577));
 sky130_fd_sc_hd__diode_2 ANTENNA__11590__A1 (.DIODE(net386));
 sky130_fd_sc_hd__diode_2 ANTENNA__11590__A2 (.DIODE(net577));
 sky130_fd_sc_hd__diode_2 ANTENNA__11596__A (.DIODE(net408));
 sky130_fd_sc_hd__diode_2 ANTENNA__11596__B (.DIODE(net404));
 sky130_fd_sc_hd__diode_2 ANTENNA__11596__C (.DIODE(net564));
 sky130_fd_sc_hd__diode_2 ANTENNA__11596__D (.DIODE(net567));
 sky130_fd_sc_hd__diode_2 ANTENNA__11597__A (.DIODE(net400));
 sky130_fd_sc_hd__diode_2 ANTENNA__11597__B (.DIODE(net572));
 sky130_fd_sc_hd__diode_2 ANTENNA__11598__A1 (.DIODE(net408));
 sky130_fd_sc_hd__diode_2 ANTENNA__11598__A2 (.DIODE(net564));
 sky130_fd_sc_hd__diode_2 ANTENNA__11598__B1 (.DIODE(net567));
 sky130_fd_sc_hd__diode_2 ANTENNA__11598__B2 (.DIODE(net404));
 sky130_fd_sc_hd__diode_2 ANTENNA__11600__A1 (.DIODE(net400));
 sky130_fd_sc_hd__diode_2 ANTENNA__11600__A2 (.DIODE(net572));
 sky130_fd_sc_hd__diode_2 ANTENNA__11603__A1 (.DIODE(net396));
 sky130_fd_sc_hd__diode_2 ANTENNA__11603__A2 (.DIODE(net572));
 sky130_fd_sc_hd__diode_2 ANTENNA__11603__B1 (.DIODE(net577));
 sky130_fd_sc_hd__diode_2 ANTENNA__11603__B2 (.DIODE(net390));
 sky130_fd_sc_hd__diode_2 ANTENNA__11604__A (.DIODE(net396));
 sky130_fd_sc_hd__diode_2 ANTENNA__11604__B (.DIODE(net390));
 sky130_fd_sc_hd__diode_2 ANTENNA__11604__C (.DIODE(net575));
 sky130_fd_sc_hd__diode_2 ANTENNA__11604__D (.DIODE(net577));
 sky130_fd_sc_hd__diode_2 ANTENNA__11606__A (.DIODE(net386));
 sky130_fd_sc_hd__diode_2 ANTENNA__11606__B (.DIODE(net581));
 sky130_fd_sc_hd__diode_2 ANTENNA__11607__A1 (.DIODE(net386));
 sky130_fd_sc_hd__diode_2 ANTENNA__11607__A2 (.DIODE(net581));
 sky130_fd_sc_hd__diode_2 ANTENNA__11613__A (.DIODE(net381));
 sky130_fd_sc_hd__diode_2 ANTENNA__11613__B (.DIODE(net581));
 sky130_fd_sc_hd__diode_2 ANTENNA__11615__A1 (.DIODE(net577));
 sky130_fd_sc_hd__diode_2 ANTENNA__11615__A2 (.DIODE(net381));
 sky130_fd_sc_hd__diode_2 ANTENNA__11615__B1 (.DIODE(net375));
 sky130_fd_sc_hd__diode_2 ANTENNA__11615__B2 (.DIODE(net584));
 sky130_fd_sc_hd__diode_2 ANTENNA__11616__A (.DIODE(net577));
 sky130_fd_sc_hd__diode_2 ANTENNA__11616__B (.DIODE(net381));
 sky130_fd_sc_hd__diode_2 ANTENNA__11616__C (.DIODE(net375));
 sky130_fd_sc_hd__diode_2 ANTENNA__11616__D (.DIODE(net581));
 sky130_fd_sc_hd__diode_2 ANTENNA__11617__A (.DIODE(net577));
 sky130_fd_sc_hd__diode_2 ANTENNA__11617__B (.DIODE(net381));
 sky130_fd_sc_hd__diode_2 ANTENNA__11617__C (.DIODE(net375));
 sky130_fd_sc_hd__diode_2 ANTENNA__11617__D (.DIODE(net582));
 sky130_fd_sc_hd__diode_2 ANTENNA__11625__D (.DIODE(net535));
 sky130_fd_sc_hd__diode_2 ANTENNA__11626__B1 (.DIODE(net536));
 sky130_fd_sc_hd__diode_2 ANTENNA__11627__C (.DIODE(net426));
 sky130_fd_sc_hd__diode_2 ANTENNA__11627__D (.DIODE(net540));
 sky130_fd_sc_hd__diode_2 ANTENNA__11628__A1 (.DIODE(net421));
 sky130_fd_sc_hd__diode_2 ANTENNA__11628__A2 (.DIODE(net540));
 sky130_fd_sc_hd__diode_2 ANTENNA__11628__B1 (.DIODE(net544));
 sky130_fd_sc_hd__diode_2 ANTENNA__11628__B2 (.DIODE(net417));
 sky130_fd_sc_hd__diode_2 ANTENNA__11629__A (.DIODE(net421));
 sky130_fd_sc_hd__diode_2 ANTENNA__11629__B (.DIODE(net417));
 sky130_fd_sc_hd__diode_2 ANTENNA__11629__C (.DIODE(net540));
 sky130_fd_sc_hd__diode_2 ANTENNA__11629__D (.DIODE(net544));
 sky130_fd_sc_hd__diode_2 ANTENNA__11630__A (.DIODE(net413));
 sky130_fd_sc_hd__diode_2 ANTENNA__11630__B (.DIODE(net548));
 sky130_fd_sc_hd__diode_2 ANTENNA__11631__A1 (.DIODE(net413));
 sky130_fd_sc_hd__diode_2 ANTENNA__11631__A2 (.DIODE(net548));
 sky130_fd_sc_hd__diode_2 ANTENNA__11633__A1 (.DIODE(net413));
 sky130_fd_sc_hd__diode_2 ANTENNA__11633__A2 (.DIODE(net552));
 sky130_fd_sc_hd__diode_2 ANTENNA__11633__B2 (.DIODE(net545));
 sky130_fd_sc_hd__diode_2 ANTENNA__11637__A (.DIODE(net400));
 sky130_fd_sc_hd__diode_2 ANTENNA__11637__B (.DIODE(net557));
 sky130_fd_sc_hd__diode_2 ANTENNA__11638__A1 (.DIODE(net548));
 sky130_fd_sc_hd__diode_2 ANTENNA__11638__A2 (.DIODE(net408));
 sky130_fd_sc_hd__diode_2 ANTENNA__11638__B1 (.DIODE(net405));
 sky130_fd_sc_hd__diode_2 ANTENNA__11638__B2 (.DIODE(net552));
 sky130_fd_sc_hd__diode_2 ANTENNA__11639__A (.DIODE(net548));
 sky130_fd_sc_hd__diode_2 ANTENNA__11639__B (.DIODE(net408));
 sky130_fd_sc_hd__diode_2 ANTENNA__11639__C (.DIODE(net405));
 sky130_fd_sc_hd__diode_2 ANTENNA__11639__D (.DIODE(net552));
 sky130_fd_sc_hd__diode_2 ANTENNA__11642__A1 (.DIODE(net400));
 sky130_fd_sc_hd__diode_2 ANTENNA__11642__A2 (.DIODE(net564));
 sky130_fd_sc_hd__diode_2 ANTENNA__11642__B2 (.DIODE(net552));
 sky130_fd_sc_hd__diode_2 ANTENNA__11645__A (.DIODE(net386));
 sky130_fd_sc_hd__diode_2 ANTENNA__11645__B (.DIODE(net572));
 sky130_fd_sc_hd__diode_2 ANTENNA__11646__A1 (.DIODE(net396));
 sky130_fd_sc_hd__diode_2 ANTENNA__11646__A2 (.DIODE(net564));
 sky130_fd_sc_hd__diode_2 ANTENNA__11646__B1 (.DIODE(net567));
 sky130_fd_sc_hd__diode_2 ANTENNA__11646__B2 (.DIODE(net390));
 sky130_fd_sc_hd__diode_2 ANTENNA__11647__A (.DIODE(net396));
 sky130_fd_sc_hd__diode_2 ANTENNA__11647__B (.DIODE(net390));
 sky130_fd_sc_hd__diode_2 ANTENNA__11647__C (.DIODE(net564));
 sky130_fd_sc_hd__diode_2 ANTENNA__11647__D (.DIODE(net567));
 sky130_fd_sc_hd__diode_2 ANTENNA__11657__A1 (.DIODE(net386));
 sky130_fd_sc_hd__diode_2 ANTENNA__11657__A2 (.DIODE(net575));
 sky130_fd_sc_hd__diode_2 ANTENNA__11658__A (.DIODE(net371));
 sky130_fd_sc_hd__diode_2 ANTENNA__11658__B (.DIODE(net581));
 sky130_fd_sc_hd__diode_2 ANTENNA__11659__A (.DIODE(net572));
 sky130_fd_sc_hd__diode_2 ANTENNA__11659__B (.DIODE(net580));
 sky130_fd_sc_hd__diode_2 ANTENNA__11659__C (.DIODE(net381));
 sky130_fd_sc_hd__diode_2 ANTENNA__11659__D (.DIODE(net375));
 sky130_fd_sc_hd__diode_2 ANTENNA__11660__A1 (.DIODE(net572));
 sky130_fd_sc_hd__diode_2 ANTENNA__11660__A2 (.DIODE(net381));
 sky130_fd_sc_hd__diode_2 ANTENNA__11660__B1 (.DIODE(net375));
 sky130_fd_sc_hd__diode_2 ANTENNA__11660__B2 (.DIODE(net580));
 sky130_fd_sc_hd__diode_2 ANTENNA__11673__C (.DIODE(net525));
 sky130_fd_sc_hd__diode_2 ANTENNA__11674__A (.DIODE(net426));
 sky130_fd_sc_hd__diode_2 ANTENNA__11674__B (.DIODE(net535));
 sky130_fd_sc_hd__diode_2 ANTENNA__11675__A2 (.DIODE(net525));
 sky130_fd_sc_hd__diode_2 ANTENNA__11677__A1 (.DIODE(net426));
 sky130_fd_sc_hd__diode_2 ANTENNA__11677__A2 (.DIODE(net535));
 sky130_fd_sc_hd__diode_2 ANTENNA__11678__A1 (.DIODE(net421));
 sky130_fd_sc_hd__diode_2 ANTENNA__11678__A2 (.DIODE(net536));
 sky130_fd_sc_hd__diode_2 ANTENNA__11678__B1 (.DIODE(net541));
 sky130_fd_sc_hd__diode_2 ANTENNA__11678__B2 (.DIODE(net417));
 sky130_fd_sc_hd__diode_2 ANTENNA__11679__A (.DIODE(net421));
 sky130_fd_sc_hd__diode_2 ANTENNA__11679__B (.DIODE(net417));
 sky130_fd_sc_hd__diode_2 ANTENNA__11679__C (.DIODE(net536));
 sky130_fd_sc_hd__diode_2 ANTENNA__11679__D (.DIODE(net540));
 sky130_fd_sc_hd__diode_2 ANTENNA__11680__A (.DIODE(net413));
 sky130_fd_sc_hd__diode_2 ANTENNA__11680__B (.DIODE(net545));
 sky130_fd_sc_hd__diode_2 ANTENNA__11681__A1 (.DIODE(net413));
 sky130_fd_sc_hd__diode_2 ANTENNA__11681__A2 (.DIODE(net545));
 sky130_fd_sc_hd__diode_2 ANTENNA__11687__A (.DIODE(net386));
 sky130_fd_sc_hd__diode_2 ANTENNA__11687__B (.DIODE(net567));
 sky130_fd_sc_hd__diode_2 ANTENNA__11688__A (.DIODE(net560));
 sky130_fd_sc_hd__diode_2 ANTENNA__11688__B (.DIODE(net396));
 sky130_fd_sc_hd__diode_2 ANTENNA__11688__C (.DIODE(net390));
 sky130_fd_sc_hd__diode_2 ANTENNA__11688__D (.DIODE(net564));
 sky130_fd_sc_hd__diode_2 ANTENNA__11689__A1 (.DIODE(net560));
 sky130_fd_sc_hd__diode_2 ANTENNA__11689__A2 (.DIODE(net396));
 sky130_fd_sc_hd__diode_2 ANTENNA__11689__B1 (.DIODE(net390));
 sky130_fd_sc_hd__diode_2 ANTENNA__11689__B2 (.DIODE(net564));
 sky130_fd_sc_hd__diode_2 ANTENNA__11692__A (.DIODE(net545));
 sky130_fd_sc_hd__diode_2 ANTENNA__11692__B (.DIODE(net548));
 sky130_fd_sc_hd__diode_2 ANTENNA__11692__C (.DIODE(net408));
 sky130_fd_sc_hd__diode_2 ANTENNA__11692__D (.DIODE(net404));
 sky130_fd_sc_hd__diode_2 ANTENNA__11693__A1 (.DIODE(net545));
 sky130_fd_sc_hd__diode_2 ANTENNA__11693__A2 (.DIODE(net408));
 sky130_fd_sc_hd__diode_2 ANTENNA__11693__B1 (.DIODE(net404));
 sky130_fd_sc_hd__diode_2 ANTENNA__11693__B2 (.DIODE(net548));
 sky130_fd_sc_hd__diode_2 ANTENNA__11694__A (.DIODE(net400));
 sky130_fd_sc_hd__diode_2 ANTENNA__11694__B (.DIODE(net552));
 sky130_fd_sc_hd__diode_2 ANTENNA__11695__A1 (.DIODE(net400));
 sky130_fd_sc_hd__diode_2 ANTENNA__11695__A2 (.DIODE(net552));
 sky130_fd_sc_hd__diode_2 ANTENNA__11706__A (.DIODE(net436));
 sky130_fd_sc_hd__diode_2 ANTENNA__11706__C (.DIODE(net520));
 sky130_fd_sc_hd__diode_2 ANTENNA__11706__D (.DIODE(net525));
 sky130_fd_sc_hd__diode_2 ANTENNA__11707__A1 (.DIODE(net436));
 sky130_fd_sc_hd__diode_2 ANTENNA__11707__A2 (.DIODE(net520));
 sky130_fd_sc_hd__diode_2 ANTENNA__11707__B1 (.DIODE(net525));
 sky130_fd_sc_hd__diode_2 ANTENNA__11708__C (.DIODE(net426));
 sky130_fd_sc_hd__diode_2 ANTENNA__11710__A (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA__11710__B (.DIODE(net541));
 sky130_fd_sc_hd__diode_2 ANTENNA__11711__B (.DIODE(net422));
 sky130_fd_sc_hd__diode_2 ANTENNA__11711__C (.DIODE(net418));
 sky130_fd_sc_hd__diode_2 ANTENNA__11711__D (.DIODE(net536));
 sky130_fd_sc_hd__diode_2 ANTENNA__11712__A2 (.DIODE(net422));
 sky130_fd_sc_hd__diode_2 ANTENNA__11712__B1 (.DIODE(net418));
 sky130_fd_sc_hd__diode_2 ANTENNA__11712__B2 (.DIODE(net536));
 sky130_fd_sc_hd__diode_2 ANTENNA__11719__A (.DIODE(net427));
 sky130_fd_sc_hd__diode_2 ANTENNA__11719__B (.DIODE(net525));
 sky130_fd_sc_hd__diode_2 ANTENNA__11720__A1 (.DIODE(net516));
 sky130_fd_sc_hd__diode_2 ANTENNA__11720__A2 (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA__11720__B1 (.DIODE(net432));
 sky130_fd_sc_hd__diode_2 ANTENNA__11720__B2 (.DIODE(net520));
 sky130_fd_sc_hd__diode_2 ANTENNA__11721__A (.DIODE(net515));
 sky130_fd_sc_hd__diode_2 ANTENNA__11721__C (.DIODE(net432));
 sky130_fd_sc_hd__diode_2 ANTENNA__11721__D (.DIODE(net520));
 sky130_fd_sc_hd__diode_2 ANTENNA__11724__A (.DIODE(net441));
 sky130_fd_sc_hd__diode_2 ANTENNA__11724__B (.DIODE(net511));
 sky130_fd_sc_hd__diode_2 ANTENNA__11725__B (.DIODE(net503));
 sky130_fd_sc_hd__diode_2 ANTENNA__11725__D (.DIODE(net507));
 sky130_fd_sc_hd__diode_2 ANTENNA__11726__A2 (.DIODE(net503));
 sky130_fd_sc_hd__diode_2 ANTENNA__11726__B2 (.DIODE(net507));
 sky130_fd_sc_hd__diode_2 ANTENNA__11729__C (.DIODE(net507));
 sky130_fd_sc_hd__diode_2 ANTENNA__11729__D (.DIODE(net511));
 sky130_fd_sc_hd__diode_2 ANTENNA__11730__A (.DIODE(net441));
 sky130_fd_sc_hd__diode_2 ANTENNA__11730__B (.DIODE(net515));
 sky130_fd_sc_hd__diode_2 ANTENNA__11731__A2 (.DIODE(net507));
 sky130_fd_sc_hd__diode_2 ANTENNA__11731__B1 (.DIODE(net511));
 sky130_fd_sc_hd__diode_2 ANTENNA__11738__C (.DIODE(net511));
 sky130_fd_sc_hd__diode_2 ANTENNA__11738__D (.DIODE(net515));
 sky130_fd_sc_hd__diode_2 ANTENNA__11739__A (.DIODE(net441));
 sky130_fd_sc_hd__diode_2 ANTENNA__11739__B (.DIODE(net520));
 sky130_fd_sc_hd__diode_2 ANTENNA__11740__A2 (.DIODE(net511));
 sky130_fd_sc_hd__diode_2 ANTENNA__11740__B1 (.DIODE(net515));
 sky130_fd_sc_hd__diode_2 ANTENNA__11746__A1_N (.DIODE(net427));
 sky130_fd_sc_hd__diode_2 ANTENNA__11755__C (.DIODE(net515));
 sky130_fd_sc_hd__diode_2 ANTENNA__11755__D (.DIODE(net520));
 sky130_fd_sc_hd__diode_2 ANTENNA__11756__A (.DIODE(net440));
 sky130_fd_sc_hd__diode_2 ANTENNA__11756__B (.DIODE(net525));
 sky130_fd_sc_hd__diode_2 ANTENNA__11757__A2 (.DIODE(net515));
 sky130_fd_sc_hd__diode_2 ANTENNA__11757__B1 (.DIODE(net520));
 sky130_fd_sc_hd__diode_2 ANTENNA__11778__C (.DIODE(net520));
 sky130_fd_sc_hd__diode_2 ANTENNA__11778__D (.DIODE(net525));
 sky130_fd_sc_hd__diode_2 ANTENNA__11779__A (.DIODE(net440));
 sky130_fd_sc_hd__diode_2 ANTENNA__11780__A2 (.DIODE(net520));
 sky130_fd_sc_hd__diode_2 ANTENNA__11780__B1 (.DIODE(net525));
 sky130_fd_sc_hd__diode_2 ANTENNA__11786__A1_N (.DIODE(net426));
 sky130_fd_sc_hd__diode_2 ANTENNA__11786__A2_N (.DIODE(net540));
 sky130_fd_sc_hd__diode_2 ANTENNA__11807__C (.DIODE(net525));
 sky130_fd_sc_hd__diode_2 ANTENNA__11808__A (.DIODE(net440));
 sky130_fd_sc_hd__diode_2 ANTENNA__11808__B (.DIODE(net535));
 sky130_fd_sc_hd__diode_2 ANTENNA__11809__A2 (.DIODE(net525));
 sky130_fd_sc_hd__diode_2 ANTENNA__11842__D (.DIODE(net535));
 sky130_fd_sc_hd__diode_2 ANTENNA__11843__A (.DIODE(net440));
 sky130_fd_sc_hd__diode_2 ANTENNA__11843__B (.DIODE(net540));
 sky130_fd_sc_hd__diode_2 ANTENNA__11844__B1 (.DIODE(net535));
 sky130_fd_sc_hd__diode_2 ANTENNA__11850__A (.DIODE(net426));
 sky130_fd_sc_hd__diode_2 ANTENNA__11850__B (.DIODE(net548));
 sky130_fd_sc_hd__diode_2 ANTENNA__11851__A1 (.DIODE(net436));
 sky130_fd_sc_hd__diode_2 ANTENNA__11851__A2 (.DIODE(net540));
 sky130_fd_sc_hd__diode_2 ANTENNA__11851__B1 (.DIODE(net544));
 sky130_fd_sc_hd__diode_2 ANTENNA__11851__B2 (.DIODE(net431));
 sky130_fd_sc_hd__diode_2 ANTENNA__11852__A1 (.DIODE(net544));
 sky130_fd_sc_hd__diode_2 ANTENNA__11859__A (.DIODE(net422));
 sky130_fd_sc_hd__diode_2 ANTENNA__11859__B (.DIODE(net418));
 sky130_fd_sc_hd__diode_2 ANTENNA__11859__C (.DIODE(net552));
 sky130_fd_sc_hd__diode_2 ANTENNA__11859__D (.DIODE(net558));
 sky130_fd_sc_hd__diode_2 ANTENNA__11860__A (.DIODE(net413));
 sky130_fd_sc_hd__diode_2 ANTENNA__11860__B (.DIODE(net565));
 sky130_fd_sc_hd__diode_2 ANTENNA__11861__A1 (.DIODE(net422));
 sky130_fd_sc_hd__diode_2 ANTENNA__11861__A2 (.DIODE(net552));
 sky130_fd_sc_hd__diode_2 ANTENNA__11861__B1 (.DIODE(net558));
 sky130_fd_sc_hd__diode_2 ANTENNA__11861__B2 (.DIODE(net418));
 sky130_fd_sc_hd__diode_2 ANTENNA__11863__A1 (.DIODE(net413));
 sky130_fd_sc_hd__diode_2 ANTENNA__11863__A2 (.DIODE(net565));
 sky130_fd_sc_hd__diode_2 ANTENNA__11864__A1 (.DIODE(net427));
 sky130_fd_sc_hd__diode_2 ANTENNA__11864__A2 (.DIODE(net548));
 sky130_fd_sc_hd__diode_2 ANTENNA__11864__B2 (.DIODE(net544));
 sky130_fd_sc_hd__diode_2 ANTENNA__11875__A (.DIODE(net408));
 sky130_fd_sc_hd__diode_2 ANTENNA__11875__B (.DIODE(net404));
 sky130_fd_sc_hd__diode_2 ANTENNA__11875__C (.DIODE(net567));
 sky130_fd_sc_hd__diode_2 ANTENNA__11875__D (.DIODE(net572));
 sky130_fd_sc_hd__diode_2 ANTENNA__11877__A1 (.DIODE(net408));
 sky130_fd_sc_hd__diode_2 ANTENNA__11877__A2 (.DIODE(net567));
 sky130_fd_sc_hd__diode_2 ANTENNA__11877__B1 (.DIODE(net572));
 sky130_fd_sc_hd__diode_2 ANTENNA__11877__B2 (.DIODE(net404));
 sky130_fd_sc_hd__diode_2 ANTENNA__11878__C (.DIODE(net400));
 sky130_fd_sc_hd__diode_2 ANTENNA__11878__D (.DIODE(net577));
 sky130_fd_sc_hd__diode_2 ANTENNA__11882__A1 (.DIODE(net396));
 sky130_fd_sc_hd__diode_2 ANTENNA__11882__A2 (.DIODE(net577));
 sky130_fd_sc_hd__diode_2 ANTENNA__11882__B1 (.DIODE(net581));
 sky130_fd_sc_hd__diode_2 ANTENNA__11882__B2 (.DIODE(net390));
 sky130_fd_sc_hd__diode_2 ANTENNA__11884__A (.DIODE(net396));
 sky130_fd_sc_hd__diode_2 ANTENNA__11884__B (.DIODE(net390));
 sky130_fd_sc_hd__diode_2 ANTENNA__11884__C (.DIODE(net577));
 sky130_fd_sc_hd__diode_2 ANTENNA__11884__D (.DIODE(net581));
 sky130_fd_sc_hd__diode_2 ANTENNA__11911__C (.DIODE(net535));
 sky130_fd_sc_hd__diode_2 ANTENNA__11911__D (.DIODE(net540));
 sky130_fd_sc_hd__diode_2 ANTENNA__11912__A (.DIODE(net440));
 sky130_fd_sc_hd__diode_2 ANTENNA__11912__B (.DIODE(net544));
 sky130_fd_sc_hd__diode_2 ANTENNA__11913__A2 (.DIODE(net535));
 sky130_fd_sc_hd__diode_2 ANTENNA__11913__B1 (.DIODE(net540));
 sky130_fd_sc_hd__diode_2 ANTENNA__11919__A (.DIODE(net427));
 sky130_fd_sc_hd__diode_2 ANTENNA__11919__B (.DIODE(net552));
 sky130_fd_sc_hd__diode_2 ANTENNA__11920__A2 (.DIODE(net544));
 sky130_fd_sc_hd__diode_2 ANTENNA__11920__B1 (.DIODE(net549));
 sky130_fd_sc_hd__diode_2 ANTENNA__11921__C (.DIODE(net544));
 sky130_fd_sc_hd__diode_2 ANTENNA__11921__D (.DIODE(net549));
 sky130_fd_sc_hd__diode_2 ANTENNA__11930__A (.DIODE(net422));
 sky130_fd_sc_hd__diode_2 ANTENNA__11930__B (.DIODE(net418));
 sky130_fd_sc_hd__diode_2 ANTENNA__11930__C (.DIODE(net558));
 sky130_fd_sc_hd__diode_2 ANTENNA__11930__D (.DIODE(net565));
 sky130_fd_sc_hd__diode_2 ANTENNA__11931__A (.DIODE(net413));
 sky130_fd_sc_hd__diode_2 ANTENNA__11931__B (.DIODE(net570));
 sky130_fd_sc_hd__diode_2 ANTENNA__11932__A1 (.DIODE(net422));
 sky130_fd_sc_hd__diode_2 ANTENNA__11932__A2 (.DIODE(net558));
 sky130_fd_sc_hd__diode_2 ANTENNA__11932__B1 (.DIODE(net561));
 sky130_fd_sc_hd__diode_2 ANTENNA__11932__B2 (.DIODE(net418));
 sky130_fd_sc_hd__diode_2 ANTENNA__11934__A1 (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA__11934__A2 (.DIODE(net566));
 sky130_fd_sc_hd__diode_2 ANTENNA__11947__A1 (.DIODE(net400));
 sky130_fd_sc_hd__diode_2 ANTENNA__11947__A2 (.DIODE(net577));
 sky130_fd_sc_hd__diode_2 ANTENNA__11949__A (.DIODE(net408));
 sky130_fd_sc_hd__diode_2 ANTENNA__11949__B (.DIODE(net404));
 sky130_fd_sc_hd__diode_2 ANTENNA__11949__C (.DIODE(net572));
 sky130_fd_sc_hd__diode_2 ANTENNA__11949__D (.DIODE(net577));
 sky130_fd_sc_hd__diode_2 ANTENNA__11951__A1 (.DIODE(net408));
 sky130_fd_sc_hd__diode_2 ANTENNA__11951__A2 (.DIODE(net572));
 sky130_fd_sc_hd__diode_2 ANTENNA__11951__B1 (.DIODE(net577));
 sky130_fd_sc_hd__diode_2 ANTENNA__11951__B2 (.DIODE(net404));
 sky130_fd_sc_hd__diode_2 ANTENNA__11952__A (.DIODE(net400));
 sky130_fd_sc_hd__diode_2 ANTENNA__11952__B (.DIODE(net581));
 sky130_fd_sc_hd__diode_2 ANTENNA__11955__A (.DIODE(net396));
 sky130_fd_sc_hd__diode_2 ANTENNA__11955__B (.DIODE(net581));
 sky130_fd_sc_hd__diode_2 ANTENNA__11983__C (.DIODE(net540));
 sky130_fd_sc_hd__diode_2 ANTENNA__11983__D (.DIODE(net544));
 sky130_fd_sc_hd__diode_2 ANTENNA__11984__A (.DIODE(net440));
 sky130_fd_sc_hd__diode_2 ANTENNA__11984__B (.DIODE(net549));
 sky130_fd_sc_hd__diode_2 ANTENNA__11985__A2 (.DIODE(net540));
 sky130_fd_sc_hd__diode_2 ANTENNA__11985__B1 (.DIODE(net544));
 sky130_fd_sc_hd__diode_2 ANTENNA__11990__A2 (.DIODE(net549));
 sky130_fd_sc_hd__diode_2 ANTENNA__11990__B1 (.DIODE(net553));
 sky130_fd_sc_hd__diode_2 ANTENNA__11991__C (.DIODE(net549));
 sky130_fd_sc_hd__diode_2 ANTENNA__11991__D (.DIODE(net553));
 sky130_fd_sc_hd__diode_2 ANTENNA__11993__A (.DIODE(net427));
 sky130_fd_sc_hd__diode_2 ANTENNA__11993__B (.DIODE(net557));
 sky130_fd_sc_hd__diode_2 ANTENNA__12004__A (.DIODE(net422));
 sky130_fd_sc_hd__diode_2 ANTENNA__12004__B (.DIODE(net417));
 sky130_fd_sc_hd__diode_2 ANTENNA__12004__C (.DIODE(net561));
 sky130_fd_sc_hd__diode_2 ANTENNA__12004__D (.DIODE(net570));
 sky130_fd_sc_hd__diode_2 ANTENNA__12005__A (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA__12005__B (.DIODE(net571));
 sky130_fd_sc_hd__diode_2 ANTENNA__12006__A1 (.DIODE(net422));
 sky130_fd_sc_hd__diode_2 ANTENNA__12006__A2 (.DIODE(net561));
 sky130_fd_sc_hd__diode_2 ANTENNA__12006__B1 (.DIODE(net570));
 sky130_fd_sc_hd__diode_2 ANTENNA__12006__B2 (.DIODE(net418));
 sky130_fd_sc_hd__diode_2 ANTENNA__12008__A1 (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA__12008__A2 (.DIODE(net575));
 sky130_fd_sc_hd__diode_2 ANTENNA__12018__A1 (.DIODE(net400));
 sky130_fd_sc_hd__diode_2 ANTENNA__12018__A2 (.DIODE(net581));
 sky130_fd_sc_hd__diode_2 ANTENNA__12020__A (.DIODE(net408));
 sky130_fd_sc_hd__diode_2 ANTENNA__12020__B (.DIODE(net404));
 sky130_fd_sc_hd__diode_2 ANTENNA__12020__C (.DIODE(net577));
 sky130_fd_sc_hd__diode_2 ANTENNA__12020__D (.DIODE(net581));
 sky130_fd_sc_hd__diode_2 ANTENNA__12037__C (.DIODE(net544));
 sky130_fd_sc_hd__diode_2 ANTENNA__12037__D (.DIODE(net549));
 sky130_fd_sc_hd__diode_2 ANTENNA__12038__A (.DIODE(net440));
 sky130_fd_sc_hd__diode_2 ANTENNA__12038__B (.DIODE(net553));
 sky130_fd_sc_hd__diode_2 ANTENNA__12039__A2 (.DIODE(net544));
 sky130_fd_sc_hd__diode_2 ANTENNA__12039__B1 (.DIODE(net549));
 sky130_fd_sc_hd__diode_2 ANTENNA__12044__C (.DIODE(net553));
 sky130_fd_sc_hd__diode_2 ANTENNA__12044__D (.DIODE(net557));
 sky130_fd_sc_hd__diode_2 ANTENNA__12045__A2 (.DIODE(net553));
 sky130_fd_sc_hd__diode_2 ANTENNA__12045__B1 (.DIODE(net557));
 sky130_fd_sc_hd__diode_2 ANTENNA__12047__A (.DIODE(net427));
 sky130_fd_sc_hd__diode_2 ANTENNA__12047__B (.DIODE(net561));
 sky130_fd_sc_hd__diode_2 ANTENNA__12054__A1 (.DIODE(net427));
 sky130_fd_sc_hd__diode_2 ANTENNA__12054__A2 (.DIODE(net561));
 sky130_fd_sc_hd__diode_2 ANTENNA__12058__A (.DIODE(net421));
 sky130_fd_sc_hd__diode_2 ANTENNA__12058__B (.DIODE(net417));
 sky130_fd_sc_hd__diode_2 ANTENNA__12058__C (.DIODE(net566));
 sky130_fd_sc_hd__diode_2 ANTENNA__12058__D (.DIODE(net571));
 sky130_fd_sc_hd__diode_2 ANTENNA__12059__A (.DIODE(net413));
 sky130_fd_sc_hd__diode_2 ANTENNA__12059__B (.DIODE(net576));
 sky130_fd_sc_hd__diode_2 ANTENNA__12060__A1 (.DIODE(net421));
 sky130_fd_sc_hd__diode_2 ANTENNA__12060__A2 (.DIODE(net566));
 sky130_fd_sc_hd__diode_2 ANTENNA__12060__B1 (.DIODE(net571));
 sky130_fd_sc_hd__diode_2 ANTENNA__12060__B2 (.DIODE(net417));
 sky130_fd_sc_hd__diode_2 ANTENNA__12062__A1 (.DIODE(net413));
 sky130_fd_sc_hd__diode_2 ANTENNA__12062__A2 (.DIODE(net576));
 sky130_fd_sc_hd__diode_2 ANTENNA__12088__C (.DIODE(net549));
 sky130_fd_sc_hd__diode_2 ANTENNA__12088__D (.DIODE(net553));
 sky130_fd_sc_hd__diode_2 ANTENNA__12089__A (.DIODE(net440));
 sky130_fd_sc_hd__diode_2 ANTENNA__12089__B (.DIODE(net557));
 sky130_fd_sc_hd__diode_2 ANTENNA__12090__A2 (.DIODE(net549));
 sky130_fd_sc_hd__diode_2 ANTENNA__12090__B1 (.DIODE(net553));
 sky130_fd_sc_hd__diode_2 ANTENNA__12094__C (.DIODE(net557));
 sky130_fd_sc_hd__diode_2 ANTENNA__12094__D (.DIODE(net561));
 sky130_fd_sc_hd__diode_2 ANTENNA__12095__A2 (.DIODE(net557));
 sky130_fd_sc_hd__diode_2 ANTENNA__12095__B1 (.DIODE(net561));
 sky130_fd_sc_hd__diode_2 ANTENNA__12097__A (.DIODE(net426));
 sky130_fd_sc_hd__diode_2 ANTENNA__12097__B (.DIODE(net566));
 sky130_fd_sc_hd__diode_2 ANTENNA__12103__A1 (.DIODE(net426));
 sky130_fd_sc_hd__diode_2 ANTENNA__12103__A2 (.DIODE(net566));
 sky130_fd_sc_hd__diode_2 ANTENNA__12107__A (.DIODE(net421));
 sky130_fd_sc_hd__diode_2 ANTENNA__12107__B (.DIODE(net417));
 sky130_fd_sc_hd__diode_2 ANTENNA__12107__C (.DIODE(net571));
 sky130_fd_sc_hd__diode_2 ANTENNA__12107__D (.DIODE(net576));
 sky130_fd_sc_hd__diode_2 ANTENNA__12108__A1 (.DIODE(net421));
 sky130_fd_sc_hd__diode_2 ANTENNA__12108__A2 (.DIODE(net571));
 sky130_fd_sc_hd__diode_2 ANTENNA__12108__B1 (.DIODE(net576));
 sky130_fd_sc_hd__diode_2 ANTENNA__12108__B2 (.DIODE(net417));
 sky130_fd_sc_hd__diode_2 ANTENNA__12109__C (.DIODE(net413));
 sky130_fd_sc_hd__diode_2 ANTENNA__12109__D (.DIODE(net582));
 sky130_fd_sc_hd__diode_2 ANTENNA__12117__A1 (.DIODE(net408));
 sky130_fd_sc_hd__diode_2 ANTENNA__12117__A2 (.DIODE(net577));
 sky130_fd_sc_hd__diode_2 ANTENNA__12117__B1 (.DIODE(net581));
 sky130_fd_sc_hd__diode_2 ANTENNA__12117__B2 (.DIODE(net404));
 sky130_fd_sc_hd__diode_2 ANTENNA__12136__C (.DIODE(net553));
 sky130_fd_sc_hd__diode_2 ANTENNA__12136__D (.DIODE(net557));
 sky130_fd_sc_hd__diode_2 ANTENNA__12137__A (.DIODE(net440));
 sky130_fd_sc_hd__diode_2 ANTENNA__12137__B (.DIODE(net561));
 sky130_fd_sc_hd__diode_2 ANTENNA__12138__A2 (.DIODE(net553));
 sky130_fd_sc_hd__diode_2 ANTENNA__12138__B1 (.DIODE(net557));
 sky130_fd_sc_hd__diode_2 ANTENNA__12142__A1 (.DIODE(net436));
 sky130_fd_sc_hd__diode_2 ANTENNA__12142__A2 (.DIODE(net561));
 sky130_fd_sc_hd__diode_2 ANTENNA__12142__B1 (.DIODE(net566));
 sky130_fd_sc_hd__diode_2 ANTENNA__12142__B2 (.DIODE(net431));
 sky130_fd_sc_hd__diode_2 ANTENNA__12143__A (.DIODE(net436));
 sky130_fd_sc_hd__diode_2 ANTENNA__12143__B (.DIODE(net431));
 sky130_fd_sc_hd__diode_2 ANTENNA__12143__C (.DIODE(net561));
 sky130_fd_sc_hd__diode_2 ANTENNA__12143__D (.DIODE(net566));
 sky130_fd_sc_hd__diode_2 ANTENNA__12145__A (.DIODE(net426));
 sky130_fd_sc_hd__diode_2 ANTENNA__12145__B (.DIODE(net571));
 sky130_fd_sc_hd__diode_2 ANTENNA__12151__A1 (.DIODE(net426));
 sky130_fd_sc_hd__diode_2 ANTENNA__12151__A2 (.DIODE(net571));
 sky130_fd_sc_hd__diode_2 ANTENNA__12152__A1_N (.DIODE(net413));
 sky130_fd_sc_hd__diode_2 ANTENNA__12152__A2_N (.DIODE(net582));
 sky130_fd_sc_hd__diode_2 ANTENNA__12155__A (.DIODE(net421));
 sky130_fd_sc_hd__diode_2 ANTENNA__12155__B (.DIODE(net417));
 sky130_fd_sc_hd__diode_2 ANTENNA__12155__C (.DIODE(net576));
 sky130_fd_sc_hd__diode_2 ANTENNA__12155__D (.DIODE(net582));
 sky130_fd_sc_hd__diode_2 ANTENNA__12162__A (.DIODE(net412));
 sky130_fd_sc_hd__diode_2 ANTENNA__12162__B (.DIODE(net582));
 sky130_fd_sc_hd__diode_2 ANTENNA__12180__C (.DIODE(net557));
 sky130_fd_sc_hd__diode_2 ANTENNA__12180__D (.DIODE(net561));
 sky130_fd_sc_hd__diode_2 ANTENNA__12181__A (.DIODE(net440));
 sky130_fd_sc_hd__diode_2 ANTENNA__12181__B (.DIODE(net566));
 sky130_fd_sc_hd__diode_2 ANTENNA__12182__A2 (.DIODE(net557));
 sky130_fd_sc_hd__diode_2 ANTENNA__12182__B1 (.DIODE(net561));
 sky130_fd_sc_hd__diode_2 ANTENNA__12186__A (.DIODE(net436));
 sky130_fd_sc_hd__diode_2 ANTENNA__12186__B (.DIODE(net431));
 sky130_fd_sc_hd__diode_2 ANTENNA__12186__C (.DIODE(net566));
 sky130_fd_sc_hd__diode_2 ANTENNA__12186__D (.DIODE(net571));
 sky130_fd_sc_hd__diode_2 ANTENNA__12187__A1 (.DIODE(net436));
 sky130_fd_sc_hd__diode_2 ANTENNA__12187__A2 (.DIODE(net566));
 sky130_fd_sc_hd__diode_2 ANTENNA__12187__B1 (.DIODE(net571));
 sky130_fd_sc_hd__diode_2 ANTENNA__12187__B2 (.DIODE(net431));
 sky130_fd_sc_hd__diode_2 ANTENNA__12189__A (.DIODE(net426));
 sky130_fd_sc_hd__diode_2 ANTENNA__12189__B (.DIODE(net576));
 sky130_fd_sc_hd__diode_2 ANTENNA__12190__A (.DIODE(net426));
 sky130_fd_sc_hd__diode_2 ANTENNA__12190__B (.DIODE(net576));
 sky130_fd_sc_hd__diode_2 ANTENNA__12196__A1 (.DIODE(net421));
 sky130_fd_sc_hd__diode_2 ANTENNA__12196__A2 (.DIODE(net576));
 sky130_fd_sc_hd__diode_2 ANTENNA__12196__B1 (.DIODE(net582));
 sky130_fd_sc_hd__diode_2 ANTENNA__12196__B2 (.DIODE(net417));
 sky130_fd_sc_hd__diode_2 ANTENNA__12214__C (.DIODE(net561));
 sky130_fd_sc_hd__diode_2 ANTENNA__12214__D (.DIODE(net566));
 sky130_fd_sc_hd__diode_2 ANTENNA__12215__A (.DIODE(net440));
 sky130_fd_sc_hd__diode_2 ANTENNA__12215__B (.DIODE(net571));
 sky130_fd_sc_hd__diode_2 ANTENNA__12216__A2 (.DIODE(net561));
 sky130_fd_sc_hd__diode_2 ANTENNA__12216__B1 (.DIODE(net566));
 sky130_fd_sc_hd__diode_2 ANTENNA__12220__A1 (.DIODE(net436));
 sky130_fd_sc_hd__diode_2 ANTENNA__12220__A2 (.DIODE(net571));
 sky130_fd_sc_hd__diode_2 ANTENNA__12220__B1 (.DIODE(net576));
 sky130_fd_sc_hd__diode_2 ANTENNA__12220__B2 (.DIODE(net431));
 sky130_fd_sc_hd__diode_2 ANTENNA__12221__A (.DIODE(net436));
 sky130_fd_sc_hd__diode_2 ANTENNA__12221__B (.DIODE(net431));
 sky130_fd_sc_hd__diode_2 ANTENNA__12221__C (.DIODE(net571));
 sky130_fd_sc_hd__diode_2 ANTENNA__12221__D (.DIODE(net576));
 sky130_fd_sc_hd__diode_2 ANTENNA__12223__A (.DIODE(net426));
 sky130_fd_sc_hd__diode_2 ANTENNA__12223__B (.DIODE(net582));
 sky130_fd_sc_hd__diode_2 ANTENNA__12229__A (.DIODE(net421));
 sky130_fd_sc_hd__diode_2 ANTENNA__12229__B (.DIODE(net582));
 sky130_fd_sc_hd__diode_2 ANTENNA__12242__A (.DIODE(net436));
 sky130_fd_sc_hd__diode_2 ANTENNA__12242__B (.DIODE(net431));
 sky130_fd_sc_hd__diode_2 ANTENNA__12242__C (.DIODE(net576));
 sky130_fd_sc_hd__diode_2 ANTENNA__12242__D (.DIODE(net582));
 sky130_fd_sc_hd__diode_2 ANTENNA__12245__C (.DIODE(net566));
 sky130_fd_sc_hd__diode_2 ANTENNA__12245__D (.DIODE(net571));
 sky130_fd_sc_hd__diode_2 ANTENNA__12246__C (.DIODE(net566));
 sky130_fd_sc_hd__diode_2 ANTENNA__12246__D (.DIODE(net571));
 sky130_fd_sc_hd__diode_2 ANTENNA__12247__A2 (.DIODE(net566));
 sky130_fd_sc_hd__diode_2 ANTENNA__12247__B1 (.DIODE(net571));
 sky130_fd_sc_hd__diode_2 ANTENNA__12248__A (.DIODE(net441));
 sky130_fd_sc_hd__diode_2 ANTENNA__12248__B (.DIODE(\mul0.a[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__12249__A (.DIODE(net440));
 sky130_fd_sc_hd__diode_2 ANTENNA__12249__B (.DIODE(\mul0.a[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__12251__A1 (.DIODE(net436));
 sky130_fd_sc_hd__diode_2 ANTENNA__12251__A2 (.DIODE(net576));
 sky130_fd_sc_hd__diode_2 ANTENNA__12251__B1 (.DIODE(net582));
 sky130_fd_sc_hd__diode_2 ANTENNA__12251__B2 (.DIODE(net431));
 sky130_fd_sc_hd__diode_2 ANTENNA__12260__A1 (.DIODE(net440));
 sky130_fd_sc_hd__diode_2 ANTENNA__12260__A2 (.DIODE(net576));
 sky130_fd_sc_hd__diode_2 ANTENNA__12261__C (.DIODE(net575));
 sky130_fd_sc_hd__diode_2 ANTENNA__12261__D (.DIODE(net576));
 sky130_fd_sc_hd__diode_2 ANTENNA__12262__A2 (.DIODE(net575));
 sky130_fd_sc_hd__diode_2 ANTENNA__12262__B1 (.DIODE(\mul0.a[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__12263__A1 (.DIODE(net440));
 sky130_fd_sc_hd__diode_2 ANTENNA__12263__A2 (.DIODE(net582));
 sky130_fd_sc_hd__diode_2 ANTENNA__12266__A1 (.DIODE(net436));
 sky130_fd_sc_hd__diode_2 ANTENNA__12266__A2 (.DIODE(net582));
 sky130_fd_sc_hd__diode_2 ANTENNA__12267__A (.DIODE(net436));
 sky130_fd_sc_hd__diode_2 ANTENNA__12267__B (.DIODE(net582));
 sky130_fd_sc_hd__diode_2 ANTENNA__12268__A (.DIODE(net440));
 sky130_fd_sc_hd__diode_2 ANTENNA__12268__B (.DIODE(net575));
 sky130_fd_sc_hd__diode_2 ANTENNA__12269__C (.DIODE(net576));
 sky130_fd_sc_hd__diode_2 ANTENNA__12269__D (.DIODE(net582));
 sky130_fd_sc_hd__diode_2 ANTENNA__12290__A (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__12290__B (.DIODE(_03792_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12291__A (.DIODE(net600));
 sky130_fd_sc_hd__diode_2 ANTENNA__12291__B (.DIODE(_03058_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12292__A1 (.DIODE(net599));
 sky130_fd_sc_hd__diode_2 ANTENNA__12292__B1 (.DIODE(_02738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12292__B2 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__12298__A1 (.DIODE(net371));
 sky130_fd_sc_hd__diode_2 ANTENNA__12298__A2 (.DIODE(net581));
 sky130_fd_sc_hd__diode_2 ANTENNA__12299__A1 (.DIODE(net386));
 sky130_fd_sc_hd__diode_2 ANTENNA__12299__A2 (.DIODE(net567));
 sky130_fd_sc_hd__diode_2 ANTENNA__12300__A (.DIODE(net567));
 sky130_fd_sc_hd__diode_2 ANTENNA__12300__B (.DIODE(net572));
 sky130_fd_sc_hd__diode_2 ANTENNA__12300__C (.DIODE(net381));
 sky130_fd_sc_hd__diode_2 ANTENNA__12300__D (.DIODE(net375));
 sky130_fd_sc_hd__diode_2 ANTENNA__12301__A1 (.DIODE(net567));
 sky130_fd_sc_hd__diode_2 ANTENNA__12301__A2 (.DIODE(net381));
 sky130_fd_sc_hd__diode_2 ANTENNA__12301__B1 (.DIODE(net375));
 sky130_fd_sc_hd__diode_2 ANTENNA__12301__B2 (.DIODE(net572));
 sky130_fd_sc_hd__diode_2 ANTENNA__12302__A (.DIODE(net577));
 sky130_fd_sc_hd__diode_2 ANTENNA__12302__B (.DIODE(net371));
 sky130_fd_sc_hd__diode_2 ANTENNA__12303__A1 (.DIODE(net580));
 sky130_fd_sc_hd__diode_2 ANTENNA__12303__A2 (.DIODE(net371));
 sky130_fd_sc_hd__diode_2 ANTENNA__12311__A (.DIODE(net581));
 sky130_fd_sc_hd__diode_2 ANTENNA__12311__B (.DIODE(net631));
 sky130_fd_sc_hd__diode_2 ANTENNA__12312__A (.DIODE(net581));
 sky130_fd_sc_hd__diode_2 ANTENNA__12312__B (.DIODE(net631));
 sky130_fd_sc_hd__diode_2 ANTENNA__12319__A (.DIODE(net554));
 sky130_fd_sc_hd__diode_2 ANTENNA__12319__B (.DIODE(net560));
 sky130_fd_sc_hd__diode_2 ANTENNA__12319__C (.DIODE(net396));
 sky130_fd_sc_hd__diode_2 ANTENNA__12319__D (.DIODE(net390));
 sky130_fd_sc_hd__diode_2 ANTENNA__12321__A1 (.DIODE(net553));
 sky130_fd_sc_hd__diode_2 ANTENNA__12321__A2 (.DIODE(net396));
 sky130_fd_sc_hd__diode_2 ANTENNA__12321__B1 (.DIODE(net390));
 sky130_fd_sc_hd__diode_2 ANTENNA__12321__B2 (.DIODE(net560));
 sky130_fd_sc_hd__diode_2 ANTENNA__12322__C (.DIODE(net564));
 sky130_fd_sc_hd__diode_2 ANTENNA__12322__D (.DIODE(net389));
 sky130_fd_sc_hd__diode_2 ANTENNA__12323__A1 (.DIODE(net564));
 sky130_fd_sc_hd__diode_2 ANTENNA__12323__A2 (.DIODE(net386));
 sky130_fd_sc_hd__diode_2 ANTENNA__12325__A (.DIODE(net549));
 sky130_fd_sc_hd__diode_2 ANTENNA__12325__B (.DIODE(net401));
 sky130_fd_sc_hd__diode_2 ANTENNA__12326__A (.DIODE(net541));
 sky130_fd_sc_hd__diode_2 ANTENNA__12326__B (.DIODE(net545));
 sky130_fd_sc_hd__diode_2 ANTENNA__12326__C (.DIODE(net409));
 sky130_fd_sc_hd__diode_2 ANTENNA__12326__D (.DIODE(net404));
 sky130_fd_sc_hd__diode_2 ANTENNA__12327__A1 (.DIODE(net541));
 sky130_fd_sc_hd__diode_2 ANTENNA__12327__A2 (.DIODE(net409));
 sky130_fd_sc_hd__diode_2 ANTENNA__12327__B1 (.DIODE(net404));
 sky130_fd_sc_hd__diode_2 ANTENNA__12327__B2 (.DIODE(net545));
 sky130_fd_sc_hd__diode_2 ANTENNA__12340__A1 (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA__12340__A2 (.DIODE(net541));
 sky130_fd_sc_hd__diode_2 ANTENNA__12342__A (.DIODE(net536));
 sky130_fd_sc_hd__diode_2 ANTENNA__12342__B (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA__12343__A (.DIODE(net525));
 sky130_fd_sc_hd__diode_2 ANTENNA__12343__C (.DIODE(net422));
 sky130_fd_sc_hd__diode_2 ANTENNA__12343__D (.DIODE(net418));
 sky130_fd_sc_hd__diode_2 ANTENNA__12344__A1 (.DIODE(net525));
 sky130_fd_sc_hd__diode_2 ANTENNA__12344__A2 (.DIODE(net422));
 sky130_fd_sc_hd__diode_2 ANTENNA__12344__B1 (.DIODE(net418));
 sky130_fd_sc_hd__diode_2 ANTENNA__12351__A (.DIODE(net520));
 sky130_fd_sc_hd__diode_2 ANTENNA__12351__B (.DIODE(net427));
 sky130_fd_sc_hd__diode_2 ANTENNA__12352__A1 (.DIODE(net511));
 sky130_fd_sc_hd__diode_2 ANTENNA__12352__A2 (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA__12352__B1 (.DIODE(net432));
 sky130_fd_sc_hd__diode_2 ANTENNA__12352__B2 (.DIODE(net515));
 sky130_fd_sc_hd__diode_2 ANTENNA__12353__A (.DIODE(net511));
 sky130_fd_sc_hd__diode_2 ANTENNA__12353__B (.DIODE(net515));
 sky130_fd_sc_hd__diode_2 ANTENNA__12353__C (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA__12353__D (.DIODE(net432));
 sky130_fd_sc_hd__diode_2 ANTENNA__12356__A (.DIODE(net507));
 sky130_fd_sc_hd__diode_2 ANTENNA__12356__B (.DIODE(net441));
 sky130_fd_sc_hd__diode_2 ANTENNA__12357__B (.DIODE(net503));
 sky130_fd_sc_hd__diode_2 ANTENNA__12357__D (.DIODE(net498));
 sky130_fd_sc_hd__diode_2 ANTENNA__12358__A1 (.DIODE(net503));
 sky130_fd_sc_hd__diode_2 ANTENNA__12358__B1 (.DIODE(net498));
 sky130_fd_sc_hd__diode_2 ANTENNA__12392__A (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__12392__B (.DIODE(_03893_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12393__A1 (.DIODE(net599));
 sky130_fd_sc_hd__diode_2 ANTENNA__12393__B1 (.DIODE(_02739_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12393__B2 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__12396__A1 (.DIODE(net580));
 sky130_fd_sc_hd__diode_2 ANTENNA__12396__A2 (.DIODE(net631));
 sky130_fd_sc_hd__diode_2 ANTENNA__12396__B1 (.DIODE(net365));
 sky130_fd_sc_hd__diode_2 ANTENNA__12396__B2 (.DIODE(net581));
 sky130_fd_sc_hd__diode_2 ANTENNA__12397__A (.DIODE(net578));
 sky130_fd_sc_hd__diode_2 ANTENNA__12397__B (.DIODE(net583));
 sky130_fd_sc_hd__diode_2 ANTENNA__12397__C (.DIODE(net631));
 sky130_fd_sc_hd__diode_2 ANTENNA__12397__D (.DIODE(net365));
 sky130_fd_sc_hd__diode_2 ANTENNA__12400__A1 (.DIODE(net567));
 sky130_fd_sc_hd__diode_2 ANTENNA__12400__A2 (.DIODE(net572));
 sky130_fd_sc_hd__diode_2 ANTENNA__12400__A3 (.DIODE(net381));
 sky130_fd_sc_hd__diode_2 ANTENNA__12400__A4 (.DIODE(net375));
 sky130_fd_sc_hd__diode_2 ANTENNA__12402__A (.DIODE(net572));
 sky130_fd_sc_hd__diode_2 ANTENNA__12402__B (.DIODE(net371));
 sky130_fd_sc_hd__diode_2 ANTENNA__12403__A (.DIODE(net564));
 sky130_fd_sc_hd__diode_2 ANTENNA__12403__B (.DIODE(net570));
 sky130_fd_sc_hd__diode_2 ANTENNA__12403__C (.DIODE(net381));
 sky130_fd_sc_hd__diode_2 ANTENNA__12403__D (.DIODE(net375));
 sky130_fd_sc_hd__diode_2 ANTENNA__12404__A1 (.DIODE(net564));
 sky130_fd_sc_hd__diode_2 ANTENNA__12404__A2 (.DIODE(net381));
 sky130_fd_sc_hd__diode_2 ANTENNA__12404__B1 (.DIODE(net375));
 sky130_fd_sc_hd__diode_2 ANTENNA__12404__B2 (.DIODE(net570));
 sky130_fd_sc_hd__diode_2 ANTENNA__12420__A (.DIODE(net549));
 sky130_fd_sc_hd__diode_2 ANTENNA__12420__B (.DIODE(net553));
 sky130_fd_sc_hd__diode_2 ANTENNA__12420__C (.DIODE(net395));
 sky130_fd_sc_hd__diode_2 ANTENNA__12420__D (.DIODE(net390));
 sky130_fd_sc_hd__diode_2 ANTENNA__12422__A1 (.DIODE(net549));
 sky130_fd_sc_hd__diode_2 ANTENNA__12422__A2 (.DIODE(net396));
 sky130_fd_sc_hd__diode_2 ANTENNA__12422__B1 (.DIODE(net390));
 sky130_fd_sc_hd__diode_2 ANTENNA__12422__B2 (.DIODE(net553));
 sky130_fd_sc_hd__diode_2 ANTENNA__12423__C (.DIODE(net557));
 sky130_fd_sc_hd__diode_2 ANTENNA__12423__D (.DIODE(net389));
 sky130_fd_sc_hd__diode_2 ANTENNA__12424__A1 (.DIODE(net557));
 sky130_fd_sc_hd__diode_2 ANTENNA__12424__A2 (.DIODE(net389));
 sky130_fd_sc_hd__diode_2 ANTENNA__12426__A (.DIODE(net545));
 sky130_fd_sc_hd__diode_2 ANTENNA__12426__B (.DIODE(net400));
 sky130_fd_sc_hd__diode_2 ANTENNA__12427__A (.DIODE(net536));
 sky130_fd_sc_hd__diode_2 ANTENNA__12427__B (.DIODE(net541));
 sky130_fd_sc_hd__diode_2 ANTENNA__12427__C (.DIODE(net409));
 sky130_fd_sc_hd__diode_2 ANTENNA__12427__D (.DIODE(net405));
 sky130_fd_sc_hd__diode_2 ANTENNA__12428__A1 (.DIODE(net536));
 sky130_fd_sc_hd__diode_2 ANTENNA__12428__A2 (.DIODE(net412));
 sky130_fd_sc_hd__diode_2 ANTENNA__12428__B1 (.DIODE(net405));
 sky130_fd_sc_hd__diode_2 ANTENNA__12428__B2 (.DIODE(net541));
 sky130_fd_sc_hd__diode_2 ANTENNA__12431__A1 (.DIODE(net548));
 sky130_fd_sc_hd__diode_2 ANTENNA__12431__A2 (.DIODE(net400));
 sky130_fd_sc_hd__diode_2 ANTENNA__12441__A1 (.DIODE(net535));
 sky130_fd_sc_hd__diode_2 ANTENNA__12441__A2 (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA__12443__B (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA__12444__A (.DIODE(net520));
 sky130_fd_sc_hd__diode_2 ANTENNA__12444__B (.DIODE(net525));
 sky130_fd_sc_hd__diode_2 ANTENNA__12444__C (.DIODE(net425));
 sky130_fd_sc_hd__diode_2 ANTENNA__12444__D (.DIODE(net418));
 sky130_fd_sc_hd__diode_2 ANTENNA__12445__A1 (.DIODE(net520));
 sky130_fd_sc_hd__diode_2 ANTENNA__12445__A2 (.DIODE(net425));
 sky130_fd_sc_hd__diode_2 ANTENNA__12445__B1 (.DIODE(net418));
 sky130_fd_sc_hd__diode_2 ANTENNA__12445__B2 (.DIODE(net525));
 sky130_fd_sc_hd__diode_2 ANTENNA__12452__A (.DIODE(net515));
 sky130_fd_sc_hd__diode_2 ANTENNA__12452__B (.DIODE(net427));
 sky130_fd_sc_hd__diode_2 ANTENNA__12453__A1 (.DIODE(net507));
 sky130_fd_sc_hd__diode_2 ANTENNA__12453__A2 (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA__12453__B1 (.DIODE(net432));
 sky130_fd_sc_hd__diode_2 ANTENNA__12453__B2 (.DIODE(net511));
 sky130_fd_sc_hd__diode_2 ANTENNA__12454__A (.DIODE(net507));
 sky130_fd_sc_hd__diode_2 ANTENNA__12454__B (.DIODE(net511));
 sky130_fd_sc_hd__diode_2 ANTENNA__12454__C (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA__12454__D (.DIODE(net432));
 sky130_fd_sc_hd__diode_2 ANTENNA__12457__A (.DIODE(net503));
 sky130_fd_sc_hd__diode_2 ANTENNA__12457__B (.DIODE(net441));
 sky130_fd_sc_hd__diode_2 ANTENNA__12458__B (.DIODE(net446));
 sky130_fd_sc_hd__diode_2 ANTENNA__12458__C (.DIODE(net498));
 sky130_fd_sc_hd__diode_2 ANTENNA__12458__D (.DIODE(net494));
 sky130_fd_sc_hd__diode_2 ANTENNA__12459__A2 (.DIODE(net498));
 sky130_fd_sc_hd__diode_2 ANTENNA__12459__B1 (.DIODE(net494));
 sky130_fd_sc_hd__diode_2 ANTENNA__12493__A (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__12493__B (.DIODE(_03993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12494__A1 (.DIODE(net599));
 sky130_fd_sc_hd__diode_2 ANTENNA__12494__B1 (.DIODE(_02741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12494__B2 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__12501__A (.DIODE(net574));
 sky130_fd_sc_hd__diode_2 ANTENNA__12501__B (.DIODE(net578));
 sky130_fd_sc_hd__diode_2 ANTENNA__12501__C (.DIODE(net631));
 sky130_fd_sc_hd__diode_2 ANTENNA__12501__D (.DIODE(net365));
 sky130_fd_sc_hd__diode_2 ANTENNA__12502__A1 (.DIODE(net574));
 sky130_fd_sc_hd__diode_2 ANTENNA__12502__A2 (.DIODE(net631));
 sky130_fd_sc_hd__diode_2 ANTENNA__12502__B1 (.DIODE(net365));
 sky130_fd_sc_hd__diode_2 ANTENNA__12502__B2 (.DIODE(net578));
 sky130_fd_sc_hd__diode_2 ANTENNA__12504__A (.DIODE(net583));
 sky130_fd_sc_hd__diode_2 ANTENNA__12504__B (.DIODE(net364));
 sky130_fd_sc_hd__diode_2 ANTENNA__12509__A1 (.DIODE(net572));
 sky130_fd_sc_hd__diode_2 ANTENNA__12509__A2 (.DIODE(net371));
 sky130_fd_sc_hd__diode_2 ANTENNA__12511__A (.DIODE(net567));
 sky130_fd_sc_hd__diode_2 ANTENNA__12511__B (.DIODE(net370));
 sky130_fd_sc_hd__diode_2 ANTENNA__12512__A (.DIODE(net557));
 sky130_fd_sc_hd__diode_2 ANTENNA__12512__B (.DIODE(net565));
 sky130_fd_sc_hd__diode_2 ANTENNA__12512__C (.DIODE(net381));
 sky130_fd_sc_hd__diode_2 ANTENNA__12512__D (.DIODE(net375));
 sky130_fd_sc_hd__diode_2 ANTENNA__12513__A1 (.DIODE(net557));
 sky130_fd_sc_hd__diode_2 ANTENNA__12513__A2 (.DIODE(net381));
 sky130_fd_sc_hd__diode_2 ANTENNA__12513__B1 (.DIODE(net375));
 sky130_fd_sc_hd__diode_2 ANTENNA__12513__B2 (.DIODE(net561));
 sky130_fd_sc_hd__diode_2 ANTENNA__12528__A (.DIODE(net545));
 sky130_fd_sc_hd__diode_2 ANTENNA__12528__B (.DIODE(net548));
 sky130_fd_sc_hd__diode_2 ANTENNA__12528__C (.DIODE(net395));
 sky130_fd_sc_hd__diode_2 ANTENNA__12529__A1 (.DIODE(net545));
 sky130_fd_sc_hd__diode_2 ANTENNA__12529__A2 (.DIODE(net395));
 sky130_fd_sc_hd__diode_2 ANTENNA__12529__B2 (.DIODE(net548));
 sky130_fd_sc_hd__diode_2 ANTENNA__12530__A (.DIODE(net553));
 sky130_fd_sc_hd__diode_2 ANTENNA__12530__B (.DIODE(net386));
 sky130_fd_sc_hd__diode_2 ANTENNA__12531__A1 (.DIODE(net553));
 sky130_fd_sc_hd__diode_2 ANTENNA__12531__A2 (.DIODE(net386));
 sky130_fd_sc_hd__diode_2 ANTENNA__12533__A (.DIODE(net541));
 sky130_fd_sc_hd__diode_2 ANTENNA__12533__B (.DIODE(net401));
 sky130_fd_sc_hd__diode_2 ANTENNA__12534__B (.DIODE(net536));
 sky130_fd_sc_hd__diode_2 ANTENNA__12534__C (.DIODE(net409));
 sky130_fd_sc_hd__diode_2 ANTENNA__12534__D (.DIODE(net405));
 sky130_fd_sc_hd__diode_2 ANTENNA__12535__A2 (.DIODE(net409));
 sky130_fd_sc_hd__diode_2 ANTENNA__12535__B1 (.DIODE(net405));
 sky130_fd_sc_hd__diode_2 ANTENNA__12535__B2 (.DIODE(net536));
 sky130_fd_sc_hd__diode_2 ANTENNA__12538__A1 (.DIODE(net545));
 sky130_fd_sc_hd__diode_2 ANTENNA__12538__A2 (.DIODE(net401));
 sky130_fd_sc_hd__diode_2 ANTENNA__12548__A2 (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA__12550__B (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA__12551__A (.DIODE(net515));
 sky130_fd_sc_hd__diode_2 ANTENNA__12551__B (.DIODE(net520));
 sky130_fd_sc_hd__diode_2 ANTENNA__12551__C (.DIODE(net422));
 sky130_fd_sc_hd__diode_2 ANTENNA__12551__D (.DIODE(net418));
 sky130_fd_sc_hd__diode_2 ANTENNA__12552__A1 (.DIODE(net515));
 sky130_fd_sc_hd__diode_2 ANTENNA__12552__A2 (.DIODE(net422));
 sky130_fd_sc_hd__diode_2 ANTENNA__12552__B1 (.DIODE(net418));
 sky130_fd_sc_hd__diode_2 ANTENNA__12552__B2 (.DIODE(net520));
 sky130_fd_sc_hd__diode_2 ANTENNA__12559__A (.DIODE(net511));
 sky130_fd_sc_hd__diode_2 ANTENNA__12559__B (.DIODE(net427));
 sky130_fd_sc_hd__diode_2 ANTENNA__12560__A (.DIODE(net503));
 sky130_fd_sc_hd__diode_2 ANTENNA__12560__B (.DIODE(net507));
 sky130_fd_sc_hd__diode_2 ANTENNA__12560__C (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA__12560__D (.DIODE(net432));
 sky130_fd_sc_hd__diode_2 ANTENNA__12561__A1 (.DIODE(net503));
 sky130_fd_sc_hd__diode_2 ANTENNA__12561__A2 (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA__12561__B1 (.DIODE(net432));
 sky130_fd_sc_hd__diode_2 ANTENNA__12561__B2 (.DIODE(net507));
 sky130_fd_sc_hd__diode_2 ANTENNA__12564__A (.DIODE(net441));
 sky130_fd_sc_hd__diode_2 ANTENNA__12564__B (.DIODE(net498));
 sky130_fd_sc_hd__diode_2 ANTENNA__12565__A (.DIODE(net452));
 sky130_fd_sc_hd__diode_2 ANTENNA__12565__B (.DIODE(net446));
 sky130_fd_sc_hd__diode_2 ANTENNA__12565__C (.DIODE(net494));
 sky130_fd_sc_hd__diode_2 ANTENNA__12565__D (.DIODE(net490));
 sky130_fd_sc_hd__diode_2 ANTENNA__12566__A1 (.DIODE(net446));
 sky130_fd_sc_hd__diode_2 ANTENNA__12566__A2 (.DIODE(net494));
 sky130_fd_sc_hd__diode_2 ANTENNA__12566__B1 (.DIODE(net490));
 sky130_fd_sc_hd__diode_2 ANTENNA__12566__B2 (.DIODE(net452));
 sky130_fd_sc_hd__diode_2 ANTENNA__12601__A (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__12601__B (.DIODE(_04100_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12602__A1 (.DIODE(net599));
 sky130_fd_sc_hd__diode_2 ANTENNA__12602__B1 (.DIODE(_02743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12602__B2 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__12607__A (.DIODE(net568));
 sky130_fd_sc_hd__diode_2 ANTENNA__12607__C (.DIODE(\mul0.b[18] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__12607__D (.DIODE(net365));
 sky130_fd_sc_hd__diode_2 ANTENNA__12609__A1 (.DIODE(net568));
 sky130_fd_sc_hd__diode_2 ANTENNA__12609__A2 (.DIODE(net631));
 sky130_fd_sc_hd__diode_2 ANTENNA__12609__B1 (.DIODE(net365));
 sky130_fd_sc_hd__diode_2 ANTENNA__12610__A (.DIODE(net578));
 sky130_fd_sc_hd__diode_2 ANTENNA__12610__B (.DIODE(net364));
 sky130_fd_sc_hd__diode_2 ANTENNA__12611__A1 (.DIODE(net578));
 sky130_fd_sc_hd__diode_2 ANTENNA__12611__A2 (.DIODE(net364));
 sky130_fd_sc_hd__diode_2 ANTENNA__12616__A (.DIODE(net583));
 sky130_fd_sc_hd__diode_2 ANTENNA__12616__B (.DIODE(net360));
 sky130_fd_sc_hd__diode_2 ANTENNA__12618__A1 (.DIODE(net568));
 sky130_fd_sc_hd__diode_2 ANTENNA__12618__A2 (.DIODE(net370));
 sky130_fd_sc_hd__diode_2 ANTENNA__12619__A (.DIODE(net552));
 sky130_fd_sc_hd__diode_2 ANTENNA__12619__B (.DIODE(net558));
 sky130_fd_sc_hd__diode_2 ANTENNA__12619__C (.DIODE(net382));
 sky130_fd_sc_hd__diode_2 ANTENNA__12619__D (.DIODE(net375));
 sky130_fd_sc_hd__diode_2 ANTENNA__12620__A1 (.DIODE(net552));
 sky130_fd_sc_hd__diode_2 ANTENNA__12620__A2 (.DIODE(net382));
 sky130_fd_sc_hd__diode_2 ANTENNA__12620__B1 (.DIODE(net375));
 sky130_fd_sc_hd__diode_2 ANTENNA__12620__B2 (.DIODE(net558));
 sky130_fd_sc_hd__diode_2 ANTENNA__12621__C (.DIODE(net565));
 sky130_fd_sc_hd__diode_2 ANTENNA__12621__D (.DIODE(net370));
 sky130_fd_sc_hd__diode_2 ANTENNA__12622__A1_N (.DIODE(net565));
 sky130_fd_sc_hd__diode_2 ANTENNA__12622__A2_N (.DIODE(net370));
 sky130_fd_sc_hd__diode_2 ANTENNA__12637__A (.DIODE(net541));
 sky130_fd_sc_hd__diode_2 ANTENNA__12637__B (.DIODE(net544));
 sky130_fd_sc_hd__diode_2 ANTENNA__12637__C (.DIODE(net395));
 sky130_fd_sc_hd__diode_2 ANTENNA__12638__A1 (.DIODE(net541));
 sky130_fd_sc_hd__diode_2 ANTENNA__12638__A2 (.DIODE(net395));
 sky130_fd_sc_hd__diode_2 ANTENNA__12638__B2 (.DIODE(net545));
 sky130_fd_sc_hd__diode_2 ANTENNA__12639__A (.DIODE(net549));
 sky130_fd_sc_hd__diode_2 ANTENNA__12639__B (.DIODE(net386));
 sky130_fd_sc_hd__diode_2 ANTENNA__12640__A1 (.DIODE(net548));
 sky130_fd_sc_hd__diode_2 ANTENNA__12640__A2 (.DIODE(net389));
 sky130_fd_sc_hd__diode_2 ANTENNA__12642__A (.DIODE(net536));
 sky130_fd_sc_hd__diode_2 ANTENNA__12642__B (.DIODE(net401));
 sky130_fd_sc_hd__diode_2 ANTENNA__12643__C (.DIODE(net409));
 sky130_fd_sc_hd__diode_2 ANTENNA__12643__D (.DIODE(net405));
 sky130_fd_sc_hd__diode_2 ANTENNA__12644__A2 (.DIODE(net409));
 sky130_fd_sc_hd__diode_2 ANTENNA__12644__B1 (.DIODE(net405));
 sky130_fd_sc_hd__diode_2 ANTENNA__12647__A1 (.DIODE(net541));
 sky130_fd_sc_hd__diode_2 ANTENNA__12647__A2 (.DIODE(net401));
 sky130_fd_sc_hd__diode_2 ANTENNA__12657__A2 (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA__12659__A (.DIODE(net521));
 sky130_fd_sc_hd__diode_2 ANTENNA__12659__B (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA__12660__A (.DIODE(net512));
 sky130_fd_sc_hd__diode_2 ANTENNA__12660__B (.DIODE(net516));
 sky130_fd_sc_hd__diode_2 ANTENNA__12660__C (.DIODE(\mul0.b[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__12661__A1 (.DIODE(net511));
 sky130_fd_sc_hd__diode_2 ANTENNA__12661__A2 (.DIODE(net425));
 sky130_fd_sc_hd__diode_2 ANTENNA__12661__B1 (.DIODE(\mul0.b[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__12661__B2 (.DIODE(net516));
 sky130_fd_sc_hd__diode_2 ANTENNA__12662__A1 (.DIODE(net422));
 sky130_fd_sc_hd__diode_2 ANTENNA__12668__A1 (.DIODE(net503));
 sky130_fd_sc_hd__diode_2 ANTENNA__12668__A2 (.DIODE(net432));
 sky130_fd_sc_hd__diode_2 ANTENNA__12668__B1 (.DIODE(net498));
 sky130_fd_sc_hd__diode_2 ANTENNA__12668__B2 (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA__12669__A (.DIODE(net503));
 sky130_fd_sc_hd__diode_2 ANTENNA__12669__B (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA__12669__C (.DIODE(net432));
 sky130_fd_sc_hd__diode_2 ANTENNA__12669__D (.DIODE(net498));
 sky130_fd_sc_hd__diode_2 ANTENNA__12670__C (.DIODE(net507));
 sky130_fd_sc_hd__diode_2 ANTENNA__12670__D (.DIODE(net427));
 sky130_fd_sc_hd__diode_2 ANTENNA__12671__A1_N (.DIODE(net507));
 sky130_fd_sc_hd__diode_2 ANTENNA__12671__A2_N (.DIODE(net427));
 sky130_fd_sc_hd__diode_2 ANTENNA__12673__A (.DIODE(net441));
 sky130_fd_sc_hd__diode_2 ANTENNA__12673__B (.DIODE(net494));
 sky130_fd_sc_hd__diode_2 ANTENNA__12674__A (.DIODE(net452));
 sky130_fd_sc_hd__diode_2 ANTENNA__12674__B (.DIODE(net446));
 sky130_fd_sc_hd__diode_2 ANTENNA__12674__C (.DIODE(net490));
 sky130_fd_sc_hd__diode_2 ANTENNA__12674__D (.DIODE(net486));
 sky130_fd_sc_hd__diode_2 ANTENNA__12675__A1 (.DIODE(net446));
 sky130_fd_sc_hd__diode_2 ANTENNA__12675__A2 (.DIODE(net490));
 sky130_fd_sc_hd__diode_2 ANTENNA__12675__B1 (.DIODE(net486));
 sky130_fd_sc_hd__diode_2 ANTENNA__12675__B2 (.DIODE(net452));
 sky130_fd_sc_hd__diode_2 ANTENNA__12711__A (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__12711__B (.DIODE(_04209_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12712__A1 (.DIODE(net599));
 sky130_fd_sc_hd__diode_2 ANTENNA__12712__B1 (.DIODE(_02744_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12712__B2 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__12714__A1 (.DIODE(net583));
 sky130_fd_sc_hd__diode_2 ANTENNA__12714__A2 (.DIODE(net360));
 sky130_fd_sc_hd__diode_2 ANTENNA__12718__A1 (.DIODE(net578));
 sky130_fd_sc_hd__diode_2 ANTENNA__12718__A2 (.DIODE(net360));
 sky130_fd_sc_hd__diode_2 ANTENNA__12718__B1 (.DIODE(net355));
 sky130_fd_sc_hd__diode_2 ANTENNA__12718__B2 (.DIODE(net583));
 sky130_fd_sc_hd__diode_2 ANTENNA__12720__A (.DIODE(net578));
 sky130_fd_sc_hd__diode_2 ANTENNA__12720__B (.DIODE(net583));
 sky130_fd_sc_hd__diode_2 ANTENNA__12720__C (.DIODE(net360));
 sky130_fd_sc_hd__diode_2 ANTENNA__12720__D (.DIODE(net355));
 sky130_fd_sc_hd__diode_2 ANTENNA__12722__B (.DIODE(net568));
 sky130_fd_sc_hd__diode_2 ANTENNA__12722__C (.DIODE(net631));
 sky130_fd_sc_hd__diode_2 ANTENNA__12722__D (.DIODE(net365));
 sky130_fd_sc_hd__diode_2 ANTENNA__12724__A2 (.DIODE(net631));
 sky130_fd_sc_hd__diode_2 ANTENNA__12724__B1 (.DIODE(net365));
 sky130_fd_sc_hd__diode_2 ANTENNA__12724__B2 (.DIODE(net568));
 sky130_fd_sc_hd__diode_2 ANTENNA__12725__B (.DIODE(net364));
 sky130_fd_sc_hd__diode_2 ANTENNA__12726__A2 (.DIODE(net364));
 sky130_fd_sc_hd__diode_2 ANTENNA__12733__A (.DIODE(net550));
 sky130_fd_sc_hd__diode_2 ANTENNA__12733__B (.DIODE(net554));
 sky130_fd_sc_hd__diode_2 ANTENNA__12733__C (.DIODE(net381));
 sky130_fd_sc_hd__diode_2 ANTENNA__12734__A1 (.DIODE(net550));
 sky130_fd_sc_hd__diode_2 ANTENNA__12734__A2 (.DIODE(net382));
 sky130_fd_sc_hd__diode_2 ANTENNA__12734__B2 (.DIODE(net554));
 sky130_fd_sc_hd__diode_2 ANTENNA__12735__C (.DIODE(net558));
 sky130_fd_sc_hd__diode_2 ANTENNA__12735__D (.DIODE(net370));
 sky130_fd_sc_hd__diode_2 ANTENNA__12736__A1_N (.DIODE(net558));
 sky130_fd_sc_hd__diode_2 ANTENNA__12736__A2_N (.DIODE(net370));
 sky130_fd_sc_hd__diode_2 ANTENNA__12750__A (.DIODE(net545));
 sky130_fd_sc_hd__diode_2 ANTENNA__12750__B (.DIODE(net389));
 sky130_fd_sc_hd__diode_2 ANTENNA__12751__A (.DIODE(net535));
 sky130_fd_sc_hd__diode_2 ANTENNA__12751__B (.DIODE(net540));
 sky130_fd_sc_hd__diode_2 ANTENNA__12752__A1 (.DIODE(net535));
 sky130_fd_sc_hd__diode_2 ANTENNA__12752__A2 (.DIODE(net395));
 sky130_fd_sc_hd__diode_2 ANTENNA__12752__B2 (.DIODE(net541));
 sky130_fd_sc_hd__diode_2 ANTENNA__12753__A1 (.DIODE(net395));
 sky130_fd_sc_hd__diode_2 ANTENNA__12755__B (.DIODE(net401));
 sky130_fd_sc_hd__diode_2 ANTENNA__12756__A (.DIODE(net521));
 sky130_fd_sc_hd__diode_2 ANTENNA__12756__C (.DIODE(net405));
 sky130_fd_sc_hd__diode_2 ANTENNA__12757__A1 (.DIODE(net521));
 sky130_fd_sc_hd__diode_2 ANTENNA__12757__A2 (.DIODE(net409));
 sky130_fd_sc_hd__diode_2 ANTENNA__12757__B1 (.DIODE(net405));
 sky130_fd_sc_hd__diode_2 ANTENNA__12758__A1 (.DIODE(net409));
 sky130_fd_sc_hd__diode_2 ANTENNA__12760__A1 (.DIODE(net536));
 sky130_fd_sc_hd__diode_2 ANTENNA__12760__A2 (.DIODE(net401));
 sky130_fd_sc_hd__diode_2 ANTENNA__12770__A1 (.DIODE(net521));
 sky130_fd_sc_hd__diode_2 ANTENNA__12770__A2 (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA__12770__B2 (.DIODE(net425));
 sky130_fd_sc_hd__diode_2 ANTENNA__12771__A (.DIODE(net507));
 sky130_fd_sc_hd__diode_2 ANTENNA__12771__B (.DIODE(net512));
 sky130_fd_sc_hd__diode_2 ANTENNA__12771__C (.DIODE(net425));
 sky130_fd_sc_hd__diode_2 ANTENNA__12771__D (.DIODE(\mul0.b[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__12772__A1 (.DIODE(net507));
 sky130_fd_sc_hd__diode_2 ANTENNA__12772__A2 (.DIODE(net425));
 sky130_fd_sc_hd__diode_2 ANTENNA__12772__B1 (.DIODE(\mul0.b[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__12772__B2 (.DIODE(net512));
 sky130_fd_sc_hd__diode_2 ANTENNA__12773__A (.DIODE(net516));
 sky130_fd_sc_hd__diode_2 ANTENNA__12773__B (.DIODE(\mul0.b[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__12774__A1 (.DIODE(net516));
 sky130_fd_sc_hd__diode_2 ANTENNA__12774__A2 (.DIODE(\mul0.b[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__12779__A1 (.DIODE(net432));
 sky130_fd_sc_hd__diode_2 ANTENNA__12779__A2 (.DIODE(net498));
 sky130_fd_sc_hd__diode_2 ANTENNA__12779__B1 (.DIODE(net494));
 sky130_fd_sc_hd__diode_2 ANTENNA__12779__B2 (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA__12780__A (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA__12780__B (.DIODE(net432));
 sky130_fd_sc_hd__diode_2 ANTENNA__12780__C (.DIODE(net498));
 sky130_fd_sc_hd__diode_2 ANTENNA__12780__D (.DIODE(net494));
 sky130_fd_sc_hd__diode_2 ANTENNA__12781__C (.DIODE(net503));
 sky130_fd_sc_hd__diode_2 ANTENNA__12781__D (.DIODE(net427));
 sky130_fd_sc_hd__diode_2 ANTENNA__12782__A1_N (.DIODE(net503));
 sky130_fd_sc_hd__diode_2 ANTENNA__12782__A2_N (.DIODE(net427));
 sky130_fd_sc_hd__diode_2 ANTENNA__12784__A (.DIODE(net441));
 sky130_fd_sc_hd__diode_2 ANTENNA__12784__B (.DIODE(net490));
 sky130_fd_sc_hd__diode_2 ANTENNA__12785__A (.DIODE(net452));
 sky130_fd_sc_hd__diode_2 ANTENNA__12785__B (.DIODE(net446));
 sky130_fd_sc_hd__diode_2 ANTENNA__12785__C (.DIODE(net486));
 sky130_fd_sc_hd__diode_2 ANTENNA__12785__D (.DIODE(net482));
 sky130_fd_sc_hd__diode_2 ANTENNA__12786__A1 (.DIODE(net446));
 sky130_fd_sc_hd__diode_2 ANTENNA__12786__A2 (.DIODE(net486));
 sky130_fd_sc_hd__diode_2 ANTENNA__12786__B1 (.DIODE(net482));
 sky130_fd_sc_hd__diode_2 ANTENNA__12786__B2 (.DIODE(net452));
 sky130_fd_sc_hd__diode_2 ANTENNA__12828__A (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__12828__B (.DIODE(_04325_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12829__A1 (.DIODE(net599));
 sky130_fd_sc_hd__diode_2 ANTENNA__12829__B1 (.DIODE(_02745_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12829__B2 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__12830__S (.DIODE(_03055_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12839__B (.DIODE(net578));
 sky130_fd_sc_hd__diode_2 ANTENNA__12839__C (.DIODE(net360));
 sky130_fd_sc_hd__diode_2 ANTENNA__12839__D (.DIODE(net355));
 sky130_fd_sc_hd__diode_2 ANTENNA__12840__A2 (.DIODE(net360));
 sky130_fd_sc_hd__diode_2 ANTENNA__12840__B1 (.DIODE(net355));
 sky130_fd_sc_hd__diode_2 ANTENNA__12840__B2 (.DIODE(net578));
 sky130_fd_sc_hd__diode_2 ANTENNA__12842__C (.DIODE(net583));
 sky130_fd_sc_hd__diode_2 ANTENNA__12842__D (.DIODE(net348));
 sky130_fd_sc_hd__diode_2 ANTENNA__12843__A1_N (.DIODE(net583));
 sky130_fd_sc_hd__diode_2 ANTENNA__12843__A2_N (.DIODE(net348));
 sky130_fd_sc_hd__diode_2 ANTENNA__12845__A (.DIODE(net559));
 sky130_fd_sc_hd__diode_2 ANTENNA__12845__C (.DIODE(net631));
 sky130_fd_sc_hd__diode_2 ANTENNA__12845__D (.DIODE(net365));
 sky130_fd_sc_hd__diode_2 ANTENNA__12846__A1 (.DIODE(net559));
 sky130_fd_sc_hd__diode_2 ANTENNA__12846__A2 (.DIODE(net631));
 sky130_fd_sc_hd__diode_2 ANTENNA__12846__B1 (.DIODE(net365));
 sky130_fd_sc_hd__diode_2 ANTENNA__12848__C (.DIODE(net568));
 sky130_fd_sc_hd__diode_2 ANTENNA__12848__D (.DIODE(net364));
 sky130_fd_sc_hd__diode_2 ANTENNA__12849__A1_N (.DIODE(net568));
 sky130_fd_sc_hd__diode_2 ANTENNA__12849__A2_N (.DIODE(net364));
 sky130_fd_sc_hd__diode_2 ANTENNA__12857__A1 (.DIODE(net546));
 sky130_fd_sc_hd__diode_2 ANTENNA__12857__A2 (.DIODE(net389));
 sky130_fd_sc_hd__diode_2 ANTENNA__12857__B2 (.DIODE(net395));
 sky130_fd_sc_hd__diode_2 ANTENNA__12858__A (.DIODE(net546));
 sky130_fd_sc_hd__diode_2 ANTENNA__12858__B (.DIODE(net550));
 sky130_fd_sc_hd__diode_2 ANTENNA__12858__C (.DIODE(net381));
 sky130_fd_sc_hd__diode_2 ANTENNA__12859__A1 (.DIODE(net546));
 sky130_fd_sc_hd__diode_2 ANTENNA__12859__A2 (.DIODE(net382));
 sky130_fd_sc_hd__diode_2 ANTENNA__12859__B2 (.DIODE(net550));
 sky130_fd_sc_hd__diode_2 ANTENNA__12860__A (.DIODE(net554));
 sky130_fd_sc_hd__diode_2 ANTENNA__12860__B (.DIODE(net370));
 sky130_fd_sc_hd__diode_2 ANTENNA__12861__A1 (.DIODE(net554));
 sky130_fd_sc_hd__diode_2 ANTENNA__12861__A2 (.DIODE(net371));
 sky130_fd_sc_hd__diode_2 ANTENNA__12876__A (.DIODE(net542));
 sky130_fd_sc_hd__diode_2 ANTENNA__12876__B (.DIODE(net386));
 sky130_fd_sc_hd__diode_2 ANTENNA__12877__B (.DIODE(net535));
 sky130_fd_sc_hd__diode_2 ANTENNA__12878__A2 (.DIODE(net395));
 sky130_fd_sc_hd__diode_2 ANTENNA__12878__B2 (.DIODE(net535));
 sky130_fd_sc_hd__diode_2 ANTENNA__12879__A1 (.DIODE(net395));
 sky130_fd_sc_hd__diode_2 ANTENNA__12881__B (.DIODE(net401));
 sky130_fd_sc_hd__diode_2 ANTENNA__12882__A (.DIODE(net515));
 sky130_fd_sc_hd__diode_2 ANTENNA__12882__B (.DIODE(net521));
 sky130_fd_sc_hd__diode_2 ANTENNA__12882__C (.DIODE(net409));
 sky130_fd_sc_hd__diode_2 ANTENNA__12882__D (.DIODE(net405));
 sky130_fd_sc_hd__diode_2 ANTENNA__12883__A1 (.DIODE(net515));
 sky130_fd_sc_hd__diode_2 ANTENNA__12883__A2 (.DIODE(net409));
 sky130_fd_sc_hd__diode_2 ANTENNA__12883__B1 (.DIODE(net405));
 sky130_fd_sc_hd__diode_2 ANTENNA__12883__B2 (.DIODE(net521));
 sky130_fd_sc_hd__diode_2 ANTENNA__12886__A2 (.DIODE(net401));
 sky130_fd_sc_hd__diode_2 ANTENNA__12886__B2 (.DIODE(net409));
 sky130_fd_sc_hd__diode_2 ANTENNA__12897__A (.DIODE(\mul0.a[17] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__12897__B (.DIODE(net508));
 sky130_fd_sc_hd__diode_2 ANTENNA__12897__C (.DIODE(net422));
 sky130_fd_sc_hd__diode_2 ANTENNA__12897__D (.DIODE(net418));
 sky130_fd_sc_hd__diode_2 ANTENNA__12898__A1 (.DIODE(\mul0.a[17] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__12898__A2 (.DIODE(net422));
 sky130_fd_sc_hd__diode_2 ANTENNA__12898__B1 (.DIODE(net418));
 sky130_fd_sc_hd__diode_2 ANTENNA__12898__B2 (.DIODE(net508));
 sky130_fd_sc_hd__diode_2 ANTENNA__12899__A (.DIODE(net512));
 sky130_fd_sc_hd__diode_2 ANTENNA__12899__B (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA__12900__A1 (.DIODE(net512));
 sky130_fd_sc_hd__diode_2 ANTENNA__12900__A2 (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA__12905__A (.DIODE(net429));
 sky130_fd_sc_hd__diode_2 ANTENNA__12905__B (.DIODE(net498));
 sky130_fd_sc_hd__diode_2 ANTENNA__12906__A1 (.DIODE(net434));
 sky130_fd_sc_hd__diode_2 ANTENNA__12906__A2 (.DIODE(net494));
 sky130_fd_sc_hd__diode_2 ANTENNA__12906__B1 (.DIODE(net490));
 sky130_fd_sc_hd__diode_2 ANTENNA__12906__B2 (.DIODE(net439));
 sky130_fd_sc_hd__diode_2 ANTENNA__12907__A (.DIODE(net439));
 sky130_fd_sc_hd__diode_2 ANTENNA__12907__B (.DIODE(net434));
 sky130_fd_sc_hd__diode_2 ANTENNA__12907__C (.DIODE(net494));
 sky130_fd_sc_hd__diode_2 ANTENNA__12908__A1 (.DIODE(net490));
 sky130_fd_sc_hd__diode_2 ANTENNA__12910__A (.DIODE(net442));
 sky130_fd_sc_hd__diode_2 ANTENNA__12910__B (.DIODE(net486));
 sky130_fd_sc_hd__diode_2 ANTENNA__12911__A (.DIODE(net451));
 sky130_fd_sc_hd__diode_2 ANTENNA__12911__B (.DIODE(net447));
 sky130_fd_sc_hd__diode_2 ANTENNA__12911__C (.DIODE(net482));
 sky130_fd_sc_hd__diode_2 ANTENNA__12911__D (.DIODE(net478));
 sky130_fd_sc_hd__diode_2 ANTENNA__12912__A1 (.DIODE(net447));
 sky130_fd_sc_hd__diode_2 ANTENNA__12912__A2 (.DIODE(net482));
 sky130_fd_sc_hd__diode_2 ANTENNA__12912__B1 (.DIODE(net478));
 sky130_fd_sc_hd__diode_2 ANTENNA__12912__B2 (.DIODE(net451));
 sky130_fd_sc_hd__diode_2 ANTENNA__12953__A (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__12953__B (.DIODE(_04449_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12954__A1 (.DIODE(net599));
 sky130_fd_sc_hd__diode_2 ANTENNA__12954__B1 (.DIODE(_02746_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12954__B2 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__12962__B1 (.DIODE(net583));
 sky130_fd_sc_hd__diode_2 ANTENNA__12962__C1 (.DIODE(net344));
 sky130_fd_sc_hd__diode_2 ANTENNA__12963__A1 (.DIODE(net583));
 sky130_fd_sc_hd__diode_2 ANTENNA__12963__A2 (.DIODE(net344));
 sky130_fd_sc_hd__diode_2 ANTENNA__12973__A (.DIODE(net569));
 sky130_fd_sc_hd__diode_2 ANTENNA__12973__C (.DIODE(net360));
 sky130_fd_sc_hd__diode_2 ANTENNA__12973__D (.DIODE(net355));
 sky130_fd_sc_hd__diode_2 ANTENNA__12975__A1 (.DIODE(net568));
 sky130_fd_sc_hd__diode_2 ANTENNA__12975__A2 (.DIODE(net360));
 sky130_fd_sc_hd__diode_2 ANTENNA__12975__B1 (.DIODE(net355));
 sky130_fd_sc_hd__diode_2 ANTENNA__12976__A (.DIODE(net580));
 sky130_fd_sc_hd__diode_2 ANTENNA__12976__B (.DIODE(net348));
 sky130_fd_sc_hd__diode_2 ANTENNA__12977__A2 (.DIODE(net348));
 sky130_fd_sc_hd__diode_2 ANTENNA__12979__B (.DIODE(net364));
 sky130_fd_sc_hd__diode_2 ANTENNA__12980__A (.DIODE(net555));
 sky130_fd_sc_hd__diode_2 ANTENNA__12980__B (.DIODE(net559));
 sky130_fd_sc_hd__diode_2 ANTENNA__12980__C (.DIODE(net631));
 sky130_fd_sc_hd__diode_2 ANTENNA__12980__D (.DIODE(net365));
 sky130_fd_sc_hd__diode_2 ANTENNA__12981__A1 (.DIODE(net555));
 sky130_fd_sc_hd__diode_2 ANTENNA__12981__A2 (.DIODE(net631));
 sky130_fd_sc_hd__diode_2 ANTENNA__12981__B1 (.DIODE(net365));
 sky130_fd_sc_hd__diode_2 ANTENNA__12981__B2 (.DIODE(net559));
 sky130_fd_sc_hd__diode_2 ANTENNA__12990__A1 (.DIODE(net542));
 sky130_fd_sc_hd__diode_2 ANTENNA__12990__A2 (.DIODE(net386));
 sky130_fd_sc_hd__diode_2 ANTENNA__12990__B2 (.DIODE(net395));
 sky130_fd_sc_hd__diode_2 ANTENNA__12991__A (.DIODE(net542));
 sky130_fd_sc_hd__diode_2 ANTENNA__12991__B (.DIODE(net546));
 sky130_fd_sc_hd__diode_2 ANTENNA__12991__C (.DIODE(net382));
 sky130_fd_sc_hd__diode_2 ANTENNA__12991__D (.DIODE(net375));
 sky130_fd_sc_hd__diode_2 ANTENNA__12992__A1 (.DIODE(\mul0.a[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__12992__A2 (.DIODE(net382));
 sky130_fd_sc_hd__diode_2 ANTENNA__12992__B2 (.DIODE(net546));
 sky130_fd_sc_hd__diode_2 ANTENNA__12993__A (.DIODE(net550));
 sky130_fd_sc_hd__diode_2 ANTENNA__12993__B (.DIODE(net370));
 sky130_fd_sc_hd__diode_2 ANTENNA__12994__A1 (.DIODE(net550));
 sky130_fd_sc_hd__diode_2 ANTENNA__12994__A2 (.DIODE(net370));
 sky130_fd_sc_hd__diode_2 ANTENNA__13012__A (.DIODE(net537));
 sky130_fd_sc_hd__diode_2 ANTENNA__13012__B (.DIODE(net386));
 sky130_fd_sc_hd__diode_2 ANTENNA__13013__B (.DIODE(net532));
 sky130_fd_sc_hd__diode_2 ANTENNA__13014__A1 (.DIODE(net525));
 sky130_fd_sc_hd__diode_2 ANTENNA__13014__A2 (.DIODE(net395));
 sky130_fd_sc_hd__diode_2 ANTENNA__13014__B2 (.DIODE(net532));
 sky130_fd_sc_hd__diode_2 ANTENNA__13015__A1 (.DIODE(net395));
 sky130_fd_sc_hd__diode_2 ANTENNA__13017__A (.DIODE(net520));
 sky130_fd_sc_hd__diode_2 ANTENNA__13017__B (.DIODE(net401));
 sky130_fd_sc_hd__diode_2 ANTENNA__13018__A (.DIODE(net511));
 sky130_fd_sc_hd__diode_2 ANTENNA__13018__B (.DIODE(net516));
 sky130_fd_sc_hd__diode_2 ANTENNA__13018__C (.DIODE(net409));
 sky130_fd_sc_hd__diode_2 ANTENNA__13018__D (.DIODE(\mul0.b[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13019__A1 (.DIODE(net511));
 sky130_fd_sc_hd__diode_2 ANTENNA__13019__A2 (.DIODE(net409));
 sky130_fd_sc_hd__diode_2 ANTENNA__13019__B1 (.DIODE(\mul0.b[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13019__B2 (.DIODE(net516));
 sky130_fd_sc_hd__diode_2 ANTENNA__13033__A1 (.DIODE(net429));
 sky130_fd_sc_hd__diode_2 ANTENNA__13033__A2 (.DIODE(net498));
 sky130_fd_sc_hd__diode_2 ANTENNA__13033__B2 (.DIODE(net490));
 sky130_fd_sc_hd__diode_2 ANTENNA__13034__A (.DIODE(net503));
 sky130_fd_sc_hd__diode_2 ANTENNA__13034__B (.DIODE(net424));
 sky130_fd_sc_hd__diode_2 ANTENNA__13034__C (.DIODE(net420));
 sky130_fd_sc_hd__diode_2 ANTENNA__13034__D (.DIODE(net498));
 sky130_fd_sc_hd__diode_2 ANTENNA__13035__A1 (.DIODE(net503));
 sky130_fd_sc_hd__diode_2 ANTENNA__13035__A2 (.DIODE(net420));
 sky130_fd_sc_hd__diode_2 ANTENNA__13035__B1 (.DIODE(net498));
 sky130_fd_sc_hd__diode_2 ANTENNA__13035__B2 (.DIODE(net424));
 sky130_fd_sc_hd__diode_2 ANTENNA__13036__A (.DIODE(net508));
 sky130_fd_sc_hd__diode_2 ANTENNA__13036__B (.DIODE(net416));
 sky130_fd_sc_hd__diode_2 ANTENNA__13037__A1 (.DIODE(net508));
 sky130_fd_sc_hd__diode_2 ANTENNA__13037__A2 (.DIODE(net416));
 sky130_fd_sc_hd__diode_2 ANTENNA__13043__A (.DIODE(net429));
 sky130_fd_sc_hd__diode_2 ANTENNA__13043__B (.DIODE(net494));
 sky130_fd_sc_hd__diode_2 ANTENNA__13044__A (.DIODE(net439));
 sky130_fd_sc_hd__diode_2 ANTENNA__13044__B (.DIODE(net434));
 sky130_fd_sc_hd__diode_2 ANTENNA__13044__C (.DIODE(net490));
 sky130_fd_sc_hd__diode_2 ANTENNA__13044__D (.DIODE(net486));
 sky130_fd_sc_hd__diode_2 ANTENNA__13045__A1 (.DIODE(net434));
 sky130_fd_sc_hd__diode_2 ANTENNA__13045__A2 (.DIODE(net490));
 sky130_fd_sc_hd__diode_2 ANTENNA__13045__B1 (.DIODE(net486));
 sky130_fd_sc_hd__diode_2 ANTENNA__13045__B2 (.DIODE(net439));
 sky130_fd_sc_hd__diode_2 ANTENNA__13048__A (.DIODE(net442));
 sky130_fd_sc_hd__diode_2 ANTENNA__13048__B (.DIODE(net482));
 sky130_fd_sc_hd__diode_2 ANTENNA__13049__A (.DIODE(net451));
 sky130_fd_sc_hd__diode_2 ANTENNA__13049__B (.DIODE(net447));
 sky130_fd_sc_hd__diode_2 ANTENNA__13049__C (.DIODE(net478));
 sky130_fd_sc_hd__diode_2 ANTENNA__13049__D (.DIODE(net474));
 sky130_fd_sc_hd__diode_2 ANTENNA__13050__A1 (.DIODE(net447));
 sky130_fd_sc_hd__diode_2 ANTENNA__13050__A2 (.DIODE(net478));
 sky130_fd_sc_hd__diode_2 ANTENNA__13050__B1 (.DIODE(net474));
 sky130_fd_sc_hd__diode_2 ANTENNA__13050__B2 (.DIODE(net451));
 sky130_fd_sc_hd__diode_2 ANTENNA__13093__A (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__13093__B (.DIODE(_04588_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13094__A1 (.DIODE(net600));
 sky130_fd_sc_hd__diode_2 ANTENNA__13094__B1 (.DIODE(_02747_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13094__B2 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__13095__S (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__13098__A2 (.DIODE(net344));
 sky130_fd_sc_hd__diode_2 ANTENNA__13098__B2 (.DIODE(net583));
 sky130_fd_sc_hd__diode_2 ANTENNA__13099__B (.DIODE(net583));
 sky130_fd_sc_hd__diode_2 ANTENNA__13099__C (.DIODE(net344));
 sky130_fd_sc_hd__diode_2 ANTENNA__13113__B (.DIODE(net569));
 sky130_fd_sc_hd__diode_2 ANTENNA__13113__C (.DIODE(net356));
 sky130_fd_sc_hd__diode_2 ANTENNA__13113__D (.DIODE(net355));
 sky130_fd_sc_hd__diode_2 ANTENNA__13114__A2 (.DIODE(net356));
 sky130_fd_sc_hd__diode_2 ANTENNA__13114__B1 (.DIODE(net355));
 sky130_fd_sc_hd__diode_2 ANTENNA__13114__B2 (.DIODE(net569));
 sky130_fd_sc_hd__diode_2 ANTENNA__13116__A (.DIODE(net574));
 sky130_fd_sc_hd__diode_2 ANTENNA__13116__B (.DIODE(net348));
 sky130_fd_sc_hd__diode_2 ANTENNA__13118__A (.DIODE(net559));
 sky130_fd_sc_hd__diode_2 ANTENNA__13118__B (.DIODE(net364));
 sky130_fd_sc_hd__diode_2 ANTENNA__13119__A (.DIODE(net551));
 sky130_fd_sc_hd__diode_2 ANTENNA__13119__B (.DIODE(net555));
 sky130_fd_sc_hd__diode_2 ANTENNA__13119__C (.DIODE(\mul0.b[18] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13119__D (.DIODE(\mul0.b[19] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13120__A1 (.DIODE(net551));
 sky130_fd_sc_hd__diode_2 ANTENNA__13120__A2 (.DIODE(\mul0.b[18] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13120__B1 (.DIODE(net365));
 sky130_fd_sc_hd__diode_2 ANTENNA__13120__B2 (.DIODE(net555));
 sky130_fd_sc_hd__diode_2 ANTENNA__13123__A2 (.DIODE(net364));
 sky130_fd_sc_hd__diode_2 ANTENNA__13129__A1 (.DIODE(net537));
 sky130_fd_sc_hd__diode_2 ANTENNA__13129__A2 (.DIODE(net389));
 sky130_fd_sc_hd__diode_2 ANTENNA__13129__B2 (.DIODE(net395));
 sky130_fd_sc_hd__diode_2 ANTENNA__13130__A (.DIODE(net537));
 sky130_fd_sc_hd__diode_2 ANTENNA__13130__B (.DIODE(net542));
 sky130_fd_sc_hd__diode_2 ANTENNA__13130__C (.DIODE(net382));
 sky130_fd_sc_hd__diode_2 ANTENNA__13131__A1 (.DIODE(net537));
 sky130_fd_sc_hd__diode_2 ANTENNA__13131__A2 (.DIODE(net382));
 sky130_fd_sc_hd__diode_2 ANTENNA__13131__B2 (.DIODE(net542));
 sky130_fd_sc_hd__diode_2 ANTENNA__13132__A (.DIODE(net546));
 sky130_fd_sc_hd__diode_2 ANTENNA__13132__B (.DIODE(net370));
 sky130_fd_sc_hd__diode_2 ANTENNA__13133__A1 (.DIODE(net546));
 sky130_fd_sc_hd__diode_2 ANTENNA__13133__A2 (.DIODE(net370));
 sky130_fd_sc_hd__diode_2 ANTENNA__13150__A (.DIODE(net532));
 sky130_fd_sc_hd__diode_2 ANTENNA__13150__B (.DIODE(net387));
 sky130_fd_sc_hd__diode_2 ANTENNA__13151__A1 (.DIODE(net521));
 sky130_fd_sc_hd__diode_2 ANTENNA__13151__A2 (.DIODE(net395));
 sky130_fd_sc_hd__diode_2 ANTENNA__13151__B1 (.DIODE(net390));
 sky130_fd_sc_hd__diode_2 ANTENNA__13151__B2 (.DIODE(net527));
 sky130_fd_sc_hd__diode_2 ANTENNA__13152__A (.DIODE(net521));
 sky130_fd_sc_hd__diode_2 ANTENNA__13152__B (.DIODE(net527));
 sky130_fd_sc_hd__diode_2 ANTENNA__13152__C (.DIODE(net395));
 sky130_fd_sc_hd__diode_2 ANTENNA__13155__A (.DIODE(net507));
 sky130_fd_sc_hd__diode_2 ANTENNA__13155__B (.DIODE(net511));
 sky130_fd_sc_hd__diode_2 ANTENNA__13155__C (.DIODE(net409));
 sky130_fd_sc_hd__diode_2 ANTENNA__13155__D (.DIODE(net405));
 sky130_fd_sc_hd__diode_2 ANTENNA__13156__A1 (.DIODE(net507));
 sky130_fd_sc_hd__diode_2 ANTENNA__13156__A2 (.DIODE(net409));
 sky130_fd_sc_hd__diode_2 ANTENNA__13156__B1 (.DIODE(net405));
 sky130_fd_sc_hd__diode_2 ANTENNA__13156__B2 (.DIODE(net511));
 sky130_fd_sc_hd__diode_2 ANTENNA__13157__A (.DIODE(net515));
 sky130_fd_sc_hd__diode_2 ANTENNA__13157__B (.DIODE(net401));
 sky130_fd_sc_hd__diode_2 ANTENNA__13158__A1 (.DIODE(net515));
 sky130_fd_sc_hd__diode_2 ANTENNA__13158__A2 (.DIODE(net401));
 sky130_fd_sc_hd__diode_2 ANTENNA__13171__A1 (.DIODE(net420));
 sky130_fd_sc_hd__diode_2 ANTENNA__13171__A2 (.DIODE(net498));
 sky130_fd_sc_hd__diode_2 ANTENNA__13171__B1 (.DIODE(net494));
 sky130_fd_sc_hd__diode_2 ANTENNA__13171__B2 (.DIODE(net424));
 sky130_fd_sc_hd__diode_2 ANTENNA__13172__A (.DIODE(net424));
 sky130_fd_sc_hd__diode_2 ANTENNA__13172__B (.DIODE(net420));
 sky130_fd_sc_hd__diode_2 ANTENNA__13172__C (.DIODE(net499));
 sky130_fd_sc_hd__diode_2 ANTENNA__13172__D (.DIODE(net494));
 sky130_fd_sc_hd__diode_2 ANTENNA__13173__C (.DIODE(net503));
 sky130_fd_sc_hd__diode_2 ANTENNA__13173__D (.DIODE(net416));
 sky130_fd_sc_hd__diode_2 ANTENNA__13174__A1_N (.DIODE(net503));
 sky130_fd_sc_hd__diode_2 ANTENNA__13174__A2_N (.DIODE(net416));
 sky130_fd_sc_hd__diode_2 ANTENNA__13180__A (.DIODE(net429));
 sky130_fd_sc_hd__diode_2 ANTENNA__13180__B (.DIODE(net490));
 sky130_fd_sc_hd__diode_2 ANTENNA__13181__A (.DIODE(net439));
 sky130_fd_sc_hd__diode_2 ANTENNA__13181__B (.DIODE(net434));
 sky130_fd_sc_hd__diode_2 ANTENNA__13181__C (.DIODE(net486));
 sky130_fd_sc_hd__diode_2 ANTENNA__13181__D (.DIODE(net482));
 sky130_fd_sc_hd__diode_2 ANTENNA__13182__A1 (.DIODE(net434));
 sky130_fd_sc_hd__diode_2 ANTENNA__13182__A2 (.DIODE(net486));
 sky130_fd_sc_hd__diode_2 ANTENNA__13182__B1 (.DIODE(net482));
 sky130_fd_sc_hd__diode_2 ANTENNA__13182__B2 (.DIODE(net439));
 sky130_fd_sc_hd__diode_2 ANTENNA__13185__A (.DIODE(net442));
 sky130_fd_sc_hd__diode_2 ANTENNA__13185__B (.DIODE(net478));
 sky130_fd_sc_hd__diode_2 ANTENNA__13186__A (.DIODE(net451));
 sky130_fd_sc_hd__diode_2 ANTENNA__13186__B (.DIODE(net447));
 sky130_fd_sc_hd__diode_2 ANTENNA__13186__C (.DIODE(net474));
 sky130_fd_sc_hd__diode_2 ANTENNA__13186__D (.DIODE(net470));
 sky130_fd_sc_hd__diode_2 ANTENNA__13187__A1 (.DIODE(net447));
 sky130_fd_sc_hd__diode_2 ANTENNA__13187__A2 (.DIODE(net474));
 sky130_fd_sc_hd__diode_2 ANTENNA__13187__B1 (.DIODE(net470));
 sky130_fd_sc_hd__diode_2 ANTENNA__13187__B2 (.DIODE(net451));
 sky130_fd_sc_hd__diode_2 ANTENNA__13225__A (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__13225__B (.DIODE(_04719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13226__A1 (.DIODE(net599));
 sky130_fd_sc_hd__diode_2 ANTENNA__13226__B1 (.DIODE(_02748_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13226__B2 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__13232__A2 (.DIODE(net348));
 sky130_fd_sc_hd__diode_2 ANTENNA__13233__C (.DIODE(net344));
 sky130_fd_sc_hd__diode_2 ANTENNA__13234__A2 (.DIODE(net344));
 sky130_fd_sc_hd__diode_2 ANTENNA__13235__C (.DIODE(net583));
 sky130_fd_sc_hd__diode_2 ANTENNA__13235__D (.DIODE(net337));
 sky130_fd_sc_hd__diode_2 ANTENNA__13236__A1_N (.DIODE(net583));
 sky130_fd_sc_hd__diode_2 ANTENNA__13236__A2_N (.DIODE(net337));
 sky130_fd_sc_hd__diode_2 ANTENNA__13253__A1 (.DIODE(net559));
 sky130_fd_sc_hd__diode_2 ANTENNA__13253__A2 (.DIODE(net356));
 sky130_fd_sc_hd__diode_2 ANTENNA__13253__B1 (.DIODE(net355));
 sky130_fd_sc_hd__diode_2 ANTENNA__13253__B2 (.DIODE(net563));
 sky130_fd_sc_hd__diode_2 ANTENNA__13254__A (.DIODE(net559));
 sky130_fd_sc_hd__diode_2 ANTENNA__13254__B (.DIODE(net563));
 sky130_fd_sc_hd__diode_2 ANTENNA__13254__C (.DIODE(net355));
 sky130_fd_sc_hd__diode_2 ANTENNA__13255__A1 (.DIODE(net356));
 sky130_fd_sc_hd__diode_2 ANTENNA__13256__A (.DIODE(net569));
 sky130_fd_sc_hd__diode_2 ANTENNA__13256__B (.DIODE(net348));
 sky130_fd_sc_hd__diode_2 ANTENNA__13258__A (.DIODE(net546));
 sky130_fd_sc_hd__diode_2 ANTENNA__13258__B (.DIODE(net550));
 sky130_fd_sc_hd__diode_2 ANTENNA__13258__C (.DIODE(net631));
 sky130_fd_sc_hd__diode_2 ANTENNA__13258__D (.DIODE(net365));
 sky130_fd_sc_hd__diode_2 ANTENNA__13259__A1 (.DIODE(net546));
 sky130_fd_sc_hd__diode_2 ANTENNA__13259__A2 (.DIODE(net631));
 sky130_fd_sc_hd__diode_2 ANTENNA__13259__B1 (.DIODE(net365));
 sky130_fd_sc_hd__diode_2 ANTENNA__13259__B2 (.DIODE(net550));
 sky130_fd_sc_hd__diode_2 ANTENNA__13260__A (.DIODE(net554));
 sky130_fd_sc_hd__diode_2 ANTENNA__13260__B (.DIODE(net364));
 sky130_fd_sc_hd__diode_2 ANTENNA__13261__A1 (.DIODE(net554));
 sky130_fd_sc_hd__diode_2 ANTENNA__13261__A2 (.DIODE(net364));
 sky130_fd_sc_hd__diode_2 ANTENNA__13269__A (.DIODE(net532));
 sky130_fd_sc_hd__diode_2 ANTENNA__13269__B (.DIODE(net537));
 sky130_fd_sc_hd__diode_2 ANTENNA__13269__C (.DIODE(net382));
 sky130_fd_sc_hd__diode_2 ANTENNA__13270__A1 (.DIODE(net532));
 sky130_fd_sc_hd__diode_2 ANTENNA__13270__A2 (.DIODE(net382));
 sky130_fd_sc_hd__diode_2 ANTENNA__13270__B2 (.DIODE(net537));
 sky130_fd_sc_hd__diode_2 ANTENNA__13271__C (.DIODE(net542));
 sky130_fd_sc_hd__diode_2 ANTENNA__13271__D (.DIODE(net370));
 sky130_fd_sc_hd__diode_2 ANTENNA__13272__A1_N (.DIODE(net542));
 sky130_fd_sc_hd__diode_2 ANTENNA__13272__A2_N (.DIODE(net370));
 sky130_fd_sc_hd__diode_2 ANTENNA__13288__A1 (.DIODE(net517));
 sky130_fd_sc_hd__diode_2 ANTENNA__13288__A2 (.DIODE(net397));
 sky130_fd_sc_hd__diode_2 ANTENNA__13288__B1 (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA__13288__B2 (.DIODE(net524));
 sky130_fd_sc_hd__diode_2 ANTENNA__13289__A (.DIODE(net517));
 sky130_fd_sc_hd__diode_2 ANTENNA__13289__B (.DIODE(net521));
 sky130_fd_sc_hd__diode_2 ANTENNA__13289__C (.DIODE(net397));
 sky130_fd_sc_hd__diode_2 ANTENNA__13289__D (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA__13290__A (.DIODE(net527));
 sky130_fd_sc_hd__diode_2 ANTENNA__13290__B (.DIODE(net387));
 sky130_fd_sc_hd__diode_2 ANTENNA__13291__A1 (.DIODE(net527));
 sky130_fd_sc_hd__diode_2 ANTENNA__13291__A2 (.DIODE(net387));
 sky130_fd_sc_hd__diode_2 ANTENNA__13293__A1 (.DIODE(net504));
 sky130_fd_sc_hd__diode_2 ANTENNA__13293__A2 (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA__13293__B1 (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA__13293__B2 (.DIODE(net508));
 sky130_fd_sc_hd__diode_2 ANTENNA__13294__A (.DIODE(net504));
 sky130_fd_sc_hd__diode_2 ANTENNA__13294__B (.DIODE(net508));
 sky130_fd_sc_hd__diode_2 ANTENNA__13294__C (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA__13294__D (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA__13295__C (.DIODE(net512));
 sky130_fd_sc_hd__diode_2 ANTENNA__13295__D (.DIODE(net403));
 sky130_fd_sc_hd__diode_2 ANTENNA__13296__A1_N (.DIODE(net512));
 sky130_fd_sc_hd__diode_2 ANTENNA__13296__A2_N (.DIODE(net403));
 sky130_fd_sc_hd__diode_2 ANTENNA__13310__A1 (.DIODE(net420));
 sky130_fd_sc_hd__diode_2 ANTENNA__13310__A2 (.DIODE(net494));
 sky130_fd_sc_hd__diode_2 ANTENNA__13310__B1 (.DIODE(net490));
 sky130_fd_sc_hd__diode_2 ANTENNA__13310__B2 (.DIODE(net424));
 sky130_fd_sc_hd__diode_2 ANTENNA__13311__A (.DIODE(net424));
 sky130_fd_sc_hd__diode_2 ANTENNA__13311__B (.DIODE(net420));
 sky130_fd_sc_hd__diode_2 ANTENNA__13311__C (.DIODE(net494));
 sky130_fd_sc_hd__diode_2 ANTENNA__13311__D (.DIODE(net490));
 sky130_fd_sc_hd__diode_2 ANTENNA__13312__C (.DIODE(net416));
 sky130_fd_sc_hd__diode_2 ANTENNA__13312__D (.DIODE(net499));
 sky130_fd_sc_hd__diode_2 ANTENNA__13313__A1_N (.DIODE(net416));
 sky130_fd_sc_hd__diode_2 ANTENNA__13313__A2_N (.DIODE(net498));
 sky130_fd_sc_hd__diode_2 ANTENNA__13319__A (.DIODE(net429));
 sky130_fd_sc_hd__diode_2 ANTENNA__13319__B (.DIODE(net486));
 sky130_fd_sc_hd__diode_2 ANTENNA__13320__A (.DIODE(net439));
 sky130_fd_sc_hd__diode_2 ANTENNA__13320__B (.DIODE(net434));
 sky130_fd_sc_hd__diode_2 ANTENNA__13320__C (.DIODE(net482));
 sky130_fd_sc_hd__diode_2 ANTENNA__13320__D (.DIODE(net478));
 sky130_fd_sc_hd__diode_2 ANTENNA__13321__A1 (.DIODE(net434));
 sky130_fd_sc_hd__diode_2 ANTENNA__13321__A2 (.DIODE(net482));
 sky130_fd_sc_hd__diode_2 ANTENNA__13321__B1 (.DIODE(net478));
 sky130_fd_sc_hd__diode_2 ANTENNA__13321__B2 (.DIODE(net439));
 sky130_fd_sc_hd__diode_2 ANTENNA__13324__A (.DIODE(net442));
 sky130_fd_sc_hd__diode_2 ANTENNA__13324__B (.DIODE(net474));
 sky130_fd_sc_hd__diode_2 ANTENNA__13325__A (.DIODE(net451));
 sky130_fd_sc_hd__diode_2 ANTENNA__13325__B (.DIODE(net447));
 sky130_fd_sc_hd__diode_2 ANTENNA__13325__C (.DIODE(net470));
 sky130_fd_sc_hd__diode_2 ANTENNA__13325__D (.DIODE(net466));
 sky130_fd_sc_hd__diode_2 ANTENNA__13326__A1 (.DIODE(net447));
 sky130_fd_sc_hd__diode_2 ANTENNA__13326__A2 (.DIODE(net470));
 sky130_fd_sc_hd__diode_2 ANTENNA__13326__B1 (.DIODE(net466));
 sky130_fd_sc_hd__diode_2 ANTENNA__13326__B2 (.DIODE(net451));
 sky130_fd_sc_hd__diode_2 ANTENNA__13369__A (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__13369__B (.DIODE(_04862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13370__A1 (.DIODE(net600));
 sky130_fd_sc_hd__diode_2 ANTENNA__13370__B1 (.DIODE(_02749_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13370__B2 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__13377__A1 (.DIODE(net568));
 sky130_fd_sc_hd__diode_2 ANTENNA__13377__A2 (.DIODE(net348));
 sky130_fd_sc_hd__diode_2 ANTENNA__13377__B2 (.DIODE(net356));
 sky130_fd_sc_hd__diode_2 ANTENNA__13378__A1 (.DIODE(net568));
 sky130_fd_sc_hd__diode_2 ANTENNA__13378__A2 (.DIODE(net344));
 sky130_fd_sc_hd__diode_2 ANTENNA__13379__A (.DIODE(net568));
 sky130_fd_sc_hd__diode_2 ANTENNA__13379__C (.DIODE(net344));
 sky130_fd_sc_hd__diode_2 ANTENNA__13380__A2_N (.DIODE(net337));
 sky130_fd_sc_hd__diode_2 ANTENNA__13381__D (.DIODE(net337));
 sky130_fd_sc_hd__diode_2 ANTENNA__13394__A (.DIODE(net583));
 sky130_fd_sc_hd__diode_2 ANTENNA__13394__B (.DIODE(net336));
 sky130_fd_sc_hd__diode_2 ANTENNA__13401__A1 (.DIODE(net554));
 sky130_fd_sc_hd__diode_2 ANTENNA__13401__A2 (.DIODE(net356));
 sky130_fd_sc_hd__diode_2 ANTENNA__13401__B1 (.DIODE(net355));
 sky130_fd_sc_hd__diode_2 ANTENNA__13401__B2 (.DIODE(net558));
 sky130_fd_sc_hd__diode_2 ANTENNA__13402__A (.DIODE(net554));
 sky130_fd_sc_hd__diode_2 ANTENNA__13402__B (.DIODE(net558));
 sky130_fd_sc_hd__diode_2 ANTENNA__13402__C (.DIODE(net356));
 sky130_fd_sc_hd__diode_2 ANTENNA__13402__D (.DIODE(net355));
 sky130_fd_sc_hd__diode_2 ANTENNA__13403__A1 (.DIODE(net563));
 sky130_fd_sc_hd__diode_2 ANTENNA__13403__A2 (.DIODE(\mul0.b[23] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13404__A (.DIODE(net563));
 sky130_fd_sc_hd__diode_2 ANTENNA__13404__B (.DIODE(net348));
 sky130_fd_sc_hd__diode_2 ANTENNA__13406__A (.DIODE(net550));
 sky130_fd_sc_hd__diode_2 ANTENNA__13406__B (.DIODE(net364));
 sky130_fd_sc_hd__diode_2 ANTENNA__13407__A1 (.DIODE(net542));
 sky130_fd_sc_hd__diode_2 ANTENNA__13407__A2 (.DIODE(net632));
 sky130_fd_sc_hd__diode_2 ANTENNA__13407__B1 (.DIODE(net367));
 sky130_fd_sc_hd__diode_2 ANTENNA__13407__B2 (.DIODE(\mul0.a[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13408__A (.DIODE(net542));
 sky130_fd_sc_hd__diode_2 ANTENNA__13408__B (.DIODE(net546));
 sky130_fd_sc_hd__diode_2 ANTENNA__13408__C (.DIODE(net632));
 sky130_fd_sc_hd__diode_2 ANTENNA__13408__D (.DIODE(net367));
 sky130_fd_sc_hd__diode_2 ANTENNA__13417__A1 (.DIODE(net527));
 sky130_fd_sc_hd__diode_2 ANTENNA__13417__A2 (.DIODE(net383));
 sky130_fd_sc_hd__diode_2 ANTENNA__13417__B1 (.DIODE(net377));
 sky130_fd_sc_hd__diode_2 ANTENNA__13417__B2 (.DIODE(net532));
 sky130_fd_sc_hd__diode_2 ANTENNA__13418__A (.DIODE(net527));
 sky130_fd_sc_hd__diode_2 ANTENNA__13418__B (.DIODE(net532));
 sky130_fd_sc_hd__diode_2 ANTENNA__13418__C (.DIODE(net383));
 sky130_fd_sc_hd__diode_2 ANTENNA__13418__D (.DIODE(net377));
 sky130_fd_sc_hd__diode_2 ANTENNA__13419__A1_N (.DIODE(net537));
 sky130_fd_sc_hd__diode_2 ANTENNA__13419__A2_N (.DIODE(net370));
 sky130_fd_sc_hd__diode_2 ANTENNA__13420__C (.DIODE(net537));
 sky130_fd_sc_hd__diode_2 ANTENNA__13420__D (.DIODE(net370));
 sky130_fd_sc_hd__diode_2 ANTENNA__13435__A1 (.DIODE(net512));
 sky130_fd_sc_hd__diode_2 ANTENNA__13435__A2 (.DIODE(net397));
 sky130_fd_sc_hd__diode_2 ANTENNA__13435__B1 (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA__13435__B2 (.DIODE(net517));
 sky130_fd_sc_hd__diode_2 ANTENNA__13436__A (.DIODE(net512));
 sky130_fd_sc_hd__diode_2 ANTENNA__13436__B (.DIODE(net517));
 sky130_fd_sc_hd__diode_2 ANTENNA__13436__C (.DIODE(net397));
 sky130_fd_sc_hd__diode_2 ANTENNA__13436__D (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA__13437__A (.DIODE(net521));
 sky130_fd_sc_hd__diode_2 ANTENNA__13437__B (.DIODE(net387));
 sky130_fd_sc_hd__diode_2 ANTENNA__13438__A1 (.DIODE(net521));
 sky130_fd_sc_hd__diode_2 ANTENNA__13438__A2 (.DIODE(net387));
 sky130_fd_sc_hd__diode_2 ANTENNA__13440__A (.DIODE(net508));
 sky130_fd_sc_hd__diode_2 ANTENNA__13440__B (.DIODE(net403));
 sky130_fd_sc_hd__diode_2 ANTENNA__13441__A1 (.DIODE(net504));
 sky130_fd_sc_hd__diode_2 ANTENNA__13441__A2 (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA__13441__B1 (.DIODE(net499));
 sky130_fd_sc_hd__diode_2 ANTENNA__13441__B2 (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA__13442__A (.DIODE(net504));
 sky130_fd_sc_hd__diode_2 ANTENNA__13442__B (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA__13442__C (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA__13442__D (.DIODE(net499));
 sky130_fd_sc_hd__diode_2 ANTENNA__13456__A1 (.DIODE(net429));
 sky130_fd_sc_hd__diode_2 ANTENNA__13456__A2 (.DIODE(net486));
 sky130_fd_sc_hd__diode_2 ANTENNA__13457__A1 (.DIODE(net420));
 sky130_fd_sc_hd__diode_2 ANTENNA__13457__A2 (.DIODE(net491));
 sky130_fd_sc_hd__diode_2 ANTENNA__13457__B1 (.DIODE(net486));
 sky130_fd_sc_hd__diode_2 ANTENNA__13457__B2 (.DIODE(net424));
 sky130_fd_sc_hd__diode_2 ANTENNA__13458__A (.DIODE(net424));
 sky130_fd_sc_hd__diode_2 ANTENNA__13458__B (.DIODE(net420));
 sky130_fd_sc_hd__diode_2 ANTENNA__13458__C (.DIODE(net491));
 sky130_fd_sc_hd__diode_2 ANTENNA__13458__D (.DIODE(net487));
 sky130_fd_sc_hd__diode_2 ANTENNA__13459__A (.DIODE(net424));
 sky130_fd_sc_hd__diode_2 ANTENNA__13459__B (.DIODE(net420));
 sky130_fd_sc_hd__diode_2 ANTENNA__13459__C (.DIODE(net491));
 sky130_fd_sc_hd__diode_2 ANTENNA__13459__D (.DIODE(net486));
 sky130_fd_sc_hd__diode_2 ANTENNA__13460__A1 (.DIODE(net416));
 sky130_fd_sc_hd__diode_2 ANTENNA__13460__A2 (.DIODE(net495));
 sky130_fd_sc_hd__diode_2 ANTENNA__13461__A (.DIODE(net416));
 sky130_fd_sc_hd__diode_2 ANTENNA__13461__B (.DIODE(net495));
 sky130_fd_sc_hd__diode_2 ANTENNA__13467__A (.DIODE(net428));
 sky130_fd_sc_hd__diode_2 ANTENNA__13467__B (.DIODE(net482));
 sky130_fd_sc_hd__diode_2 ANTENNA__13468__A (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA__13468__B (.DIODE(net433));
 sky130_fd_sc_hd__diode_2 ANTENNA__13468__C (.DIODE(net478));
 sky130_fd_sc_hd__diode_2 ANTENNA__13468__D (.DIODE(net474));
 sky130_fd_sc_hd__diode_2 ANTENNA__13469__A1 (.DIODE(net433));
 sky130_fd_sc_hd__diode_2 ANTENNA__13469__A2 (.DIODE(net478));
 sky130_fd_sc_hd__diode_2 ANTENNA__13469__B1 (.DIODE(net474));
 sky130_fd_sc_hd__diode_2 ANTENNA__13469__B2 (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA__13472__A (.DIODE(net442));
 sky130_fd_sc_hd__diode_2 ANTENNA__13472__B (.DIODE(net470));
 sky130_fd_sc_hd__diode_2 ANTENNA__13473__A (.DIODE(net451));
 sky130_fd_sc_hd__diode_2 ANTENNA__13473__B (.DIODE(net447));
 sky130_fd_sc_hd__diode_2 ANTENNA__13473__C (.DIODE(net466));
 sky130_fd_sc_hd__diode_2 ANTENNA__13473__D (.DIODE(net463));
 sky130_fd_sc_hd__diode_2 ANTENNA__13474__A1 (.DIODE(net447));
 sky130_fd_sc_hd__diode_2 ANTENNA__13474__A2 (.DIODE(net466));
 sky130_fd_sc_hd__diode_2 ANTENNA__13474__B1 (.DIODE(net463));
 sky130_fd_sc_hd__diode_2 ANTENNA__13474__B2 (.DIODE(net451));
 sky130_fd_sc_hd__diode_2 ANTENNA__13514__A (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__13514__B (.DIODE(_05006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13515__A1 (.DIODE(net600));
 sky130_fd_sc_hd__diode_2 ANTENNA__13515__B1 (.DIODE(_02751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13515__B2 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__13516__S (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__13524__A1 (.DIODE(net580));
 sky130_fd_sc_hd__diode_2 ANTENNA__13524__A2 (.DIODE(net336));
 sky130_fd_sc_hd__diode_2 ANTENNA__13524__B1 (.DIODE(net333));
 sky130_fd_sc_hd__diode_2 ANTENNA__13524__B2 (.DIODE(net583));
 sky130_fd_sc_hd__diode_2 ANTENNA__13525__A (.DIODE(net580));
 sky130_fd_sc_hd__diode_2 ANTENNA__13525__B (.DIODE(net584));
 sky130_fd_sc_hd__diode_2 ANTENNA__13525__C (.DIODE(net336));
 sky130_fd_sc_hd__diode_2 ANTENNA__13525__D (.DIODE(net333));
 sky130_fd_sc_hd__diode_2 ANTENNA__13528__A2 (.DIODE(net344));
 sky130_fd_sc_hd__diode_2 ANTENNA__13528__B2 (.DIODE(net568));
 sky130_fd_sc_hd__diode_2 ANTENNA__13529__B (.DIODE(net568));
 sky130_fd_sc_hd__diode_2 ANTENNA__13529__C (.DIODE(net344));
 sky130_fd_sc_hd__diode_2 ANTENNA__13530__A2_N (.DIODE(net337));
 sky130_fd_sc_hd__diode_2 ANTENNA__13531__D (.DIODE(net337));
 sky130_fd_sc_hd__diode_2 ANTENNA__13553__A1 (.DIODE(net550));
 sky130_fd_sc_hd__diode_2 ANTENNA__13553__A2 (.DIODE(net356));
 sky130_fd_sc_hd__diode_2 ANTENNA__13553__B1 (.DIODE(net355));
 sky130_fd_sc_hd__diode_2 ANTENNA__13553__B2 (.DIODE(net554));
 sky130_fd_sc_hd__diode_2 ANTENNA__13554__A (.DIODE(net550));
 sky130_fd_sc_hd__diode_2 ANTENNA__13554__B (.DIODE(net554));
 sky130_fd_sc_hd__diode_2 ANTENNA__13554__C (.DIODE(net356));
 sky130_fd_sc_hd__diode_2 ANTENNA__13554__D (.DIODE(net354));
 sky130_fd_sc_hd__diode_2 ANTENNA__13555__A1 (.DIODE(net558));
 sky130_fd_sc_hd__diode_2 ANTENNA__13555__A2 (.DIODE(net348));
 sky130_fd_sc_hd__diode_2 ANTENNA__13556__A (.DIODE(net558));
 sky130_fd_sc_hd__diode_2 ANTENNA__13556__B (.DIODE(net348));
 sky130_fd_sc_hd__diode_2 ANTENNA__13558__A1 (.DIODE(net537));
 sky130_fd_sc_hd__diode_2 ANTENNA__13558__A2 (.DIODE(net632));
 sky130_fd_sc_hd__diode_2 ANTENNA__13558__B1 (.DIODE(net367));
 sky130_fd_sc_hd__diode_2 ANTENNA__13558__B2 (.DIODE(net542));
 sky130_fd_sc_hd__diode_2 ANTENNA__13559__A (.DIODE(net537));
 sky130_fd_sc_hd__diode_2 ANTENNA__13559__B (.DIODE(net542));
 sky130_fd_sc_hd__diode_2 ANTENNA__13559__C (.DIODE(net632));
 sky130_fd_sc_hd__diode_2 ANTENNA__13559__D (.DIODE(net367));
 sky130_fd_sc_hd__diode_2 ANTENNA__13560__A1_N (.DIODE(net546));
 sky130_fd_sc_hd__diode_2 ANTENNA__13560__A2_N (.DIODE(net363));
 sky130_fd_sc_hd__diode_2 ANTENNA__13561__C (.DIODE(\mul0.a[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13561__D (.DIODE(net363));
 sky130_fd_sc_hd__diode_2 ANTENNA__13570__A1 (.DIODE(net521));
 sky130_fd_sc_hd__diode_2 ANTENNA__13570__A2 (.DIODE(net383));
 sky130_fd_sc_hd__diode_2 ANTENNA__13570__B1 (.DIODE(net377));
 sky130_fd_sc_hd__diode_2 ANTENNA__13570__B2 (.DIODE(net527));
 sky130_fd_sc_hd__diode_2 ANTENNA__13571__A (.DIODE(net524));
 sky130_fd_sc_hd__diode_2 ANTENNA__13571__B (.DIODE(net527));
 sky130_fd_sc_hd__diode_2 ANTENNA__13571__C (.DIODE(net383));
 sky130_fd_sc_hd__diode_2 ANTENNA__13571__D (.DIODE(net377));
 sky130_fd_sc_hd__diode_2 ANTENNA__13572__A1_N (.DIODE(net532));
 sky130_fd_sc_hd__diode_2 ANTENNA__13572__A2_N (.DIODE(net374));
 sky130_fd_sc_hd__diode_2 ANTENNA__13573__C (.DIODE(net532));
 sky130_fd_sc_hd__diode_2 ANTENNA__13573__D (.DIODE(net370));
 sky130_fd_sc_hd__diode_2 ANTENNA__13588__A1 (.DIODE(net508));
 sky130_fd_sc_hd__diode_2 ANTENNA__13588__A2 (.DIODE(net397));
 sky130_fd_sc_hd__diode_2 ANTENNA__13588__B1 (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA__13588__B2 (.DIODE(net512));
 sky130_fd_sc_hd__diode_2 ANTENNA__13589__A (.DIODE(\mul0.a[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13589__B (.DIODE(net512));
 sky130_fd_sc_hd__diode_2 ANTENNA__13589__C (.DIODE(net397));
 sky130_fd_sc_hd__diode_2 ANTENNA__13589__D (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA__13590__A1 (.DIODE(net517));
 sky130_fd_sc_hd__diode_2 ANTENNA__13590__A2 (.DIODE(net387));
 sky130_fd_sc_hd__diode_2 ANTENNA__13591__A (.DIODE(net517));
 sky130_fd_sc_hd__diode_2 ANTENNA__13591__B (.DIODE(net387));
 sky130_fd_sc_hd__diode_2 ANTENNA__13593__A1 (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA__13593__A2 (.DIODE(net499));
 sky130_fd_sc_hd__diode_2 ANTENNA__13593__B1 (.DIODE(net495));
 sky130_fd_sc_hd__diode_2 ANTENNA__13593__B2 (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA__13594__A (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA__13594__B (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA__13594__C (.DIODE(net499));
 sky130_fd_sc_hd__diode_2 ANTENNA__13594__D (.DIODE(net495));
 sky130_fd_sc_hd__diode_2 ANTENNA__13595__A1_N (.DIODE(net504));
 sky130_fd_sc_hd__diode_2 ANTENNA__13595__A2_N (.DIODE(net403));
 sky130_fd_sc_hd__diode_2 ANTENNA__13596__C (.DIODE(net504));
 sky130_fd_sc_hd__diode_2 ANTENNA__13596__D (.DIODE(net403));
 sky130_fd_sc_hd__diode_2 ANTENNA__13609__A1 (.DIODE(net428));
 sky130_fd_sc_hd__diode_2 ANTENNA__13609__A2 (.DIODE(net483));
 sky130_fd_sc_hd__diode_2 ANTENNA__13610__A1 (.DIODE(net419));
 sky130_fd_sc_hd__diode_2 ANTENNA__13610__A2 (.DIODE(net487));
 sky130_fd_sc_hd__diode_2 ANTENNA__13610__B1 (.DIODE(net483));
 sky130_fd_sc_hd__diode_2 ANTENNA__13610__B2 (.DIODE(net423));
 sky130_fd_sc_hd__diode_2 ANTENNA__13611__A (.DIODE(net423));
 sky130_fd_sc_hd__diode_2 ANTENNA__13611__B (.DIODE(net419));
 sky130_fd_sc_hd__diode_2 ANTENNA__13611__C (.DIODE(net487));
 sky130_fd_sc_hd__diode_2 ANTENNA__13611__D (.DIODE(net483));
 sky130_fd_sc_hd__diode_2 ANTENNA__13612__A1 (.DIODE(net416));
 sky130_fd_sc_hd__diode_2 ANTENNA__13612__A2 (.DIODE(net491));
 sky130_fd_sc_hd__diode_2 ANTENNA__13613__A (.DIODE(net416));
 sky130_fd_sc_hd__diode_2 ANTENNA__13613__B (.DIODE(net491));
 sky130_fd_sc_hd__diode_2 ANTENNA__13619__A (.DIODE(net428));
 sky130_fd_sc_hd__diode_2 ANTENNA__13619__B (.DIODE(net478));
 sky130_fd_sc_hd__diode_2 ANTENNA__13620__A (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA__13620__B (.DIODE(net433));
 sky130_fd_sc_hd__diode_2 ANTENNA__13620__C (.DIODE(net474));
 sky130_fd_sc_hd__diode_2 ANTENNA__13620__D (.DIODE(net470));
 sky130_fd_sc_hd__diode_2 ANTENNA__13621__A1 (.DIODE(net433));
 sky130_fd_sc_hd__diode_2 ANTENNA__13621__A2 (.DIODE(net474));
 sky130_fd_sc_hd__diode_2 ANTENNA__13621__B1 (.DIODE(net470));
 sky130_fd_sc_hd__diode_2 ANTENNA__13621__B2 (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA__13624__A (.DIODE(net442));
 sky130_fd_sc_hd__diode_2 ANTENNA__13624__B (.DIODE(net466));
 sky130_fd_sc_hd__diode_2 ANTENNA__13625__A (.DIODE(net451));
 sky130_fd_sc_hd__diode_2 ANTENNA__13625__B (.DIODE(net447));
 sky130_fd_sc_hd__diode_2 ANTENNA__13625__C (.DIODE(net463));
 sky130_fd_sc_hd__diode_2 ANTENNA__13625__D (.DIODE(net460));
 sky130_fd_sc_hd__diode_2 ANTENNA__13626__A1 (.DIODE(net447));
 sky130_fd_sc_hd__diode_2 ANTENNA__13626__A2 (.DIODE(net463));
 sky130_fd_sc_hd__diode_2 ANTENNA__13626__B1 (.DIODE(net460));
 sky130_fd_sc_hd__diode_2 ANTENNA__13626__B2 (.DIODE(net451));
 sky130_fd_sc_hd__diode_2 ANTENNA__13665__A (.DIODE(_03057_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13665__B (.DIODE(_05156_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13666__A1 (.DIODE(net600));
 sky130_fd_sc_hd__diode_2 ANTENNA__13666__B1 (.DIODE(_02619_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13666__B2 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__13670__A1 (.DIODE(net574));
 sky130_fd_sc_hd__diode_2 ANTENNA__13670__A2 (.DIODE(net336));
 sky130_fd_sc_hd__diode_2 ANTENNA__13670__B1 (.DIODE(net333));
 sky130_fd_sc_hd__diode_2 ANTENNA__13670__B2 (.DIODE(net578));
 sky130_fd_sc_hd__diode_2 ANTENNA__13671__A (.DIODE(net574));
 sky130_fd_sc_hd__diode_2 ANTENNA__13671__B (.DIODE(net578));
 sky130_fd_sc_hd__diode_2 ANTENNA__13671__C (.DIODE(net333));
 sky130_fd_sc_hd__diode_2 ANTENNA__13672__A1 (.DIODE(net336));
 sky130_fd_sc_hd__diode_2 ANTENNA__13673__A (.DIODE(net584));
 sky130_fd_sc_hd__diode_2 ANTENNA__13673__B (.DIODE(net330));
 sky130_fd_sc_hd__diode_2 ANTENNA__13679__A1 (.DIODE(net559));
 sky130_fd_sc_hd__diode_2 ANTENNA__13679__A2 (.DIODE(net344));
 sky130_fd_sc_hd__diode_2 ANTENNA__13680__A (.DIODE(net559));
 sky130_fd_sc_hd__diode_2 ANTENNA__13680__C (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA__13680__D (.DIODE(net341));
 sky130_fd_sc_hd__diode_2 ANTENNA__13681__A1_N (.DIODE(net568));
 sky130_fd_sc_hd__diode_2 ANTENNA__13681__A2_N (.DIODE(net337));
 sky130_fd_sc_hd__diode_2 ANTENNA__13682__C (.DIODE(net568));
 sky130_fd_sc_hd__diode_2 ANTENNA__13682__D (.DIODE(net337));
 sky130_fd_sc_hd__diode_2 ANTENNA__13704__A1 (.DIODE(net546));
 sky130_fd_sc_hd__diode_2 ANTENNA__13704__A2 (.DIODE(net356));
 sky130_fd_sc_hd__diode_2 ANTENNA__13704__B1 (.DIODE(net355));
 sky130_fd_sc_hd__diode_2 ANTENNA__13704__B2 (.DIODE(net551));
 sky130_fd_sc_hd__diode_2 ANTENNA__13705__A (.DIODE(net546));
 sky130_fd_sc_hd__diode_2 ANTENNA__13705__B (.DIODE(net550));
 sky130_fd_sc_hd__diode_2 ANTENNA__13705__C (.DIODE(net356));
 sky130_fd_sc_hd__diode_2 ANTENNA__13705__D (.DIODE(net354));
 sky130_fd_sc_hd__diode_2 ANTENNA__13706__A1 (.DIODE(net555));
 sky130_fd_sc_hd__diode_2 ANTENNA__13706__A2 (.DIODE(net348));
 sky130_fd_sc_hd__diode_2 ANTENNA__13707__A (.DIODE(net555));
 sky130_fd_sc_hd__diode_2 ANTENNA__13707__B (.DIODE(net348));
 sky130_fd_sc_hd__diode_2 ANTENNA__13709__A1 (.DIODE(net532));
 sky130_fd_sc_hd__diode_2 ANTENNA__13709__A2 (.DIODE(net632));
 sky130_fd_sc_hd__diode_2 ANTENNA__13709__B1 (.DIODE(net367));
 sky130_fd_sc_hd__diode_2 ANTENNA__13709__B2 (.DIODE(net537));
 sky130_fd_sc_hd__diode_2 ANTENNA__13710__A (.DIODE(net532));
 sky130_fd_sc_hd__diode_2 ANTENNA__13710__B (.DIODE(net537));
 sky130_fd_sc_hd__diode_2 ANTENNA__13710__C (.DIODE(net632));
 sky130_fd_sc_hd__diode_2 ANTENNA__13710__D (.DIODE(net367));
 sky130_fd_sc_hd__diode_2 ANTENNA__13711__A1_N (.DIODE(net542));
 sky130_fd_sc_hd__diode_2 ANTENNA__13711__A2_N (.DIODE(net363));
 sky130_fd_sc_hd__diode_2 ANTENNA__13712__C (.DIODE(net542));
 sky130_fd_sc_hd__diode_2 ANTENNA__13712__D (.DIODE(net363));
 sky130_fd_sc_hd__diode_2 ANTENNA__13721__A1 (.DIODE(net517));
 sky130_fd_sc_hd__diode_2 ANTENNA__13721__A2 (.DIODE(net383));
 sky130_fd_sc_hd__diode_2 ANTENNA__13721__B1 (.DIODE(net377));
 sky130_fd_sc_hd__diode_2 ANTENNA__13721__B2 (.DIODE(net524));
 sky130_fd_sc_hd__diode_2 ANTENNA__13722__A (.DIODE(net517));
 sky130_fd_sc_hd__diode_2 ANTENNA__13722__B (.DIODE(net524));
 sky130_fd_sc_hd__diode_2 ANTENNA__13722__C (.DIODE(net383));
 sky130_fd_sc_hd__diode_2 ANTENNA__13722__D (.DIODE(net377));
 sky130_fd_sc_hd__diode_2 ANTENNA__13723__A1 (.DIODE(net527));
 sky130_fd_sc_hd__diode_2 ANTENNA__13723__A2 (.DIODE(net374));
 sky130_fd_sc_hd__diode_2 ANTENNA__13724__A (.DIODE(net527));
 sky130_fd_sc_hd__diode_2 ANTENNA__13724__B (.DIODE(net374));
 sky130_fd_sc_hd__diode_2 ANTENNA__13741__A1 (.DIODE(net504));
 sky130_fd_sc_hd__diode_2 ANTENNA__13741__A2 (.DIODE(net397));
 sky130_fd_sc_hd__diode_2 ANTENNA__13741__B1 (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA__13741__B2 (.DIODE(net508));
 sky130_fd_sc_hd__diode_2 ANTENNA__13742__A (.DIODE(net504));
 sky130_fd_sc_hd__diode_2 ANTENNA__13742__B (.DIODE(net508));
 sky130_fd_sc_hd__diode_2 ANTENNA__13742__C (.DIODE(net397));
 sky130_fd_sc_hd__diode_2 ANTENNA__13742__D (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA__13745__A (.DIODE(net512));
 sky130_fd_sc_hd__diode_2 ANTENNA__13745__B (.DIODE(net387));
 sky130_fd_sc_hd__diode_2 ANTENNA__13747__A1 (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA__13747__A2 (.DIODE(net495));
 sky130_fd_sc_hd__diode_2 ANTENNA__13747__B1 (.DIODE(net491));
 sky130_fd_sc_hd__diode_2 ANTENNA__13747__B2 (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA__13748__A (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA__13748__B (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA__13748__C (.DIODE(net495));
 sky130_fd_sc_hd__diode_2 ANTENNA__13748__D (.DIODE(net491));
 sky130_fd_sc_hd__diode_2 ANTENNA__13749__A1 (.DIODE(net403));
 sky130_fd_sc_hd__diode_2 ANTENNA__13749__A2 (.DIODE(net499));
 sky130_fd_sc_hd__diode_2 ANTENNA__13750__A (.DIODE(net403));
 sky130_fd_sc_hd__diode_2 ANTENNA__13750__B (.DIODE(net499));
 sky130_fd_sc_hd__diode_2 ANTENNA__13761__A1 (.DIODE(net423));
 sky130_fd_sc_hd__diode_2 ANTENNA__13761__A2 (.DIODE(net419));
 sky130_fd_sc_hd__diode_2 ANTENNA__13761__A3 (.DIODE(net487));
 sky130_fd_sc_hd__diode_2 ANTENNA__13761__A4 (.DIODE(net482));
 sky130_fd_sc_hd__diode_2 ANTENNA__13762__A1 (.DIODE(net428));
 sky130_fd_sc_hd__diode_2 ANTENNA__13762__A2 (.DIODE(net478));
 sky130_fd_sc_hd__diode_2 ANTENNA__13763__A1 (.DIODE(net419));
 sky130_fd_sc_hd__diode_2 ANTENNA__13763__A2 (.DIODE(net483));
 sky130_fd_sc_hd__diode_2 ANTENNA__13763__B1 (.DIODE(net478));
 sky130_fd_sc_hd__diode_2 ANTENNA__13763__B2 (.DIODE(net423));
 sky130_fd_sc_hd__diode_2 ANTENNA__13764__A (.DIODE(net423));
 sky130_fd_sc_hd__diode_2 ANTENNA__13764__B (.DIODE(net419));
 sky130_fd_sc_hd__diode_2 ANTENNA__13764__C (.DIODE(net483));
 sky130_fd_sc_hd__diode_2 ANTENNA__13764__D (.DIODE(net478));
 sky130_fd_sc_hd__diode_2 ANTENNA__13765__A1 (.DIODE(net415));
 sky130_fd_sc_hd__diode_2 ANTENNA__13765__A2 (.DIODE(net487));
 sky130_fd_sc_hd__diode_2 ANTENNA__13766__A (.DIODE(net415));
 sky130_fd_sc_hd__diode_2 ANTENNA__13766__B (.DIODE(net487));
 sky130_fd_sc_hd__diode_2 ANTENNA__13771__A (.DIODE(net428));
 sky130_fd_sc_hd__diode_2 ANTENNA__13771__B (.DIODE(net474));
 sky130_fd_sc_hd__diode_2 ANTENNA__13772__A1 (.DIODE(net433));
 sky130_fd_sc_hd__diode_2 ANTENNA__13772__A2 (.DIODE(net470));
 sky130_fd_sc_hd__diode_2 ANTENNA__13772__B1 (.DIODE(net466));
 sky130_fd_sc_hd__diode_2 ANTENNA__13772__B2 (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA__13773__A (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA__13773__B (.DIODE(net433));
 sky130_fd_sc_hd__diode_2 ANTENNA__13773__C (.DIODE(net470));
 sky130_fd_sc_hd__diode_2 ANTENNA__13774__A1 (.DIODE(net466));
 sky130_fd_sc_hd__diode_2 ANTENNA__13776__A (.DIODE(net442));
 sky130_fd_sc_hd__diode_2 ANTENNA__13776__B (.DIODE(net463));
 sky130_fd_sc_hd__diode_2 ANTENNA__13777__A1 (.DIODE(net447));
 sky130_fd_sc_hd__diode_2 ANTENNA__13777__A2 (.DIODE(net460));
 sky130_fd_sc_hd__diode_2 ANTENNA__13777__B1 (.DIODE(net459));
 sky130_fd_sc_hd__diode_2 ANTENNA__13777__B2 (.DIODE(net451));
 sky130_fd_sc_hd__diode_2 ANTENNA__13778__A (.DIODE(net451));
 sky130_fd_sc_hd__diode_2 ANTENNA__13778__B (.DIODE(net447));
 sky130_fd_sc_hd__diode_2 ANTENNA__13778__C (.DIODE(net460));
 sky130_fd_sc_hd__diode_2 ANTENNA__13778__D (.DIODE(net459));
 sky130_fd_sc_hd__diode_2 ANTENNA__13815__A (.DIODE(_03057_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13815__B (.DIODE(_05305_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13816__A1 (.DIODE(net600));
 sky130_fd_sc_hd__diode_2 ANTENNA__13816__B1 (.DIODE(_02626_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13816__B2 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__13820__A1 (.DIODE(net569));
 sky130_fd_sc_hd__diode_2 ANTENNA__13820__A2 (.DIODE(net336));
 sky130_fd_sc_hd__diode_2 ANTENNA__13820__B1 (.DIODE(net333));
 sky130_fd_sc_hd__diode_2 ANTENNA__13820__B2 (.DIODE(net574));
 sky130_fd_sc_hd__diode_2 ANTENNA__13822__A (.DIODE(net569));
 sky130_fd_sc_hd__diode_2 ANTENNA__13822__C (.DIODE(net336));
 sky130_fd_sc_hd__diode_2 ANTENNA__13822__D (.DIODE(net333));
 sky130_fd_sc_hd__diode_2 ANTENNA__13823__A1_N (.DIODE(net578));
 sky130_fd_sc_hd__diode_2 ANTENNA__13823__A2_N (.DIODE(net330));
 sky130_fd_sc_hd__diode_2 ANTENNA__13824__B (.DIODE(net330));
 sky130_fd_sc_hd__diode_2 ANTENNA__13824__C (.DIODE(net578));
 sky130_fd_sc_hd__diode_2 ANTENNA__13826__A1 (.DIODE(net584));
 sky130_fd_sc_hd__diode_2 ANTENNA__13826__A2 (.DIODE(net330));
 sky130_fd_sc_hd__diode_2 ANTENNA__13826__B2 (.DIODE(net336));
 sky130_fd_sc_hd__diode_2 ANTENNA__13829__A (.DIODE(net584));
 sky130_fd_sc_hd__diode_2 ANTENNA__13829__B (.DIODE(net328));
 sky130_fd_sc_hd__diode_2 ANTENNA__13836__A1 (.DIODE(net555));
 sky130_fd_sc_hd__diode_2 ANTENNA__13836__A2 (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA__13836__B2 (.DIODE(net559));
 sky130_fd_sc_hd__diode_2 ANTENNA__13837__A (.DIODE(net555));
 sky130_fd_sc_hd__diode_2 ANTENNA__13837__B (.DIODE(net559));
 sky130_fd_sc_hd__diode_2 ANTENNA__13837__C (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA__13838__A2 (.DIODE(net337));
 sky130_fd_sc_hd__diode_2 ANTENNA__13839__B (.DIODE(net337));
 sky130_fd_sc_hd__diode_2 ANTENNA__13857__A1 (.DIODE(net542));
 sky130_fd_sc_hd__diode_2 ANTENNA__13857__A2 (.DIODE(net356));
 sky130_fd_sc_hd__diode_2 ANTENNA__13857__B1 (.DIODE(net354));
 sky130_fd_sc_hd__diode_2 ANTENNA__13857__B2 (.DIODE(net546));
 sky130_fd_sc_hd__diode_2 ANTENNA__13858__A (.DIODE(net542));
 sky130_fd_sc_hd__diode_2 ANTENNA__13858__B (.DIODE(net546));
 sky130_fd_sc_hd__diode_2 ANTENNA__13858__C (.DIODE(net356));
 sky130_fd_sc_hd__diode_2 ANTENNA__13858__D (.DIODE(net354));
 sky130_fd_sc_hd__diode_2 ANTENNA__13860__A (.DIODE(net550));
 sky130_fd_sc_hd__diode_2 ANTENNA__13860__B (.DIODE(net348));
 sky130_fd_sc_hd__diode_2 ANTENNA__13862__A1 (.DIODE(net527));
 sky130_fd_sc_hd__diode_2 ANTENNA__13862__A2 (.DIODE(net632));
 sky130_fd_sc_hd__diode_2 ANTENNA__13862__B1 (.DIODE(net367));
 sky130_fd_sc_hd__diode_2 ANTENNA__13862__B2 (.DIODE(net532));
 sky130_fd_sc_hd__diode_2 ANTENNA__13863__A (.DIODE(net527));
 sky130_fd_sc_hd__diode_2 ANTENNA__13863__B (.DIODE(net532));
 sky130_fd_sc_hd__diode_2 ANTENNA__13863__C (.DIODE(net632));
 sky130_fd_sc_hd__diode_2 ANTENNA__13863__D (.DIODE(net367));
 sky130_fd_sc_hd__diode_2 ANTENNA__13864__A (.DIODE(\mul0.a[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13864__B (.DIODE(net532));
 sky130_fd_sc_hd__diode_2 ANTENNA__13864__C (.DIODE(net632));
 sky130_fd_sc_hd__diode_2 ANTENNA__13864__D (.DIODE(net367));
 sky130_fd_sc_hd__diode_2 ANTENNA__13865__A1 (.DIODE(net537));
 sky130_fd_sc_hd__diode_2 ANTENNA__13865__A2 (.DIODE(net363));
 sky130_fd_sc_hd__diode_2 ANTENNA__13866__A (.DIODE(net537));
 sky130_fd_sc_hd__diode_2 ANTENNA__13866__B (.DIODE(net363));
 sky130_fd_sc_hd__diode_2 ANTENNA__13867__A (.DIODE(net537));
 sky130_fd_sc_hd__diode_2 ANTENNA__13867__B (.DIODE(net363));
 sky130_fd_sc_hd__diode_2 ANTENNA__13872__A1 (.DIODE(net517));
 sky130_fd_sc_hd__diode_2 ANTENNA__13872__A2 (.DIODE(net521));
 sky130_fd_sc_hd__diode_2 ANTENNA__13872__A3 (.DIODE(net383));
 sky130_fd_sc_hd__diode_2 ANTENNA__13872__A4 (.DIODE(net377));
 sky130_fd_sc_hd__diode_2 ANTENNA__13873__A1 (.DIODE(net512));
 sky130_fd_sc_hd__diode_2 ANTENNA__13873__A2 (.DIODE(net387));
 sky130_fd_sc_hd__diode_2 ANTENNA__13874__A1 (.DIODE(\mul0.a[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13874__A2 (.DIODE(net383));
 sky130_fd_sc_hd__diode_2 ANTENNA__13874__B1 (.DIODE(net377));
 sky130_fd_sc_hd__diode_2 ANTENNA__13874__B2 (.DIODE(net517));
 sky130_fd_sc_hd__diode_2 ANTENNA__13875__A (.DIODE(\mul0.a[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13875__B (.DIODE(net517));
 sky130_fd_sc_hd__diode_2 ANTENNA__13875__C (.DIODE(net383));
 sky130_fd_sc_hd__diode_2 ANTENNA__13875__D (.DIODE(net377));
 sky130_fd_sc_hd__diode_2 ANTENNA__13876__A1 (.DIODE(net524));
 sky130_fd_sc_hd__diode_2 ANTENNA__13876__A2 (.DIODE(net374));
 sky130_fd_sc_hd__diode_2 ANTENNA__13877__A (.DIODE(net524));
 sky130_fd_sc_hd__diode_2 ANTENNA__13877__B (.DIODE(net374));
 sky130_fd_sc_hd__diode_2 ANTENNA__13892__A1 (.DIODE(net504));
 sky130_fd_sc_hd__diode_2 ANTENNA__13892__A2 (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA__13892__B1 (.DIODE(net499));
 sky130_fd_sc_hd__diode_2 ANTENNA__13892__B2 (.DIODE(net397));
 sky130_fd_sc_hd__diode_2 ANTENNA__13893__A (.DIODE(net504));
 sky130_fd_sc_hd__diode_2 ANTENNA__13893__B (.DIODE(net397));
 sky130_fd_sc_hd__diode_2 ANTENNA__13893__C (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA__13894__A1 (.DIODE(net499));
 sky130_fd_sc_hd__diode_2 ANTENNA__13895__A (.DIODE(net508));
 sky130_fd_sc_hd__diode_2 ANTENNA__13895__B (.DIODE(net387));
 sky130_fd_sc_hd__diode_2 ANTENNA__13897__A1 (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA__13897__A2 (.DIODE(net491));
 sky130_fd_sc_hd__diode_2 ANTENNA__13897__B1 (.DIODE(net487));
 sky130_fd_sc_hd__diode_2 ANTENNA__13897__B2 (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA__13898__A (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA__13898__B (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA__13898__C (.DIODE(net491));
 sky130_fd_sc_hd__diode_2 ANTENNA__13898__D (.DIODE(net487));
 sky130_fd_sc_hd__diode_2 ANTENNA__13899__A (.DIODE(net403));
 sky130_fd_sc_hd__diode_2 ANTENNA__13899__B (.DIODE(net495));
 sky130_fd_sc_hd__diode_2 ANTENNA__13911__A1 (.DIODE(net428));
 sky130_fd_sc_hd__diode_2 ANTENNA__13911__A2 (.DIODE(net474));
 sky130_fd_sc_hd__diode_2 ANTENNA__13911__B2 (.DIODE(net466));
 sky130_fd_sc_hd__diode_2 ANTENNA__13912__A1 (.DIODE(net419));
 sky130_fd_sc_hd__diode_2 ANTENNA__13912__A2 (.DIODE(net478));
 sky130_fd_sc_hd__diode_2 ANTENNA__13912__B1 (.DIODE(net474));
 sky130_fd_sc_hd__diode_2 ANTENNA__13912__B2 (.DIODE(net423));
 sky130_fd_sc_hd__diode_2 ANTENNA__13913__A (.DIODE(net423));
 sky130_fd_sc_hd__diode_2 ANTENNA__13913__B (.DIODE(net419));
 sky130_fd_sc_hd__diode_2 ANTENNA__13913__C (.DIODE(net478));
 sky130_fd_sc_hd__diode_2 ANTENNA__13913__D (.DIODE(net474));
 sky130_fd_sc_hd__diode_2 ANTENNA__13914__A1 (.DIODE(net415));
 sky130_fd_sc_hd__diode_2 ANTENNA__13914__A2 (.DIODE(net482));
 sky130_fd_sc_hd__diode_2 ANTENNA__13915__A (.DIODE(net415));
 sky130_fd_sc_hd__diode_2 ANTENNA__13915__B (.DIODE(net482));
 sky130_fd_sc_hd__diode_2 ANTENNA__13920__A1 (.DIODE(net433));
 sky130_fd_sc_hd__diode_2 ANTENNA__13920__A2 (.DIODE(net466));
 sky130_fd_sc_hd__diode_2 ANTENNA__13920__B1 (.DIODE(net463));
 sky130_fd_sc_hd__diode_2 ANTENNA__13920__B2 (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA__13921__A (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA__13921__B (.DIODE(net433));
 sky130_fd_sc_hd__diode_2 ANTENNA__13921__C (.DIODE(net466));
 sky130_fd_sc_hd__diode_2 ANTENNA__13921__D (.DIODE(net463));
 sky130_fd_sc_hd__diode_2 ANTENNA__13922__C (.DIODE(net428));
 sky130_fd_sc_hd__diode_2 ANTENNA__13922__D (.DIODE(net470));
 sky130_fd_sc_hd__diode_2 ANTENNA__13923__A1_N (.DIODE(net428));
 sky130_fd_sc_hd__diode_2 ANTENNA__13923__A2_N (.DIODE(net470));
 sky130_fd_sc_hd__diode_2 ANTENNA__13925__A (.DIODE(net442));
 sky130_fd_sc_hd__diode_2 ANTENNA__13925__B (.DIODE(net460));
 sky130_fd_sc_hd__diode_2 ANTENNA__13926__A1 (.DIODE(net447));
 sky130_fd_sc_hd__diode_2 ANTENNA__13926__A2 (.DIODE(net459));
 sky130_fd_sc_hd__diode_2 ANTENNA__13926__B2 (.DIODE(net452));
 sky130_fd_sc_hd__diode_2 ANTENNA__13927__A (.DIODE(net452));
 sky130_fd_sc_hd__diode_2 ANTENNA__13927__B (.DIODE(\mul0.b[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13927__C (.DIODE(net459));
 sky130_fd_sc_hd__diode_2 ANTENNA__13968__A1 (.DIODE(net600));
 sky130_fd_sc_hd__diode_2 ANTENNA__13968__B1 (.DIODE(_02632_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13968__B2 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__13969__A1 (.DIODE(_03058_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13969__A2 (.DIODE(_05457_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13970__S (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__13974__A1 (.DIODE(net559));
 sky130_fd_sc_hd__diode_2 ANTENNA__13974__A2 (.DIODE(net337));
 sky130_fd_sc_hd__diode_2 ANTENNA__13974__B1 (.DIODE(net336));
 sky130_fd_sc_hd__diode_2 ANTENNA__13975__A (.DIODE(net559));
 sky130_fd_sc_hd__diode_2 ANTENNA__13975__C (.DIODE(net337));
 sky130_fd_sc_hd__diode_2 ANTENNA__13975__D (.DIODE(net336));
 sky130_fd_sc_hd__diode_2 ANTENNA__13976__A1_N (.DIODE(net568));
 sky130_fd_sc_hd__diode_2 ANTENNA__13976__A2_N (.DIODE(net333));
 sky130_fd_sc_hd__diode_2 ANTENNA__13977__C (.DIODE(net569));
 sky130_fd_sc_hd__diode_2 ANTENNA__13977__D (.DIODE(net333));
 sky130_fd_sc_hd__diode_2 ANTENNA__13982__A1 (.DIODE(net574));
 sky130_fd_sc_hd__diode_2 ANTENNA__13982__A2 (.DIODE(net330));
 sky130_fd_sc_hd__diode_2 ANTENNA__13982__B1 (.DIODE(net328));
 sky130_fd_sc_hd__diode_2 ANTENNA__13982__B2 (.DIODE(net578));
 sky130_fd_sc_hd__diode_2 ANTENNA__13983__A (.DIODE(net574));
 sky130_fd_sc_hd__diode_2 ANTENNA__13983__B (.DIODE(net578));
 sky130_fd_sc_hd__diode_2 ANTENNA__13983__C (.DIODE(net330));
 sky130_fd_sc_hd__diode_2 ANTENNA__13983__D (.DIODE(net328));
 sky130_fd_sc_hd__diode_2 ANTENNA__13984__A1 (.DIODE(net584));
 sky130_fd_sc_hd__diode_2 ANTENNA__13984__A2 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__13985__A (.DIODE(net584));
 sky130_fd_sc_hd__diode_2 ANTENNA__13985__B (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__13994__A1 (.DIODE(net555));
 sky130_fd_sc_hd__diode_2 ANTENNA__13994__A2 (.DIODE(net559));
 sky130_fd_sc_hd__diode_2 ANTENNA__13994__A3 (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA__13994__A4 (.DIODE(net341));
 sky130_fd_sc_hd__diode_2 ANTENNA__13996__A1 (.DIODE(net546));
 sky130_fd_sc_hd__diode_2 ANTENNA__13996__A2 (.DIODE(net348));
 sky130_fd_sc_hd__diode_2 ANTENNA__13996__B1 (.DIODE(net344));
 sky130_fd_sc_hd__diode_2 ANTENNA__13996__B2 (.DIODE(net551));
 sky130_fd_sc_hd__diode_2 ANTENNA__13997__A (.DIODE(net547));
 sky130_fd_sc_hd__diode_2 ANTENNA__13997__B (.DIODE(net551));
 sky130_fd_sc_hd__diode_2 ANTENNA__13997__C (.DIODE(net348));
 sky130_fd_sc_hd__diode_2 ANTENNA__13997__D (.DIODE(net344));
 sky130_fd_sc_hd__diode_2 ANTENNA__13998__A1 (.DIODE(net555));
 sky130_fd_sc_hd__diode_2 ANTENNA__13999__A (.DIODE(net555));
 sky130_fd_sc_hd__diode_2 ANTENNA__14017__A1 (.DIODE(net533));
 sky130_fd_sc_hd__diode_2 ANTENNA__14017__A2 (.DIODE(net364));
 sky130_fd_sc_hd__diode_2 ANTENNA__14017__B1 (.DIODE(net356));
 sky130_fd_sc_hd__diode_2 ANTENNA__14017__B2 (.DIODE(net538));
 sky130_fd_sc_hd__diode_2 ANTENNA__14018__A (.DIODE(net533));
 sky130_fd_sc_hd__diode_2 ANTENNA__14018__B (.DIODE(net538));
 sky130_fd_sc_hd__diode_2 ANTENNA__14018__C (.DIODE(net364));
 sky130_fd_sc_hd__diode_2 ANTENNA__14018__D (.DIODE(net360));
 sky130_fd_sc_hd__diode_2 ANTENNA__14019__A1 (.DIODE(net543));
 sky130_fd_sc_hd__diode_2 ANTENNA__14019__A2 (.DIODE(net354));
 sky130_fd_sc_hd__diode_2 ANTENNA__14020__A (.DIODE(net543));
 sky130_fd_sc_hd__diode_2 ANTENNA__14020__B (.DIODE(net352));
 sky130_fd_sc_hd__diode_2 ANTENNA__14022__A1 (.DIODE(net519));
 sky130_fd_sc_hd__diode_2 ANTENNA__14022__A2 (.DIODE(net372));
 sky130_fd_sc_hd__diode_2 ANTENNA__14022__B1 (.DIODE(net632));
 sky130_fd_sc_hd__diode_2 ANTENNA__14022__B2 (.DIODE(net521));
 sky130_fd_sc_hd__diode_2 ANTENNA__14023__A (.DIODE(net519));
 sky130_fd_sc_hd__diode_2 ANTENNA__14023__B (.DIODE(net523));
 sky130_fd_sc_hd__diode_2 ANTENNA__14023__C (.DIODE(net372));
 sky130_fd_sc_hd__diode_2 ANTENNA__14024__A (.DIODE(net519));
 sky130_fd_sc_hd__diode_2 ANTENNA__14024__B (.DIODE(net521));
 sky130_fd_sc_hd__diode_2 ANTENNA__14024__C (.DIODE(net372));
 sky130_fd_sc_hd__diode_2 ANTENNA__14024__D (.DIODE(net632));
 sky130_fd_sc_hd__diode_2 ANTENNA__14025__A1 (.DIODE(net529));
 sky130_fd_sc_hd__diode_2 ANTENNA__14026__A (.DIODE(net527));
 sky130_fd_sc_hd__diode_2 ANTENNA__14026__B (.DIODE(net367));
 sky130_fd_sc_hd__diode_2 ANTENNA__14027__A (.DIODE(net527));
 sky130_fd_sc_hd__diode_2 ANTENNA__14033__A1 (.DIODE(\mul0.a[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14033__A2 (.DIODE(net387));
 sky130_fd_sc_hd__diode_2 ANTENNA__14033__B2 (.DIODE(net499));
 sky130_fd_sc_hd__diode_2 ANTENNA__14034__A1 (.DIODE(net504));
 sky130_fd_sc_hd__diode_2 ANTENNA__14034__A2 (.DIODE(net387));
 sky130_fd_sc_hd__diode_2 ANTENNA__14034__B1 (.DIODE(net383));
 sky130_fd_sc_hd__diode_2 ANTENNA__14034__B2 (.DIODE(\mul0.a[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14035__A (.DIODE(net504));
 sky130_fd_sc_hd__diode_2 ANTENNA__14035__B (.DIODE(\mul0.a[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14035__C (.DIODE(net387));
 sky130_fd_sc_hd__diode_2 ANTENNA__14035__D (.DIODE(net383));
 sky130_fd_sc_hd__diode_2 ANTENNA__14036__A1 (.DIODE(\mul0.a[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14036__A2 (.DIODE(net377));
 sky130_fd_sc_hd__diode_2 ANTENNA__14037__A (.DIODE(\mul0.a[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14037__B (.DIODE(net377));
 sky130_fd_sc_hd__diode_2 ANTENNA__14053__A (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA__14053__B (.DIODE(net499));
 sky130_fd_sc_hd__diode_2 ANTENNA__14054__A1 (.DIODE(net397));
 sky130_fd_sc_hd__diode_2 ANTENNA__14054__A2 (.DIODE(net495));
 sky130_fd_sc_hd__diode_2 ANTENNA__14054__B1 (.DIODE(net491));
 sky130_fd_sc_hd__diode_2 ANTENNA__14054__B2 (.DIODE(net403));
 sky130_fd_sc_hd__diode_2 ANTENNA__14055__A (.DIODE(net403));
 sky130_fd_sc_hd__diode_2 ANTENNA__14055__B (.DIODE(net397));
 sky130_fd_sc_hd__diode_2 ANTENNA__14055__C (.DIODE(net491));
 sky130_fd_sc_hd__diode_2 ANTENNA__14056__A1 (.DIODE(net495));
 sky130_fd_sc_hd__diode_2 ANTENNA__14058__A (.DIODE(net406));
 sky130_fd_sc_hd__diode_2 ANTENNA__14058__B (.DIODE(net487));
 sky130_fd_sc_hd__diode_2 ANTENNA__14059__A1 (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA__14059__A2 (.DIODE(net483));
 sky130_fd_sc_hd__diode_2 ANTENNA__14059__B1 (.DIODE(net481));
 sky130_fd_sc_hd__diode_2 ANTENNA__14059__B2 (.DIODE(net415));
 sky130_fd_sc_hd__diode_2 ANTENNA__14060__A (.DIODE(net415));
 sky130_fd_sc_hd__diode_2 ANTENNA__14060__B (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA__14060__C (.DIODE(net483));
 sky130_fd_sc_hd__diode_2 ANTENNA__14060__D (.DIODE(net481));
 sky130_fd_sc_hd__diode_2 ANTENNA__14074__A1 (.DIODE(net423));
 sky130_fd_sc_hd__diode_2 ANTENNA__14074__A2 (.DIODE(net470));
 sky130_fd_sc_hd__diode_2 ANTENNA__14074__B2 (.DIODE(net428));
 sky130_fd_sc_hd__diode_2 ANTENNA__14075__A (.DIODE(net428));
 sky130_fd_sc_hd__diode_2 ANTENNA__14075__B (.DIODE(net423));
 sky130_fd_sc_hd__diode_2 ANTENNA__14075__C (.DIODE(net470));
 sky130_fd_sc_hd__diode_2 ANTENNA__14076__A1 (.DIODE(net419));
 sky130_fd_sc_hd__diode_2 ANTENNA__14076__A2 (.DIODE(net474));
 sky130_fd_sc_hd__diode_2 ANTENNA__14077__A (.DIODE(net419));
 sky130_fd_sc_hd__diode_2 ANTENNA__14077__B (.DIODE(net474));
 sky130_fd_sc_hd__diode_2 ANTENNA__14082__A (.DIODE(net433));
 sky130_fd_sc_hd__diode_2 ANTENNA__14082__B (.DIODE(net463));
 sky130_fd_sc_hd__diode_2 ANTENNA__14083__A1 (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA__14083__A2 (.DIODE(net460));
 sky130_fd_sc_hd__diode_2 ANTENNA__14083__B1 (.DIODE(net459));
 sky130_fd_sc_hd__diode_2 ANTENNA__14083__B2 (.DIODE(net442));
 sky130_fd_sc_hd__diode_2 ANTENNA__14084__A (.DIODE(net442));
 sky130_fd_sc_hd__diode_2 ANTENNA__14084__B (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA__14084__C (.DIODE(net459));
 sky130_fd_sc_hd__diode_2 ANTENNA__14085__A1 (.DIODE(net460));
 sky130_fd_sc_hd__diode_2 ANTENNA__14087__A (.DIODE(net447));
 sky130_fd_sc_hd__diode_2 ANTENNA__14088__A1 (.DIODE(net451));
 sky130_fd_sc_hd__diode_2 ANTENNA__14088__A2 (.DIODE(\mul0.a[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14088__B1 (.DIODE(\mul0.b[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14089__A (.DIODE(net451));
 sky130_fd_sc_hd__diode_2 ANTENNA__14089__B (.DIODE(\mul0.a[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14089__C (.DIODE(\mul0.b[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14127__A1 (.DIODE(net600));
 sky130_fd_sc_hd__diode_2 ANTENNA__14127__B1 (.DIODE(_02638_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14127__B2 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__14128__A1 (.DIODE(_03058_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14128__A2 (.DIODE(_05615_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14133__B (.DIODE(net328));
 sky130_fd_sc_hd__diode_2 ANTENNA__14133__C (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA__14133__D (.DIODE(net574));
 sky130_fd_sc_hd__diode_2 ANTENNA__14134__A1_N (.DIODE(net574));
 sky130_fd_sc_hd__diode_2 ANTENNA__14134__A2_N (.DIODE(net328));
 sky130_fd_sc_hd__diode_2 ANTENNA__14134__B1 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__14134__B2 (.DIODE(net578));
 sky130_fd_sc_hd__diode_2 ANTENNA__14137__A1 (.DIODE(net559));
 sky130_fd_sc_hd__diode_2 ANTENNA__14137__A2 (.DIODE(net335));
 sky130_fd_sc_hd__diode_2 ANTENNA__14137__B1 (.DIODE(net332));
 sky130_fd_sc_hd__diode_2 ANTENNA__14137__B2 (.DIODE(net563));
 sky130_fd_sc_hd__diode_2 ANTENNA__14138__A (.DIODE(net559));
 sky130_fd_sc_hd__diode_2 ANTENNA__14138__B (.DIODE(net563));
 sky130_fd_sc_hd__diode_2 ANTENNA__14138__C (.DIODE(net335));
 sky130_fd_sc_hd__diode_2 ANTENNA__14139__A1 (.DIODE(net332));
 sky130_fd_sc_hd__diode_2 ANTENNA__14140__A (.DIODE(net569));
 sky130_fd_sc_hd__diode_2 ANTENNA__14140__B (.DIODE(net330));
 sky130_fd_sc_hd__diode_2 ANTENNA__14154__A1 (.DIODE(net547));
 sky130_fd_sc_hd__diode_2 ANTENNA__14154__A2 (.DIODE(net344));
 sky130_fd_sc_hd__diode_2 ANTENNA__14154__B2 (.DIODE(net551));
 sky130_fd_sc_hd__diode_2 ANTENNA__14155__A (.DIODE(net547));
 sky130_fd_sc_hd__diode_2 ANTENNA__14155__B (.DIODE(net551));
 sky130_fd_sc_hd__diode_2 ANTENNA__14155__C (.DIODE(net344));
 sky130_fd_sc_hd__diode_2 ANTENNA__14156__A1 (.DIODE(net555));
 sky130_fd_sc_hd__diode_2 ANTENNA__14156__A2 (.DIODE(net337));
 sky130_fd_sc_hd__diode_2 ANTENNA__14157__A (.DIODE(net555));
 sky130_fd_sc_hd__diode_2 ANTENNA__14157__B (.DIODE(net337));
 sky130_fd_sc_hd__diode_2 ANTENNA__14175__A1 (.DIODE(net533));
 sky130_fd_sc_hd__diode_2 ANTENNA__14175__A2 (.DIODE(net360));
 sky130_fd_sc_hd__diode_2 ANTENNA__14175__B1 (.DIODE(net352));
 sky130_fd_sc_hd__diode_2 ANTENNA__14175__B2 (.DIODE(net538));
 sky130_fd_sc_hd__diode_2 ANTENNA__14176__A (.DIODE(net533));
 sky130_fd_sc_hd__diode_2 ANTENNA__14176__B (.DIODE(net538));
 sky130_fd_sc_hd__diode_2 ANTENNA__14176__C (.DIODE(net360));
 sky130_fd_sc_hd__diode_2 ANTENNA__14177__A1 (.DIODE(net352));
 sky130_fd_sc_hd__diode_2 ANTENNA__14178__A (.DIODE(net543));
 sky130_fd_sc_hd__diode_2 ANTENNA__14178__B (.DIODE(net351));
 sky130_fd_sc_hd__diode_2 ANTENNA__14180__A1 (.DIODE(net519));
 sky130_fd_sc_hd__diode_2 ANTENNA__14180__B2 (.DIODE(net523));
 sky130_fd_sc_hd__diode_2 ANTENNA__14181__A (.DIODE(net519));
 sky130_fd_sc_hd__diode_2 ANTENNA__14181__B (.DIODE(net523));
 sky130_fd_sc_hd__diode_2 ANTENNA__14181__C (.DIODE(net632));
 sky130_fd_sc_hd__diode_2 ANTENNA__14182__A (.DIODE(net519));
 sky130_fd_sc_hd__diode_2 ANTENNA__14182__B (.DIODE(net523));
 sky130_fd_sc_hd__diode_2 ANTENNA__14183__A1 (.DIODE(net529));
 sky130_fd_sc_hd__diode_2 ANTENNA__14184__A (.DIODE(net529));
 sky130_fd_sc_hd__diode_2 ANTENNA__14185__A (.DIODE(net529));
 sky130_fd_sc_hd__diode_2 ANTENNA__14191__A1 (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA__14191__A2 (.DIODE(net499));
 sky130_fd_sc_hd__diode_2 ANTENNA__14191__B2 (.DIODE(net495));
 sky130_fd_sc_hd__diode_2 ANTENNA__14192__A1 (.DIODE(\mul0.a[17] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14192__A2 (.DIODE(net383));
 sky130_fd_sc_hd__diode_2 ANTENNA__14192__B1 (.DIODE(net377));
 sky130_fd_sc_hd__diode_2 ANTENNA__14192__B2 (.DIODE(net508));
 sky130_fd_sc_hd__diode_2 ANTENNA__14193__A (.DIODE(net504));
 sky130_fd_sc_hd__diode_2 ANTENNA__14193__B (.DIODE(net508));
 sky130_fd_sc_hd__diode_2 ANTENNA__14193__C (.DIODE(net383));
 sky130_fd_sc_hd__diode_2 ANTENNA__14193__D (.DIODE(net377));
 sky130_fd_sc_hd__diode_2 ANTENNA__14194__A1 (.DIODE(net512));
 sky130_fd_sc_hd__diode_2 ANTENNA__14194__A2 (.DIODE(net374));
 sky130_fd_sc_hd__diode_2 ANTENNA__14195__A (.DIODE(net512));
 sky130_fd_sc_hd__diode_2 ANTENNA__14195__B (.DIODE(net374));
 sky130_fd_sc_hd__diode_2 ANTENNA__14203__A (.DIODE(_05677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14204__B1 (.DIODE(_05677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14211__A1 (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA__14211__A2 (.DIODE(net495));
 sky130_fd_sc_hd__diode_2 ANTENNA__14211__B1 (.DIODE(net491));
 sky130_fd_sc_hd__diode_2 ANTENNA__14211__B2 (.DIODE(net397));
 sky130_fd_sc_hd__diode_2 ANTENNA__14212__A (.DIODE(net397));
 sky130_fd_sc_hd__diode_2 ANTENNA__14212__B (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA__14212__C (.DIODE(net495));
 sky130_fd_sc_hd__diode_2 ANTENNA__14212__D (.DIODE(net491));
 sky130_fd_sc_hd__diode_2 ANTENNA__14214__A (.DIODE(net387));
 sky130_fd_sc_hd__diode_2 ANTENNA__14214__B (.DIODE(net499));
 sky130_fd_sc_hd__diode_2 ANTENNA__14216__A1 (.DIODE(net406));
 sky130_fd_sc_hd__diode_2 ANTENNA__14216__A2 (.DIODE(net483));
 sky130_fd_sc_hd__diode_2 ANTENNA__14216__B1 (.DIODE(net481));
 sky130_fd_sc_hd__diode_2 ANTENNA__14216__B2 (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA__14217__A (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA__14217__B (.DIODE(net406));
 sky130_fd_sc_hd__diode_2 ANTENNA__14217__C (.DIODE(net483));
 sky130_fd_sc_hd__diode_2 ANTENNA__14217__D (.DIODE(net481));
 sky130_fd_sc_hd__diode_2 ANTENNA__14218__A (.DIODE(net402));
 sky130_fd_sc_hd__diode_2 ANTENNA__14218__B (.DIODE(net487));
 sky130_fd_sc_hd__diode_2 ANTENNA__14232__A1 (.DIODE(net433));
 sky130_fd_sc_hd__diode_2 ANTENNA__14232__A2 (.DIODE(net463));
 sky130_fd_sc_hd__diode_2 ANTENNA__14232__B2 (.DIODE(net460));
 sky130_fd_sc_hd__diode_2 ANTENNA__14233__A1 (.DIODE(net419));
 sky130_fd_sc_hd__diode_2 ANTENNA__14233__A2 (.DIODE(net473));
 sky130_fd_sc_hd__diode_2 ANTENNA__14233__B2 (.DIODE(net423));
 sky130_fd_sc_hd__diode_2 ANTENNA__14234__A (.DIODE(net423));
 sky130_fd_sc_hd__diode_2 ANTENNA__14234__B (.DIODE(net419));
 sky130_fd_sc_hd__diode_2 ANTENNA__14234__C (.DIODE(net470));
 sky130_fd_sc_hd__diode_2 ANTENNA__14235__A1 (.DIODE(net415));
 sky130_fd_sc_hd__diode_2 ANTENNA__14235__A2 (.DIODE(net477));
 sky130_fd_sc_hd__diode_2 ANTENNA__14236__A (.DIODE(net415));
 sky130_fd_sc_hd__diode_2 ANTENNA__14236__B (.DIODE(net477));
 sky130_fd_sc_hd__diode_2 ANTENNA__14241__A1 (.DIODE(net433));
 sky130_fd_sc_hd__diode_2 ANTENNA__14241__A2 (.DIODE(net460));
 sky130_fd_sc_hd__diode_2 ANTENNA__14241__B1 (.DIODE(net459));
 sky130_fd_sc_hd__diode_2 ANTENNA__14241__B2 (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA__14242__A (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA__14242__B (.DIODE(net433));
 sky130_fd_sc_hd__diode_2 ANTENNA__14242__C (.DIODE(net459));
 sky130_fd_sc_hd__diode_2 ANTENNA__14243__A1 (.DIODE(net460));
 sky130_fd_sc_hd__diode_2 ANTENNA__14244__A (.DIODE(net428));
 sky130_fd_sc_hd__diode_2 ANTENNA__14244__B (.DIODE(net463));
 sky130_fd_sc_hd__diode_2 ANTENNA__14247__A (.DIODE(net452));
 sky130_fd_sc_hd__diode_2 ANTENNA__14247__B (.DIODE(\mul0.b[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14248__A (.DIODE(net452));
 sky130_fd_sc_hd__diode_2 ANTENNA__14248__B (.DIODE(\mul0.b[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14248__C (.DIODE(net453));
 sky130_fd_sc_hd__diode_2 ANTENNA__14249__A1 (.DIODE(net452));
 sky130_fd_sc_hd__diode_2 ANTENNA__14249__A2 (.DIODE(\mul0.b[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14249__B1_N (.DIODE(\mul0.a[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14250__A (.DIODE(net442));
 sky130_fd_sc_hd__diode_2 ANTENNA__14297__A1 (.DIODE(net599));
 sky130_fd_sc_hd__diode_2 ANTENNA__14297__B1 (.DIODE(_02644_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14297__B2 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__14298__A1 (.DIODE(_03058_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14298__A2 (.DIODE(_05784_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14305__A1 (.DIODE(net555));
 sky130_fd_sc_hd__diode_2 ANTENNA__14305__A2 (.DIODE(net335));
 sky130_fd_sc_hd__diode_2 ANTENNA__14305__B1 (.DIODE(net332));
 sky130_fd_sc_hd__diode_2 ANTENNA__14305__B2 (.DIODE(net560));
 sky130_fd_sc_hd__diode_2 ANTENNA__14306__A (.DIODE(net555));
 sky130_fd_sc_hd__diode_2 ANTENNA__14306__B (.DIODE(net560));
 sky130_fd_sc_hd__diode_2 ANTENNA__14306__C (.DIODE(net332));
 sky130_fd_sc_hd__diode_2 ANTENNA__14307__A1 (.DIODE(net335));
 sky130_fd_sc_hd__diode_2 ANTENNA__14308__A (.DIODE(net563));
 sky130_fd_sc_hd__diode_2 ANTENNA__14308__B (.DIODE(net329));
 sky130_fd_sc_hd__diode_2 ANTENNA__14310__A1_N (.DIODE(net332));
 sky130_fd_sc_hd__diode_2 ANTENNA__14312__A_N (.DIODE(net574));
 sky130_fd_sc_hd__diode_2 ANTENNA__14312__B (.DIODE(net328));
 sky130_fd_sc_hd__diode_2 ANTENNA__14312__C (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA__14312__D (.DIODE(net569));
 sky130_fd_sc_hd__diode_2 ANTENNA__14314__A1_N (.DIODE(net569));
 sky130_fd_sc_hd__diode_2 ANTENNA__14314__A2_N (.DIODE(net328));
 sky130_fd_sc_hd__diode_2 ANTENNA__14314__B1 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__14314__B2 (.DIODE(net574));
 sky130_fd_sc_hd__diode_2 ANTENNA__14323__A1 (.DIODE(net547));
 sky130_fd_sc_hd__diode_2 ANTENNA__14323__A2 (.DIODE(net551));
 sky130_fd_sc_hd__diode_2 ANTENNA__14323__A3 (.DIODE(net344));
 sky130_fd_sc_hd__diode_2 ANTENNA__14324__A1 (.DIODE(net543));
 sky130_fd_sc_hd__diode_2 ANTENNA__14324__A2 (.DIODE(net349));
 sky130_fd_sc_hd__diode_2 ANTENNA__14324__B2 (.DIODE(net352));
 sky130_fd_sc_hd__diode_2 ANTENNA__14325__A1 (.DIODE(net543));
 sky130_fd_sc_hd__diode_2 ANTENNA__14325__A2 (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA__14325__B1 (.DIODE(net341));
 sky130_fd_sc_hd__diode_2 ANTENNA__14325__B2 (.DIODE(net547));
 sky130_fd_sc_hd__diode_2 ANTENNA__14326__A (.DIODE(net543));
 sky130_fd_sc_hd__diode_2 ANTENNA__14326__B (.DIODE(net547));
 sky130_fd_sc_hd__diode_2 ANTENNA__14326__C (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA__14326__D (.DIODE(net341));
 sky130_fd_sc_hd__diode_2 ANTENNA__14327__A1 (.DIODE(net551));
 sky130_fd_sc_hd__diode_2 ANTENNA__14327__A2 (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA__14328__A (.DIODE(net551));
 sky130_fd_sc_hd__diode_2 ANTENNA__14328__B (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA__14347__A1 (.DIODE(net529));
 sky130_fd_sc_hd__diode_2 ANTENNA__14347__A2 (.DIODE(net360));
 sky130_fd_sc_hd__diode_2 ANTENNA__14347__B1 (.DIODE(net352));
 sky130_fd_sc_hd__diode_2 ANTENNA__14347__B2 (.DIODE(net533));
 sky130_fd_sc_hd__diode_2 ANTENNA__14348__A (.DIODE(net529));
 sky130_fd_sc_hd__diode_2 ANTENNA__14348__B (.DIODE(net533));
 sky130_fd_sc_hd__diode_2 ANTENNA__14348__C (.DIODE(net352));
 sky130_fd_sc_hd__diode_2 ANTENNA__14349__A1 (.DIODE(net360));
 sky130_fd_sc_hd__diode_2 ANTENNA__14350__A (.DIODE(net538));
 sky130_fd_sc_hd__diode_2 ANTENNA__14350__B (.DIODE(net349));
 sky130_fd_sc_hd__diode_2 ANTENNA__14352__A1 (.DIODE(net514));
 sky130_fd_sc_hd__diode_2 ANTENNA__14352__A2 (.DIODE(net632));
 sky130_fd_sc_hd__diode_2 ANTENNA__14352__B2 (.DIODE(net519));
 sky130_fd_sc_hd__diode_2 ANTENNA__14353__A (.DIODE(net514));
 sky130_fd_sc_hd__diode_2 ANTENNA__14353__B (.DIODE(net519));
 sky130_fd_sc_hd__diode_2 ANTENNA__14353__C (.DIODE(net632));
 sky130_fd_sc_hd__diode_2 ANTENNA__14354__A (.DIODE(net514));
 sky130_fd_sc_hd__diode_2 ANTENNA__14354__B (.DIODE(net519));
 sky130_fd_sc_hd__diode_2 ANTENNA__14354__C (.DIODE(net632));
 sky130_fd_sc_hd__diode_2 ANTENNA__14355__A1 (.DIODE(net523));
 sky130_fd_sc_hd__diode_2 ANTENNA__14356__A (.DIODE(net523));
 sky130_fd_sc_hd__diode_2 ANTENNA__14357__A (.DIODE(net523));
 sky130_fd_sc_hd__diode_2 ANTENNA__14357__B (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 ANTENNA__14364__A1 (.DIODE(net504));
 sky130_fd_sc_hd__diode_2 ANTENNA__14364__A2 (.DIODE(net377));
 sky130_fd_sc_hd__diode_2 ANTENNA__14364__B1 (.DIODE(\mul0.a[18] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14364__B2 (.DIODE(net383));
 sky130_fd_sc_hd__diode_2 ANTENNA__14365__A (.DIODE(net504));
 sky130_fd_sc_hd__diode_2 ANTENNA__14365__B (.DIODE(net383));
 sky130_fd_sc_hd__diode_2 ANTENNA__14365__C (.DIODE(net377));
 sky130_fd_sc_hd__diode_2 ANTENNA__14365__D (.DIODE(net499));
 sky130_fd_sc_hd__diode_2 ANTENNA__14366__A1 (.DIODE(net508));
 sky130_fd_sc_hd__diode_2 ANTENNA__14366__A2 (.DIODE(net374));
 sky130_fd_sc_hd__diode_2 ANTENNA__14367__A (.DIODE(net508));
 sky130_fd_sc_hd__diode_2 ANTENNA__14367__B (.DIODE(net374));
 sky130_fd_sc_hd__diode_2 ANTENNA__14383__A1 (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA__14383__A2 (.DIODE(net490));
 sky130_fd_sc_hd__diode_2 ANTENNA__14383__B1 (.DIODE(net486));
 sky130_fd_sc_hd__diode_2 ANTENNA__14383__B2 (.DIODE(net397));
 sky130_fd_sc_hd__diode_2 ANTENNA__14384__A (.DIODE(net397));
 sky130_fd_sc_hd__diode_2 ANTENNA__14384__B (.DIODE(net394));
 sky130_fd_sc_hd__diode_2 ANTENNA__14384__C (.DIODE(net490));
 sky130_fd_sc_hd__diode_2 ANTENNA__14384__D (.DIODE(net486));
 sky130_fd_sc_hd__diode_2 ANTENNA__14386__A (.DIODE(net387));
 sky130_fd_sc_hd__diode_2 ANTENNA__14386__B (.DIODE(net494));
 sky130_fd_sc_hd__diode_2 ANTENNA__14388__A1 (.DIODE(net406));
 sky130_fd_sc_hd__diode_2 ANTENNA__14388__A2 (.DIODE(net481));
 sky130_fd_sc_hd__diode_2 ANTENNA__14388__B1 (.DIODE(net477));
 sky130_fd_sc_hd__diode_2 ANTENNA__14388__B2 (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA__14389__A (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA__14389__B (.DIODE(net406));
 sky130_fd_sc_hd__diode_2 ANTENNA__14389__C (.DIODE(net479));
 sky130_fd_sc_hd__diode_2 ANTENNA__14390__A1 (.DIODE(net402));
 sky130_fd_sc_hd__diode_2 ANTENNA__14390__A2 (.DIODE(net482));
 sky130_fd_sc_hd__diode_2 ANTENNA__14391__A (.DIODE(net402));
 sky130_fd_sc_hd__diode_2 ANTENNA__14391__B (.DIODE(net482));
 sky130_fd_sc_hd__diode_2 ANTENNA__14397__A (.DIODE(_05869_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14398__A (.DIODE(_05869_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14399__B1 (.DIODE(_05869_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14404__A1 (.DIODE(net428));
 sky130_fd_sc_hd__diode_2 ANTENNA__14404__A2 (.DIODE(net463));
 sky130_fd_sc_hd__diode_2 ANTENNA__14404__B2 (.DIODE(net460));
 sky130_fd_sc_hd__diode_2 ANTENNA__14405__A1 (.DIODE(net419));
 sky130_fd_sc_hd__diode_2 ANTENNA__14405__B2 (.DIODE(net423));
 sky130_fd_sc_hd__diode_2 ANTENNA__14406__A (.DIODE(net423));
 sky130_fd_sc_hd__diode_2 ANTENNA__14406__B (.DIODE(net419));
 sky130_fd_sc_hd__diode_2 ANTENNA__14407__A1 (.DIODE(net415));
 sky130_fd_sc_hd__diode_2 ANTENNA__14407__A2 (.DIODE(net473));
 sky130_fd_sc_hd__diode_2 ANTENNA__14408__A (.DIODE(net415));
 sky130_fd_sc_hd__diode_2 ANTENNA__14408__B (.DIODE(net473));
 sky130_fd_sc_hd__diode_2 ANTENNA__14413__A1 (.DIODE(net433));
 sky130_fd_sc_hd__diode_2 ANTENNA__14413__A2 (.DIODE(net459));
 sky130_fd_sc_hd__diode_2 ANTENNA__14413__B2 (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA__14415__A (.DIODE(net428));
 sky130_fd_sc_hd__diode_2 ANTENNA__14415__B (.DIODE(net460));
 sky130_fd_sc_hd__diode_2 ANTENNA__14417__S (.DIODE(net442));
 sky130_fd_sc_hd__diode_2 ANTENNA__14449__A (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__14449__B (.DIODE(_05935_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14450__A1 (.DIODE(net599));
 sky130_fd_sc_hd__diode_2 ANTENNA__14450__B1 (.DIODE(_02648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14450__B2 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__14456__A1 (.DIODE(net551));
 sky130_fd_sc_hd__diode_2 ANTENNA__14456__A2 (.DIODE(net335));
 sky130_fd_sc_hd__diode_2 ANTENNA__14456__B1 (.DIODE(net332));
 sky130_fd_sc_hd__diode_2 ANTENNA__14456__B2 (.DIODE(net555));
 sky130_fd_sc_hd__diode_2 ANTENNA__14457__A (.DIODE(net551));
 sky130_fd_sc_hd__diode_2 ANTENNA__14457__B (.DIODE(net556));
 sky130_fd_sc_hd__diode_2 ANTENNA__14457__C (.DIODE(net332));
 sky130_fd_sc_hd__diode_2 ANTENNA__14458__A1 (.DIODE(net335));
 sky130_fd_sc_hd__diode_2 ANTENNA__14459__A (.DIODE(net560));
 sky130_fd_sc_hd__diode_2 ANTENNA__14459__B (.DIODE(net329));
 sky130_fd_sc_hd__diode_2 ANTENNA__14461__A1_N (.DIODE(net335));
 sky130_fd_sc_hd__diode_2 ANTENNA__14463__A_N (.DIODE(net569));
 sky130_fd_sc_hd__diode_2 ANTENNA__14463__B (.DIODE(net328));
 sky130_fd_sc_hd__diode_2 ANTENNA__14463__C (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA__14463__D (.DIODE(net563));
 sky130_fd_sc_hd__diode_2 ANTENNA__14465__A1_N (.DIODE(net563));
 sky130_fd_sc_hd__diode_2 ANTENNA__14465__A2_N (.DIODE(net328));
 sky130_fd_sc_hd__diode_2 ANTENNA__14465__B1 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__14465__B2 (.DIODE(net569));
 sky130_fd_sc_hd__diode_2 ANTENNA__14475__A1 (.DIODE(net538));
 sky130_fd_sc_hd__diode_2 ANTENNA__14475__A2 (.DIODE(net349));
 sky130_fd_sc_hd__diode_2 ANTENNA__14475__B2 (.DIODE(net356));
 sky130_fd_sc_hd__diode_2 ANTENNA__14476__A1 (.DIODE(net538));
 sky130_fd_sc_hd__diode_2 ANTENNA__14476__A2 (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA__14476__B1 (.DIODE(net341));
 sky130_fd_sc_hd__diode_2 ANTENNA__14476__B2 (.DIODE(net543));
 sky130_fd_sc_hd__diode_2 ANTENNA__14477__A (.DIODE(net538));
 sky130_fd_sc_hd__diode_2 ANTENNA__14477__B (.DIODE(net543));
 sky130_fd_sc_hd__diode_2 ANTENNA__14477__C (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA__14477__D (.DIODE(net341));
 sky130_fd_sc_hd__diode_2 ANTENNA__14478__A1 (.DIODE(net547));
 sky130_fd_sc_hd__diode_2 ANTENNA__14478__A2 (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA__14479__A (.DIODE(net547));
 sky130_fd_sc_hd__diode_2 ANTENNA__14479__B (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA__14493__B (.DIODE(_05941_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14494__A (.DIODE(_05941_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14498__A1 (.DIODE(net523));
 sky130_fd_sc_hd__diode_2 ANTENNA__14498__B1 (.DIODE(net352));
 sky130_fd_sc_hd__diode_2 ANTENNA__14498__B2 (.DIODE(net529));
 sky130_fd_sc_hd__diode_2 ANTENNA__14499__A (.DIODE(net523));
 sky130_fd_sc_hd__diode_2 ANTENNA__14499__B (.DIODE(net529));
 sky130_fd_sc_hd__diode_2 ANTENNA__14499__C (.DIODE(net352));
 sky130_fd_sc_hd__diode_2 ANTENNA__14500__A1 (.DIODE(net356));
 sky130_fd_sc_hd__diode_2 ANTENNA__14501__A (.DIODE(net533));
 sky130_fd_sc_hd__diode_2 ANTENNA__14501__B (.DIODE(net349));
 sky130_fd_sc_hd__diode_2 ANTENNA__14503__A1 (.DIODE(net510));
 sky130_fd_sc_hd__diode_2 ANTENNA__14503__A2 (.DIODE(net632));
 sky130_fd_sc_hd__diode_2 ANTENNA__14503__B2 (.DIODE(net514));
 sky130_fd_sc_hd__diode_2 ANTENNA__14504__B (.DIODE(net514));
 sky130_fd_sc_hd__diode_2 ANTENNA__14505__A (.DIODE(net510));
 sky130_fd_sc_hd__diode_2 ANTENNA__14505__B (.DIODE(net514));
 sky130_fd_sc_hd__diode_2 ANTENNA__14506__A1 (.DIODE(net519));
 sky130_fd_sc_hd__diode_2 ANTENNA__14507__A (.DIODE(net519));
 sky130_fd_sc_hd__diode_2 ANTENNA__14508__A (.DIODE(net519));
 sky130_fd_sc_hd__diode_2 ANTENNA__14515__A1 (.DIODE(net377));
 sky130_fd_sc_hd__diode_2 ANTENNA__14515__B1 (.DIODE(net497));
 sky130_fd_sc_hd__diode_2 ANTENNA__14515__B2 (.DIODE(net385));
 sky130_fd_sc_hd__diode_2 ANTENNA__14516__A (.DIODE(net383));
 sky130_fd_sc_hd__diode_2 ANTENNA__14516__B (.DIODE(net380));
 sky130_fd_sc_hd__diode_2 ANTENNA__14516__D (.DIODE(net497));
 sky130_fd_sc_hd__diode_2 ANTENNA__14517__A1 (.DIODE(net504));
 sky130_fd_sc_hd__diode_2 ANTENNA__14517__A2 (.DIODE(net372));
 sky130_fd_sc_hd__diode_2 ANTENNA__14518__A (.DIODE(\mul0.a[17] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14518__B (.DIODE(net372));
 sky130_fd_sc_hd__diode_2 ANTENNA__14534__A1 (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA__14534__A2 (.DIODE(net488));
 sky130_fd_sc_hd__diode_2 ANTENNA__14534__B1 (.DIODE(net484));
 sky130_fd_sc_hd__diode_2 ANTENNA__14535__B (.DIODE(net394));
 sky130_fd_sc_hd__diode_2 ANTENNA__14535__C (.DIODE(net488));
 sky130_fd_sc_hd__diode_2 ANTENNA__14536__A1 (.DIODE(net484));
 sky130_fd_sc_hd__diode_2 ANTENNA__14537__A (.DIODE(net387));
 sky130_fd_sc_hd__diode_2 ANTENNA__14537__B (.DIODE(net493));
 sky130_fd_sc_hd__diode_2 ANTENNA__14539__A1 (.DIODE(net406));
 sky130_fd_sc_hd__diode_2 ANTENNA__14539__B1 (.DIODE(net471));
 sky130_fd_sc_hd__diode_2 ANTENNA__14539__B2 (.DIODE(net412));
 sky130_fd_sc_hd__diode_2 ANTENNA__14540__A (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA__14540__B (.DIODE(net406));
 sky130_fd_sc_hd__diode_2 ANTENNA__14540__D (.DIODE(net471));
 sky130_fd_sc_hd__diode_2 ANTENNA__14542__A1 (.DIODE(net402));
 sky130_fd_sc_hd__diode_2 ANTENNA__14542__A2 (.DIODE(net479));
 sky130_fd_sc_hd__diode_2 ANTENNA__14543__A (.DIODE(net402));
 sky130_fd_sc_hd__diode_2 ANTENNA__14543__B (.DIODE(net479));
 sky130_fd_sc_hd__diode_2 ANTENNA__14548__A (.DIODE(_06019_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14550__B1 (.DIODE(_06019_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14555__A1 (.DIODE(net428));
 sky130_fd_sc_hd__diode_2 ANTENNA__14555__A2 (.DIODE(net460));
 sky130_fd_sc_hd__diode_2 ANTENNA__14556__A1 (.DIODE(net419));
 sky130_fd_sc_hd__diode_2 ANTENNA__14556__B1 (.DIODE(net460));
 sky130_fd_sc_hd__diode_2 ANTENNA__14556__B2 (.DIODE(net423));
 sky130_fd_sc_hd__diode_2 ANTENNA__14557__A (.DIODE(net423));
 sky130_fd_sc_hd__diode_2 ANTENNA__14557__B (.DIODE(net419));
 sky130_fd_sc_hd__diode_2 ANTENNA__14557__D (.DIODE(net460));
 sky130_fd_sc_hd__diode_2 ANTENNA__14558__A1 (.DIODE(net415));
 sky130_fd_sc_hd__diode_2 ANTENNA__14558__A2 (.DIODE(net466));
 sky130_fd_sc_hd__diode_2 ANTENNA__14559__A (.DIODE(net415));
 sky130_fd_sc_hd__diode_2 ANTENNA__14564__A1 (.DIODE(net433));
 sky130_fd_sc_hd__diode_2 ANTENNA__14564__A2 (.DIODE(net456));
 sky130_fd_sc_hd__diode_2 ANTENNA__14564__B1 (.DIODE(net453));
 sky130_fd_sc_hd__diode_2 ANTENNA__14564__B2 (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA__14565__A (.DIODE(net439));
 sky130_fd_sc_hd__diode_2 ANTENNA__14565__B (.DIODE(net434));
 sky130_fd_sc_hd__diode_2 ANTENNA__14565__C (.DIODE(net456));
 sky130_fd_sc_hd__diode_2 ANTENNA__14565__D (.DIODE(net453));
 sky130_fd_sc_hd__diode_2 ANTENNA__14566__A (.DIODE(net429));
 sky130_fd_sc_hd__diode_2 ANTENNA__14566__B (.DIODE(net459));
 sky130_fd_sc_hd__diode_2 ANTENNA__14572__A (.DIODE(net442));
 sky130_fd_sc_hd__diode_2 ANTENNA__14605__A (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__14605__B (.DIODE(_06090_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14606__A1 (.DIODE(net599));
 sky130_fd_sc_hd__diode_2 ANTENNA__14606__B1 (.DIODE(_02653_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14606__B2 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__14614__A1 (.DIODE(net547));
 sky130_fd_sc_hd__diode_2 ANTENNA__14614__A2 (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA__14614__B1 (.DIODE(net331));
 sky130_fd_sc_hd__diode_2 ANTENNA__14614__B2 (.DIODE(net551));
 sky130_fd_sc_hd__diode_2 ANTENNA__14615__A (.DIODE(net547));
 sky130_fd_sc_hd__diode_2 ANTENNA__14615__B (.DIODE(net551));
 sky130_fd_sc_hd__diode_2 ANTENNA__14615__C (.DIODE(net331));
 sky130_fd_sc_hd__diode_2 ANTENNA__14616__A1 (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA__14617__A (.DIODE(net556));
 sky130_fd_sc_hd__diode_2 ANTENNA__14617__B (.DIODE(net329));
 sky130_fd_sc_hd__diode_2 ANTENNA__14619__A1_N (.DIODE(net335));
 sky130_fd_sc_hd__diode_2 ANTENNA__14621__A_N (.DIODE(net563));
 sky130_fd_sc_hd__diode_2 ANTENNA__14621__B (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA__14621__C (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA__14621__D (.DIODE(net560));
 sky130_fd_sc_hd__diode_2 ANTENNA__14623__A1_N (.DIODE(net560));
 sky130_fd_sc_hd__diode_2 ANTENNA__14623__A2_N (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA__14623__B1 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__14623__B2 (.DIODE(net563));
 sky130_fd_sc_hd__diode_2 ANTENNA__14633__A1 (.DIODE(net533));
 sky130_fd_sc_hd__diode_2 ANTENNA__14633__A2 (.DIODE(net349));
 sky130_fd_sc_hd__diode_2 ANTENNA__14634__B1 (.DIODE(net342));
 sky130_fd_sc_hd__diode_2 ANTENNA__14634__B2 (.DIODE(net538));
 sky130_fd_sc_hd__diode_2 ANTENNA__14635__B (.DIODE(net538));
 sky130_fd_sc_hd__diode_2 ANTENNA__14635__D (.DIODE(net341));
 sky130_fd_sc_hd__diode_2 ANTENNA__14636__A1 (.DIODE(net543));
 sky130_fd_sc_hd__diode_2 ANTENNA__14636__A2 (.DIODE(net338));
 sky130_fd_sc_hd__diode_2 ANTENNA__14637__A (.DIODE(net543));
 sky130_fd_sc_hd__diode_2 ANTENNA__14637__B (.DIODE(net338));
 sky130_fd_sc_hd__diode_2 ANTENNA__14651__B (.DIODE(_06098_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14652__A (.DIODE(_06098_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14656__B1 (.DIODE(net352));
 sky130_fd_sc_hd__diode_2 ANTENNA__14657__C (.DIODE(net352));
 sky130_fd_sc_hd__diode_2 ANTENNA__14659__A (.DIODE(net529));
 sky130_fd_sc_hd__diode_2 ANTENNA__14659__B (.DIODE(net349));
 sky130_fd_sc_hd__diode_2 ANTENNA__14661__A1 (.DIODE(net506));
 sky130_fd_sc_hd__diode_2 ANTENNA__14661__B2 (.DIODE(net510));
 sky130_fd_sc_hd__diode_2 ANTENNA__14662__A (.DIODE(net506));
 sky130_fd_sc_hd__diode_2 ANTENNA__14662__B (.DIODE(net510));
 sky130_fd_sc_hd__diode_2 ANTENNA__14663__B (.DIODE(net510));
 sky130_fd_sc_hd__diode_2 ANTENNA__14663__D (.DIODE(net367));
 sky130_fd_sc_hd__diode_2 ANTENNA__14664__A1 (.DIODE(net514));
 sky130_fd_sc_hd__diode_2 ANTENNA__14665__A (.DIODE(net514));
 sky130_fd_sc_hd__diode_2 ANTENNA__14666__A (.DIODE(net514));
 sky130_fd_sc_hd__diode_2 ANTENNA__14672__A1 (.DIODE(net389));
 sky130_fd_sc_hd__diode_2 ANTENNA__14672__A2 (.DIODE(net493));
 sky130_fd_sc_hd__diode_2 ANTENNA__14672__B2 (.DIODE(net484));
 sky130_fd_sc_hd__diode_2 ANTENNA__14673__A1 (.DIODE(net380));
 sky130_fd_sc_hd__diode_2 ANTENNA__14673__A2 (.DIODE(net497));
 sky130_fd_sc_hd__diode_2 ANTENNA__14673__B1 (.DIODE(net493));
 sky130_fd_sc_hd__diode_2 ANTENNA__14673__B2 (.DIODE(net385));
 sky130_fd_sc_hd__diode_2 ANTENNA__14674__A (.DIODE(net385));
 sky130_fd_sc_hd__diode_2 ANTENNA__14674__B (.DIODE(net380));
 sky130_fd_sc_hd__diode_2 ANTENNA__14674__C (.DIODE(net497));
 sky130_fd_sc_hd__diode_2 ANTENNA__14674__D (.DIODE(net493));
 sky130_fd_sc_hd__diode_2 ANTENNA__14675__A1 (.DIODE(net372));
 sky130_fd_sc_hd__diode_2 ANTENNA__14676__A (.DIODE(net372));
 sky130_fd_sc_hd__diode_2 ANTENNA__14692__A1 (.DIODE(net393));
 sky130_fd_sc_hd__diode_2 ANTENNA__14692__A2 (.DIODE(net484));
 sky130_fd_sc_hd__diode_2 ANTENNA__14692__B1 (.DIODE(net479));
 sky130_fd_sc_hd__diode_2 ANTENNA__14692__B2 (.DIODE(net398));
 sky130_fd_sc_hd__diode_2 ANTENNA__14693__A (.DIODE(net398));
 sky130_fd_sc_hd__diode_2 ANTENNA__14693__B (.DIODE(net393));
 sky130_fd_sc_hd__diode_2 ANTENNA__14693__C (.DIODE(net484));
 sky130_fd_sc_hd__diode_2 ANTENNA__14694__A1 (.DIODE(net479));
 sky130_fd_sc_hd__diode_2 ANTENNA__14695__A (.DIODE(net388));
 sky130_fd_sc_hd__diode_2 ANTENNA__14695__B (.DIODE(net488));
 sky130_fd_sc_hd__diode_2 ANTENNA__14697__A1 (.DIODE(\mul0.b[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14697__A2 (.DIODE(net471));
 sky130_fd_sc_hd__diode_2 ANTENNA__14697__B1 (.DIODE(net469));
 sky130_fd_sc_hd__diode_2 ANTENNA__14697__B2 (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA__14698__A (.DIODE(net412));
 sky130_fd_sc_hd__diode_2 ANTENNA__14698__B (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA__14698__C (.DIODE(net471));
 sky130_fd_sc_hd__diode_2 ANTENNA__14698__D (.DIODE(net469));
 sky130_fd_sc_hd__diode_2 ANTENNA__14700__A1 (.DIODE(net402));
 sky130_fd_sc_hd__diode_2 ANTENNA__14701__A (.DIODE(net402));
 sky130_fd_sc_hd__diode_2 ANTENNA__14702__A (.DIODE(net402));
 sky130_fd_sc_hd__diode_2 ANTENNA__14712__A (.DIODE(net439));
 sky130_fd_sc_hd__diode_2 ANTENNA__14712__B (.DIODE(net434));
 sky130_fd_sc_hd__diode_2 ANTENNA__14712__C (.DIODE(net453));
 sky130_fd_sc_hd__diode_2 ANTENNA__14713__A (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA__14713__B (.DIODE(net433));
 sky130_fd_sc_hd__diode_2 ANTENNA__14713__C (.DIODE(net453));
 sky130_fd_sc_hd__diode_2 ANTENNA__14714__A1 (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA__14714__A2 (.DIODE(net433));
 sky130_fd_sc_hd__diode_2 ANTENNA__14714__B1 (.DIODE(net453));
 sky130_fd_sc_hd__diode_2 ANTENNA__14715__A1 (.DIODE(net429));
 sky130_fd_sc_hd__diode_2 ANTENNA__14715__A2 (.DIODE(net456));
 sky130_fd_sc_hd__diode_2 ANTENNA__14716__A (.DIODE(net429));
 sky130_fd_sc_hd__diode_2 ANTENNA__14716__B (.DIODE(net456));
 sky130_fd_sc_hd__diode_2 ANTENNA__14726__A1 (.DIODE(net420));
 sky130_fd_sc_hd__diode_2 ANTENNA__14726__B1 (.DIODE(net459));
 sky130_fd_sc_hd__diode_2 ANTENNA__14726__B2 (.DIODE(net423));
 sky130_fd_sc_hd__diode_2 ANTENNA__14727__A (.DIODE(net424));
 sky130_fd_sc_hd__diode_2 ANTENNA__14727__B (.DIODE(net420));
 sky130_fd_sc_hd__diode_2 ANTENNA__14727__D (.DIODE(net459));
 sky130_fd_sc_hd__diode_2 ANTENNA__14728__A1 (.DIODE(net415));
 sky130_fd_sc_hd__diode_2 ANTENNA__14729__A (.DIODE(net416));
 sky130_fd_sc_hd__diode_2 ANTENNA__14760__A (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__14760__B (.DIODE(_06244_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14761__B1 (.DIODE(_02663_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14761__B2 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__14762__S (.DIODE(_03055_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14767__A1 (.DIODE(net543));
 sky130_fd_sc_hd__diode_2 ANTENNA__14767__A2 (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA__14767__B1 (.DIODE(net331));
 sky130_fd_sc_hd__diode_2 ANTENNA__14767__B2 (.DIODE(net547));
 sky130_fd_sc_hd__diode_2 ANTENNA__14768__A (.DIODE(net543));
 sky130_fd_sc_hd__diode_2 ANTENNA__14768__B (.DIODE(net547));
 sky130_fd_sc_hd__diode_2 ANTENNA__14768__C (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA__14768__D (.DIODE(net331));
 sky130_fd_sc_hd__diode_2 ANTENNA__14770__A (.DIODE(net551));
 sky130_fd_sc_hd__diode_2 ANTENNA__14770__B (.DIODE(net329));
 sky130_fd_sc_hd__diode_2 ANTENNA__14772__A1_N (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA__14774__A_N (.DIODE(net560));
 sky130_fd_sc_hd__diode_2 ANTENNA__14774__B (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA__14774__C (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA__14774__D (.DIODE(net556));
 sky130_fd_sc_hd__diode_2 ANTENNA__14776__A1_N (.DIODE(net556));
 sky130_fd_sc_hd__diode_2 ANTENNA__14776__A2_N (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA__14776__B1 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__14776__B2 (.DIODE(net560));
 sky130_fd_sc_hd__diode_2 ANTENNA__14786__A1 (.DIODE(net528));
 sky130_fd_sc_hd__diode_2 ANTENNA__14786__A2 (.DIODE(net349));
 sky130_fd_sc_hd__diode_2 ANTENNA__14787__A1 (.DIODE(net528));
 sky130_fd_sc_hd__diode_2 ANTENNA__14787__B1 (.DIODE(net342));
 sky130_fd_sc_hd__diode_2 ANTENNA__14788__A (.DIODE(net528));
 sky130_fd_sc_hd__diode_2 ANTENNA__14788__D (.DIODE(net342));
 sky130_fd_sc_hd__diode_2 ANTENNA__14789__A1 (.DIODE(net538));
 sky130_fd_sc_hd__diode_2 ANTENNA__14789__A2 (.DIODE(net338));
 sky130_fd_sc_hd__diode_2 ANTENNA__14790__A (.DIODE(net538));
 sky130_fd_sc_hd__diode_2 ANTENNA__14790__B (.DIODE(net338));
 sky130_fd_sc_hd__diode_2 ANTENNA__14805__A_N (.DIODE(_06250_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14806__A (.DIODE(_06250_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14810__B1 (.DIODE(net352));
 sky130_fd_sc_hd__diode_2 ANTENNA__14811__C (.DIODE(net352));
 sky130_fd_sc_hd__diode_2 ANTENNA__14813__A (.DIODE(net523));
 sky130_fd_sc_hd__diode_2 ANTENNA__14813__B (.DIODE(net349));
 sky130_fd_sc_hd__diode_2 ANTENNA__14815__B2 (.DIODE(net506));
 sky130_fd_sc_hd__diode_2 ANTENNA__14817__A (.DIODE(net506));
 sky130_fd_sc_hd__diode_2 ANTENNA__14818__A1 (.DIODE(net510));
 sky130_fd_sc_hd__diode_2 ANTENNA__14819__A (.DIODE(net510));
 sky130_fd_sc_hd__diode_2 ANTENNA__14820__A (.DIODE(net510));
 sky130_fd_sc_hd__diode_2 ANTENNA__14826__A1 (.DIODE(net388));
 sky130_fd_sc_hd__diode_2 ANTENNA__14826__A2 (.DIODE(net488));
 sky130_fd_sc_hd__diode_2 ANTENNA__14826__B2 (.DIODE(net479));
 sky130_fd_sc_hd__diode_2 ANTENNA__14827__A1 (.DIODE(net378));
 sky130_fd_sc_hd__diode_2 ANTENNA__14827__A2 (.DIODE(net493));
 sky130_fd_sc_hd__diode_2 ANTENNA__14827__B1 (.DIODE(net488));
 sky130_fd_sc_hd__diode_2 ANTENNA__14827__B2 (.DIODE(net384));
 sky130_fd_sc_hd__diode_2 ANTENNA__14828__A (.DIODE(net385));
 sky130_fd_sc_hd__diode_2 ANTENNA__14828__B (.DIODE(net380));
 sky130_fd_sc_hd__diode_2 ANTENNA__14828__C (.DIODE(net493));
 sky130_fd_sc_hd__diode_2 ANTENNA__14828__D (.DIODE(net488));
 sky130_fd_sc_hd__diode_2 ANTENNA__14829__A1 (.DIODE(net372));
 sky130_fd_sc_hd__diode_2 ANTENNA__14829__A2 (.DIODE(net497));
 sky130_fd_sc_hd__diode_2 ANTENNA__14830__A (.DIODE(net372));
 sky130_fd_sc_hd__diode_2 ANTENNA__14830__B (.DIODE(net497));
 sky130_fd_sc_hd__diode_2 ANTENNA__14847__A1 (.DIODE(net428));
 sky130_fd_sc_hd__diode_2 ANTENNA__14847__A2 (.DIODE(net453));
 sky130_fd_sc_hd__diode_2 ANTENNA__14848__A (.DIODE(net428));
 sky130_fd_sc_hd__diode_2 ANTENNA__14855__A1 (.DIODE(net429));
 sky130_fd_sc_hd__diode_2 ANTENNA__14855__A2 (.DIODE(net456));
 sky130_fd_sc_hd__diode_2 ANTENNA__14856__A1 (.DIODE(net419));
 sky130_fd_sc_hd__diode_2 ANTENNA__14856__A2 (.DIODE(\mul0.a[29] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14856__B1 (.DIODE(net456));
 sky130_fd_sc_hd__diode_2 ANTENNA__14856__B2 (.DIODE(net425));
 sky130_fd_sc_hd__diode_2 ANTENNA__14857__A (.DIODE(net424));
 sky130_fd_sc_hd__diode_2 ANTENNA__14857__B (.DIODE(\mul0.b[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14857__C (.DIODE(\mul0.a[29] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14857__D (.DIODE(net456));
 sky130_fd_sc_hd__diode_2 ANTENNA__14858__A1 (.DIODE(net415));
 sky130_fd_sc_hd__diode_2 ANTENNA__14859__A (.DIODE(net415));
 sky130_fd_sc_hd__diode_2 ANTENNA__14870__A1 (.DIODE(net393));
 sky130_fd_sc_hd__diode_2 ANTENNA__14870__A2 (.DIODE(net481));
 sky130_fd_sc_hd__diode_2 ANTENNA__14871__B (.DIODE(net393));
 sky130_fd_sc_hd__diode_2 ANTENNA__14871__C (.DIODE(net479));
 sky130_fd_sc_hd__diode_2 ANTENNA__14872__A1 (.DIODE(net477));
 sky130_fd_sc_hd__diode_2 ANTENNA__14873__A (.DIODE(net388));
 sky130_fd_sc_hd__diode_2 ANTENNA__14873__B (.DIODE(net483));
 sky130_fd_sc_hd__diode_2 ANTENNA__14875__A1 (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA__14875__A2 (.DIODE(net468));
 sky130_fd_sc_hd__diode_2 ANTENNA__14875__B1 (.DIODE(net465));
 sky130_fd_sc_hd__diode_2 ANTENNA__14875__B2 (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA__14876__A (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA__14876__B (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA__14876__C (.DIODE(net468));
 sky130_fd_sc_hd__diode_2 ANTENNA__14876__D (.DIODE(net465));
 sky130_fd_sc_hd__diode_2 ANTENNA__14877__A1 (.DIODE(\mul0.b[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14877__A2 (.DIODE(net471));
 sky130_fd_sc_hd__diode_2 ANTENNA__14878__A (.DIODE(\mul0.b[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14878__B (.DIODE(net471));
 sky130_fd_sc_hd__diode_2 ANTENNA__14916__A (.DIODE(_06398_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14919__B1 (.DIODE(_02671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14919__B2 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__14920__A1 (.DIODE(_03058_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14920__A2 (.DIODE(_06402_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14927__A1 (.DIODE(net538));
 sky130_fd_sc_hd__diode_2 ANTENNA__14927__A2 (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA__14927__B1 (.DIODE(net331));
 sky130_fd_sc_hd__diode_2 ANTENNA__14927__B2 (.DIODE(net543));
 sky130_fd_sc_hd__diode_2 ANTENNA__14928__A (.DIODE(net538));
 sky130_fd_sc_hd__diode_2 ANTENNA__14928__B (.DIODE(net543));
 sky130_fd_sc_hd__diode_2 ANTENNA__14928__C (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA__14928__D (.DIODE(net331));
 sky130_fd_sc_hd__diode_2 ANTENNA__14929__A1 (.DIODE(net547));
 sky130_fd_sc_hd__diode_2 ANTENNA__14929__A2 (.DIODE(net329));
 sky130_fd_sc_hd__diode_2 ANTENNA__14930__A (.DIODE(net547));
 sky130_fd_sc_hd__diode_2 ANTENNA__14930__B (.DIODE(net329));
 sky130_fd_sc_hd__diode_2 ANTENNA__14936__A_N (.DIODE(net556));
 sky130_fd_sc_hd__diode_2 ANTENNA__14936__B (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA__14936__C (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA__14936__D (.DIODE(net551));
 sky130_fd_sc_hd__diode_2 ANTENNA__14938__A1_N (.DIODE(\mul0.a[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14938__A2_N (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA__14938__B1 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__14938__B2 (.DIODE(net556));
 sky130_fd_sc_hd__diode_2 ANTENNA__14947__A2 (.DIODE(net349));
 sky130_fd_sc_hd__diode_2 ANTENNA__14948__B1 (.DIODE(net342));
 sky130_fd_sc_hd__diode_2 ANTENNA__14948__B2 (.DIODE(net528));
 sky130_fd_sc_hd__diode_2 ANTENNA__14949__B (.DIODE(net528));
 sky130_fd_sc_hd__diode_2 ANTENNA__14949__D (.DIODE(net342));
 sky130_fd_sc_hd__diode_2 ANTENNA__14950__A2 (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA__14951__B (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA__14968__A (.DIODE(_06409_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14977__A1 (.DIODE(net429));
 sky130_fd_sc_hd__diode_2 ANTENNA__14978__A1 (.DIODE(net420));
 sky130_fd_sc_hd__diode_2 ANTENNA__14978__A2 (.DIODE(net456));
 sky130_fd_sc_hd__diode_2 ANTENNA__14978__B1 (.DIODE(net453));
 sky130_fd_sc_hd__diode_2 ANTENNA__14978__B2 (.DIODE(net424));
 sky130_fd_sc_hd__diode_2 ANTENNA__14979__A (.DIODE(net424));
 sky130_fd_sc_hd__diode_2 ANTENNA__14979__B (.DIODE(net420));
 sky130_fd_sc_hd__diode_2 ANTENNA__14979__C (.DIODE(net456));
 sky130_fd_sc_hd__diode_2 ANTENNA__14979__D (.DIODE(net453));
 sky130_fd_sc_hd__diode_2 ANTENNA__14980__A1 (.DIODE(net415));
 sky130_fd_sc_hd__diode_2 ANTENNA__14980__A2 (.DIODE(\mul0.a[29] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14981__A (.DIODE(\mul0.b[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14981__B (.DIODE(\mul0.a[29] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__14992__A1 (.DIODE(net393));
 sky130_fd_sc_hd__diode_2 ANTENNA__14992__B1 (.DIODE(net471));
 sky130_fd_sc_hd__diode_2 ANTENNA__14993__B (.DIODE(net394));
 sky130_fd_sc_hd__diode_2 ANTENNA__14993__D (.DIODE(net471));
 sky130_fd_sc_hd__diode_2 ANTENNA__14995__A (.DIODE(net389));
 sky130_fd_sc_hd__diode_2 ANTENNA__14995__B (.DIODE(net479));
 sky130_fd_sc_hd__diode_2 ANTENNA__14997__A1 (.DIODE(net406));
 sky130_fd_sc_hd__diode_2 ANTENNA__14997__A2 (.DIODE(net463));
 sky130_fd_sc_hd__diode_2 ANTENNA__14997__B2 (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA__14998__A (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA__14998__B (.DIODE(net406));
 sky130_fd_sc_hd__diode_2 ANTENNA__14999__A (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA__14999__B (.DIODE(net406));
 sky130_fd_sc_hd__diode_2 ANTENNA__14999__C (.DIODE(net463));
 sky130_fd_sc_hd__diode_2 ANTENNA__15000__A1 (.DIODE(net402));
 sky130_fd_sc_hd__diode_2 ANTENNA__15000__A2 (.DIODE(net466));
 sky130_fd_sc_hd__diode_2 ANTENNA__15001__A (.DIODE(net402));
 sky130_fd_sc_hd__diode_2 ANTENNA__15015__B1 (.DIODE(net352));
 sky130_fd_sc_hd__diode_2 ANTENNA__15016__D (.DIODE(net352));
 sky130_fd_sc_hd__diode_2 ANTENNA__15018__B (.DIODE(net349));
 sky130_fd_sc_hd__diode_2 ANTENNA__15020__B1 (.DIODE(net368));
 sky130_fd_sc_hd__diode_2 ANTENNA__15021__D (.DIODE(net368));
 sky130_fd_sc_hd__diode_2 ANTENNA__15030__A1 (.DIODE(net389));
 sky130_fd_sc_hd__diode_2 ANTENNA__15030__A2 (.DIODE(net483));
 sky130_fd_sc_hd__diode_2 ANTENNA__15031__A1 (.DIODE(net378));
 sky130_fd_sc_hd__diode_2 ANTENNA__15031__A2 (.DIODE(net488));
 sky130_fd_sc_hd__diode_2 ANTENNA__15031__B1 (.DIODE(net484));
 sky130_fd_sc_hd__diode_2 ANTENNA__15031__B2 (.DIODE(net384));
 sky130_fd_sc_hd__diode_2 ANTENNA__15032__A (.DIODE(net384));
 sky130_fd_sc_hd__diode_2 ANTENNA__15032__B (.DIODE(net378));
 sky130_fd_sc_hd__diode_2 ANTENNA__15032__C (.DIODE(net488));
 sky130_fd_sc_hd__diode_2 ANTENNA__15032__D (.DIODE(net484));
 sky130_fd_sc_hd__diode_2 ANTENNA__15033__A1 (.DIODE(net373));
 sky130_fd_sc_hd__diode_2 ANTENNA__15033__A2 (.DIODE(net493));
 sky130_fd_sc_hd__diode_2 ANTENNA__15034__A (.DIODE(net373));
 sky130_fd_sc_hd__diode_2 ANTENNA__15034__B (.DIODE(net493));
 sky130_fd_sc_hd__diode_2 ANTENNA__15048__B1 (.DIODE(_06529_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15049__A1 (.DIODE(_06529_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15050__C (.DIODE(_06531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15051__B1 (.DIODE(_06531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15070__A (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__15070__B (.DIODE(_06552_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15071__B1 (.DIODE(_02677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15071__B2 (.DIODE(_03794_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15072__S (.DIODE(_03055_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15074__A1 (.DIODE(_06409_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15076__A (.DIODE(net424));
 sky130_fd_sc_hd__diode_2 ANTENNA__15076__B (.DIODE(net420));
 sky130_fd_sc_hd__diode_2 ANTENNA__15076__C (.DIODE(net453));
 sky130_fd_sc_hd__diode_2 ANTENNA__15077__A1 (.DIODE(net424));
 sky130_fd_sc_hd__diode_2 ANTENNA__15077__A2 (.DIODE(net420));
 sky130_fd_sc_hd__diode_2 ANTENNA__15077__B1 (.DIODE(net453));
 sky130_fd_sc_hd__diode_2 ANTENNA__15078__A1 (.DIODE(net416));
 sky130_fd_sc_hd__diode_2 ANTENNA__15078__A2 (.DIODE(net456));
 sky130_fd_sc_hd__diode_2 ANTENNA__15079__A (.DIODE(net416));
 sky130_fd_sc_hd__diode_2 ANTENNA__15079__B (.DIODE(net456));
 sky130_fd_sc_hd__diode_2 ANTENNA__15090__A1 (.DIODE(net393));
 sky130_fd_sc_hd__diode_2 ANTENNA__15090__A2 (.DIODE(net473));
 sky130_fd_sc_hd__diode_2 ANTENNA__15090__B2 (.DIODE(net398));
 sky130_fd_sc_hd__diode_2 ANTENNA__15091__A (.DIODE(net398));
 sky130_fd_sc_hd__diode_2 ANTENNA__15091__B (.DIODE(net393));
 sky130_fd_sc_hd__diode_2 ANTENNA__15091__C (.DIODE(net473));
 sky130_fd_sc_hd__diode_2 ANTENNA__15093__A (.DIODE(net388));
 sky130_fd_sc_hd__diode_2 ANTENNA__15093__B (.DIODE(net477));
 sky130_fd_sc_hd__diode_2 ANTENNA__15095__A1 (.DIODE(net406));
 sky130_fd_sc_hd__diode_2 ANTENNA__15095__B1 (.DIODE(net459));
 sky130_fd_sc_hd__diode_2 ANTENNA__15095__B2 (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA__15096__A (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA__15096__B (.DIODE(net406));
 sky130_fd_sc_hd__diode_2 ANTENNA__15096__D (.DIODE(net459));
 sky130_fd_sc_hd__diode_2 ANTENNA__15097__A1 (.DIODE(net402));
 sky130_fd_sc_hd__diode_2 ANTENNA__15097__A2 (.DIODE(net463));
 sky130_fd_sc_hd__diode_2 ANTENNA__15098__A (.DIODE(net402));
 sky130_fd_sc_hd__diode_2 ANTENNA__15098__B (.DIODE(net463));
 sky130_fd_sc_hd__diode_2 ANTENNA__15111__B1 (.DIODE(net352));
 sky130_fd_sc_hd__diode_2 ANTENNA__15112__D (.DIODE(net352));
 sky130_fd_sc_hd__diode_2 ANTENNA__15114__A2 (.DIODE(net349));
 sky130_fd_sc_hd__diode_2 ANTENNA__15115__B (.DIODE(net349));
 sky130_fd_sc_hd__diode_2 ANTENNA__15117__A2 (.DIODE(net368));
 sky130_fd_sc_hd__diode_2 ANTENNA__15118__C (.DIODE(net368));
 sky130_fd_sc_hd__diode_2 ANTENNA__15120__B (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 ANTENNA__15129__A1 (.DIODE(net378));
 sky130_fd_sc_hd__diode_2 ANTENNA__15129__A2 (.DIODE(net484));
 sky130_fd_sc_hd__diode_2 ANTENNA__15129__B1 (.DIODE(net479));
 sky130_fd_sc_hd__diode_2 ANTENNA__15129__B2 (.DIODE(net384));
 sky130_fd_sc_hd__diode_2 ANTENNA__15130__A (.DIODE(net385));
 sky130_fd_sc_hd__diode_2 ANTENNA__15130__B (.DIODE(net379));
 sky130_fd_sc_hd__diode_2 ANTENNA__15130__C (.DIODE(net484));
 sky130_fd_sc_hd__diode_2 ANTENNA__15130__D (.DIODE(net479));
 sky130_fd_sc_hd__diode_2 ANTENNA__15131__A1_N (.DIODE(net373));
 sky130_fd_sc_hd__diode_2 ANTENNA__15131__A2_N (.DIODE(net488));
 sky130_fd_sc_hd__diode_2 ANTENNA__15132__C (.DIODE(net373));
 sky130_fd_sc_hd__diode_2 ANTENNA__15132__D (.DIODE(net488));
 sky130_fd_sc_hd__diode_2 ANTENNA__15151__A (.DIODE(_06631_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15152__A2 (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA__15152__B1 (.DIODE(net331));
 sky130_fd_sc_hd__diode_2 ANTENNA__15152__B2 (.DIODE(net538));
 sky130_fd_sc_hd__diode_2 ANTENNA__15153__A (.DIODE(net533));
 sky130_fd_sc_hd__diode_2 ANTENNA__15153__B (.DIODE(net538));
 sky130_fd_sc_hd__diode_2 ANTENNA__15153__C (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA__15153__D (.DIODE(net331));
 sky130_fd_sc_hd__diode_2 ANTENNA__15154__A1_N (.DIODE(net543));
 sky130_fd_sc_hd__diode_2 ANTENNA__15154__A2_N (.DIODE(net329));
 sky130_fd_sc_hd__diode_2 ANTENNA__15155__C (.DIODE(net543));
 sky130_fd_sc_hd__diode_2 ANTENNA__15155__D (.DIODE(net329));
 sky130_fd_sc_hd__diode_2 ANTENNA__15159__A_N (.DIODE(\mul0.a[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15159__B (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA__15159__C (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA__15159__D (.DIODE(net547));
 sky130_fd_sc_hd__diode_2 ANTENNA__15161__A1_N (.DIODE(\mul0.a[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15161__A2_N (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA__15161__B1 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__15161__B2 (.DIODE(\mul0.a[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15171__B1 (.DIODE(net342));
 sky130_fd_sc_hd__diode_2 ANTENNA__15172__D (.DIODE(net342));
 sky130_fd_sc_hd__diode_2 ANTENNA__15173__A1_N (.DIODE(net528));
 sky130_fd_sc_hd__diode_2 ANTENNA__15173__A2_N (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA__15174__C (.DIODE(net528));
 sky130_fd_sc_hd__diode_2 ANTENNA__15174__D (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA__15187__A1 (.DIODE(_06529_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15187__A2 (.DIODE(_06531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15188__B1 (.DIODE(_06529_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15188__C1 (.DIODE(_06531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15192__A (.DIODE(_06633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15210__A (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__15210__B (.DIODE(_06691_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15211__B1 (.DIODE(_02683_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15211__B2 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__15216__A1 (.DIODE(net416));
 sky130_fd_sc_hd__diode_2 ANTENNA__15217__A (.DIODE(net416));
 sky130_fd_sc_hd__diode_2 ANTENNA__15228__A1 (.DIODE(net393));
 sky130_fd_sc_hd__diode_2 ANTENNA__15228__A2 (.DIODE(net468));
 sky130_fd_sc_hd__diode_2 ANTENNA__15228__B1 (.DIODE(net465));
 sky130_fd_sc_hd__diode_2 ANTENNA__15228__B2 (.DIODE(net398));
 sky130_fd_sc_hd__diode_2 ANTENNA__15229__A (.DIODE(net398));
 sky130_fd_sc_hd__diode_2 ANTENNA__15229__B (.DIODE(net393));
 sky130_fd_sc_hd__diode_2 ANTENNA__15229__C (.DIODE(net466));
 sky130_fd_sc_hd__diode_2 ANTENNA__15229__D (.DIODE(net465));
 sky130_fd_sc_hd__diode_2 ANTENNA__15230__A1 (.DIODE(net388));
 sky130_fd_sc_hd__diode_2 ANTENNA__15230__A2 (.DIODE(net470));
 sky130_fd_sc_hd__diode_2 ANTENNA__15231__A (.DIODE(net388));
 sky130_fd_sc_hd__diode_2 ANTENNA__15231__B (.DIODE(net471));
 sky130_fd_sc_hd__diode_2 ANTENNA__15233__A1 (.DIODE(net406));
 sky130_fd_sc_hd__diode_2 ANTENNA__15233__B2 (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA__15234__A (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA__15234__B (.DIODE(net406));
 sky130_fd_sc_hd__diode_2 ANTENNA__15234__C (.DIODE(net459));
 sky130_fd_sc_hd__diode_2 ANTENNA__15235__A1_N (.DIODE(net402));
 sky130_fd_sc_hd__diode_2 ANTENNA__15236__C (.DIODE(net402));
 sky130_fd_sc_hd__diode_2 ANTENNA__15246__A (.DIODE(_06726_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15255__B2 (.DIODE(net506));
 sky130_fd_sc_hd__diode_2 ANTENNA__15260__A1 (.DIODE(net368));
 sky130_fd_sc_hd__diode_2 ANTENNA__15261__B (.DIODE(net368));
 sky130_fd_sc_hd__diode_2 ANTENNA__15263__A2 (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 ANTENNA__15264__A (.DIODE(net497));
 sky130_fd_sc_hd__diode_2 ANTENNA__15264__B (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 ANTENNA__15273__A1 (.DIODE(net378));
 sky130_fd_sc_hd__diode_2 ANTENNA__15273__B2 (.DIODE(net384));
 sky130_fd_sc_hd__diode_2 ANTENNA__15274__A (.DIODE(net384));
 sky130_fd_sc_hd__diode_2 ANTENNA__15274__B (.DIODE(net378));
 sky130_fd_sc_hd__diode_2 ANTENNA__15275__A1_N (.DIODE(net373));
 sky130_fd_sc_hd__diode_2 ANTENNA__15276__C (.DIODE(net372));
 sky130_fd_sc_hd__diode_2 ANTENNA__15278__A (.DIODE(_06753_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15279__A (.DIODE(_06753_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15280__A (.DIODE(_06752_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15281__A (.DIODE(_06752_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15283__B (.DIODE(_06763_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15284__B (.DIODE(_06763_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15299__A1 (.DIODE(net528));
 sky130_fd_sc_hd__diode_2 ANTENNA__15299__A2 (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA__15299__B1 (.DIODE(net331));
 sky130_fd_sc_hd__diode_2 ANTENNA__15299__B2 (.DIODE(net533));
 sky130_fd_sc_hd__diode_2 ANTENNA__15300__A (.DIODE(net528));
 sky130_fd_sc_hd__diode_2 ANTENNA__15300__B (.DIODE(net533));
 sky130_fd_sc_hd__diode_2 ANTENNA__15300__C (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA__15300__D (.DIODE(net331));
 sky130_fd_sc_hd__diode_2 ANTENNA__15302__A1 (.DIODE(net539));
 sky130_fd_sc_hd__diode_2 ANTENNA__15302__A2 (.DIODE(net329));
 sky130_fd_sc_hd__diode_2 ANTENNA__15303__A (.DIODE(net539));
 sky130_fd_sc_hd__diode_2 ANTENNA__15303__B (.DIODE(net329));
 sky130_fd_sc_hd__diode_2 ANTENNA__15308__A_N (.DIODE(\mul0.a[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15308__B (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA__15308__C (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA__15308__D (.DIODE(\mul0.a[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15309__A1_N (.DIODE(\mul0.a[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15309__A2_N (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA__15309__B1 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__15309__B2 (.DIODE(net547));
 sky130_fd_sc_hd__diode_2 ANTENNA__15317__A2 (.DIODE(net349));
 sky130_fd_sc_hd__diode_2 ANTENNA__15318__B1 (.DIODE(net342));
 sky130_fd_sc_hd__diode_2 ANTENNA__15319__D (.DIODE(net342));
 sky130_fd_sc_hd__diode_2 ANTENNA__15320__A2_N (.DIODE(net338));
 sky130_fd_sc_hd__diode_2 ANTENNA__15321__D (.DIODE(net338));
 sky130_fd_sc_hd__diode_2 ANTENNA__15336__A (.DIODE(_06779_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15337__B1 (.DIODE(_06779_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15343__A1 (.DIODE(_06633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15343__B1 (.DIODE(_06631_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15357__B1 (.DIODE(_02690_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15357__B2 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__15358__A1 (.DIODE(_03058_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15358__A2 (.DIODE(_06837_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15367__A1 (.DIODE(net393));
 sky130_fd_sc_hd__diode_2 ANTENNA__15367__B2 (.DIODE(net398));
 sky130_fd_sc_hd__diode_2 ANTENNA__15368__A (.DIODE(net398));
 sky130_fd_sc_hd__diode_2 ANTENNA__15368__B (.DIODE(net393));
 sky130_fd_sc_hd__diode_2 ANTENNA__15369__A1 (.DIODE(net388));
 sky130_fd_sc_hd__diode_2 ANTENNA__15369__A2 (.DIODE(net466));
 sky130_fd_sc_hd__diode_2 ANTENNA__15370__A (.DIODE(net388));
 sky130_fd_sc_hd__diode_2 ANTENNA__15370__B (.DIODE(net466));
 sky130_fd_sc_hd__diode_2 ANTENNA__15372__A1 (.DIODE(net406));
 sky130_fd_sc_hd__diode_2 ANTENNA__15372__B2 (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA__15373__A (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA__15373__B (.DIODE(net406));
 sky130_fd_sc_hd__diode_2 ANTENNA__15375__A (.DIODE(net402));
 sky130_fd_sc_hd__diode_2 ANTENNA__15385__A1 (.DIODE(_06863_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15386__B (.DIODE(_06863_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15394__A1 (.DIODE(net368));
 sky130_fd_sc_hd__diode_2 ANTENNA__15395__B (.DIODE(net368));
 sky130_fd_sc_hd__diode_2 ANTENNA__15397__A2 (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 ANTENNA__15398__B (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 ANTENNA__15408__A1 (.DIODE(net378));
 sky130_fd_sc_hd__diode_2 ANTENNA__15408__B1 (.DIODE(net471));
 sky130_fd_sc_hd__diode_2 ANTENNA__15408__B2 (.DIODE(net384));
 sky130_fd_sc_hd__diode_2 ANTENNA__15410__A (.DIODE(net384));
 sky130_fd_sc_hd__diode_2 ANTENNA__15410__B (.DIODE(net378));
 sky130_fd_sc_hd__diode_2 ANTENNA__15410__D (.DIODE(net471));
 sky130_fd_sc_hd__diode_2 ANTENNA__15411__A1_N (.DIODE(net372));
 sky130_fd_sc_hd__diode_2 ANTENNA__15412__C (.DIODE(net373));
 sky130_fd_sc_hd__diode_2 ANTENNA__15414__B (.DIODE(_06887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15415__A (.DIODE(_06887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15422__A1 (.DIODE(_06724_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15423__B1 (.DIODE(_06724_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15426__A (.DIODE(_06867_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15426__B (.DIODE(_06868_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15427__A1 (.DIODE(_06867_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15427__A2 (.DIODE(_06868_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15431__A1 (.DIODE(net523));
 sky130_fd_sc_hd__diode_2 ANTENNA__15431__A2 (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA__15431__B1 (.DIODE(net331));
 sky130_fd_sc_hd__diode_2 ANTENNA__15431__B2 (.DIODE(net528));
 sky130_fd_sc_hd__diode_2 ANTENNA__15432__B (.DIODE(net528));
 sky130_fd_sc_hd__diode_2 ANTENNA__15432__C (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA__15432__D (.DIODE(net331));
 sky130_fd_sc_hd__diode_2 ANTENNA__15434__A1 (.DIODE(net533));
 sky130_fd_sc_hd__diode_2 ANTENNA__15434__A2 (.DIODE(net329));
 sky130_fd_sc_hd__diode_2 ANTENNA__15435__A (.DIODE(net533));
 sky130_fd_sc_hd__diode_2 ANTENNA__15435__B (.DIODE(net329));
 sky130_fd_sc_hd__diode_2 ANTENNA__15439__A_N (.DIODE(\mul0.a[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15439__B (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA__15439__C (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA__15439__D (.DIODE(net539));
 sky130_fd_sc_hd__diode_2 ANTENNA__15441__A1_N (.DIODE(net539));
 sky130_fd_sc_hd__diode_2 ANTENNA__15441__A2_N (.DIODE(net328));
 sky130_fd_sc_hd__diode_2 ANTENNA__15441__B1 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__15441__B2 (.DIODE(\mul0.a[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15452__B1 (.DIODE(net342));
 sky130_fd_sc_hd__diode_2 ANTENNA__15454__B (.DIODE(net514));
 sky130_fd_sc_hd__diode_2 ANTENNA__15454__D (.DIODE(net342));
 sky130_fd_sc_hd__diode_2 ANTENNA__15455__A2_N (.DIODE(net338));
 sky130_fd_sc_hd__diode_2 ANTENNA__15456__B (.DIODE(net338));
 sky130_fd_sc_hd__diode_2 ANTENNA__15493__A1 (.DIODE(_06398_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15498__B1 (.DIODE(_02696_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15498__B2 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__15499__A1 (.DIODE(_03058_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15499__A2 (.DIODE(_06977_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15503__A (.DIODE(_06980_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15504__A (.DIODE(_06980_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15507__A1 (.DIODE(net393));
 sky130_fd_sc_hd__diode_2 ANTENNA__15507__A2 (.DIODE(net462));
 sky130_fd_sc_hd__diode_2 ANTENNA__15507__B2 (.DIODE(net398));
 sky130_fd_sc_hd__diode_2 ANTENNA__15508__A (.DIODE(net398));
 sky130_fd_sc_hd__diode_2 ANTENNA__15508__B (.DIODE(net393));
 sky130_fd_sc_hd__diode_2 ANTENNA__15508__C (.DIODE(net462));
 sky130_fd_sc_hd__diode_2 ANTENNA__15509__A1 (.DIODE(net388));
 sky130_fd_sc_hd__diode_2 ANTENNA__15509__A2 (.DIODE(net465));
 sky130_fd_sc_hd__diode_2 ANTENNA__15510__A (.DIODE(net388));
 sky130_fd_sc_hd__diode_2 ANTENNA__15512__A1 (.DIODE(net402));
 sky130_fd_sc_hd__diode_2 ANTENNA__15513__A (.DIODE(net403));
 sky130_fd_sc_hd__diode_2 ANTENNA__15514__A (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA__15514__B (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA__15514__C (.DIODE(net453));
 sky130_fd_sc_hd__diode_2 ANTENNA__15515__A1 (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA__15515__A2 (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA__15515__B1 (.DIODE(net453));
 sky130_fd_sc_hd__diode_2 ANTENNA__15520__A (.DIODE(_06985_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15520__B (.DIODE(_06998_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15521__A (.DIODE(_06985_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15521__B (.DIODE(_06998_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15522__B (.DIODE(_06984_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15523__A (.DIODE(_06984_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15524__A (.DIODE(_06983_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15525__A (.DIODE(_06983_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15528__B (.DIODE(_07006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15529__B (.DIODE(_07006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15531__A (.DIODE(net497));
 sky130_fd_sc_hd__diode_2 ANTENNA__15535__A1 (.DIODE(net369));
 sky130_fd_sc_hd__diode_2 ANTENNA__15535__B1 (.DIODE(net479));
 sky130_fd_sc_hd__diode_2 ANTENNA__15536__B (.DIODE(net369));
 sky130_fd_sc_hd__diode_2 ANTENNA__15538__A1 (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 ANTENNA__15539__A (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 ANTENNA__15549__A1 (.DIODE(net378));
 sky130_fd_sc_hd__diode_2 ANTENNA__15549__A2 (.DIODE(net471));
 sky130_fd_sc_hd__diode_2 ANTENNA__15549__B1 (.DIODE(net469));
 sky130_fd_sc_hd__diode_2 ANTENNA__15549__B2 (.DIODE(net384));
 sky130_fd_sc_hd__diode_2 ANTENNA__15551__A (.DIODE(net384));
 sky130_fd_sc_hd__diode_2 ANTENNA__15551__B (.DIODE(net378));
 sky130_fd_sc_hd__diode_2 ANTENNA__15551__D (.DIODE(net468));
 sky130_fd_sc_hd__diode_2 ANTENNA__15552__A1_N (.DIODE(net372));
 sky130_fd_sc_hd__diode_2 ANTENNA__15553__C (.DIODE(net372));
 sky130_fd_sc_hd__diode_2 ANTENNA__15555__B (.DIODE(_07027_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15556__A (.DIODE(_07027_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15563__A1 (.DIODE(_06861_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15563__A2 (.DIODE(_06863_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15564__B1 (.DIODE(_06861_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15564__C1 (.DIODE(_06863_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15569__A1 (.DIODE(_06868_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15570__B1 (.DIODE(_06868_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15571__A1 (.DIODE(net519));
 sky130_fd_sc_hd__diode_2 ANTENNA__15571__A2 (.DIODE(net335));
 sky130_fd_sc_hd__diode_2 ANTENNA__15571__B1 (.DIODE(net331));
 sky130_fd_sc_hd__diode_2 ANTENNA__15572__A (.DIODE(\mul0.a[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15572__C (.DIODE(net335));
 sky130_fd_sc_hd__diode_2 ANTENNA__15572__D (.DIODE(net332));
 sky130_fd_sc_hd__diode_2 ANTENNA__15574__A1 (.DIODE(net528));
 sky130_fd_sc_hd__diode_2 ANTENNA__15574__A2 (.DIODE(net329));
 sky130_fd_sc_hd__diode_2 ANTENNA__15575__A (.DIODE(net528));
 sky130_fd_sc_hd__diode_2 ANTENNA__15575__B (.DIODE(\mul0.b[29] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15579__A_N (.DIODE(net539));
 sky130_fd_sc_hd__diode_2 ANTENNA__15579__C (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA__15580__A1_N (.DIODE(net533));
 sky130_fd_sc_hd__diode_2 ANTENNA__15580__B1 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__15580__B2 (.DIODE(net539));
 sky130_fd_sc_hd__diode_2 ANTENNA__15589__A1 (.DIODE(net506));
 sky130_fd_sc_hd__diode_2 ANTENNA__15589__B1 (.DIODE(net342));
 sky130_fd_sc_hd__diode_2 ANTENNA__15591__A (.DIODE(net506));
 sky130_fd_sc_hd__diode_2 ANTENNA__15591__D (.DIODE(net342));
 sky130_fd_sc_hd__diode_2 ANTENNA__15592__A1_N (.DIODE(net514));
 sky130_fd_sc_hd__diode_2 ANTENNA__15592__A2_N (.DIODE(net338));
 sky130_fd_sc_hd__diode_2 ANTENNA__15593__B (.DIODE(net338));
 sky130_fd_sc_hd__diode_2 ANTENNA__15627__A1 (.DIODE(net599));
 sky130_fd_sc_hd__diode_2 ANTENNA__15627__B1 (.DIODE(_02700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15627__B2 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__15628__A1 (.DIODE(_03058_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15628__A2 (.DIODE(_07105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15631__A1 (.DIODE(net393));
 sky130_fd_sc_hd__diode_2 ANTENNA__15631__B2 (.DIODE(net398));
 sky130_fd_sc_hd__diode_2 ANTENNA__15632__A (.DIODE(net398));
 sky130_fd_sc_hd__diode_2 ANTENNA__15632__B (.DIODE(net393));
 sky130_fd_sc_hd__diode_2 ANTENNA__15632__D (.DIODE(net456));
 sky130_fd_sc_hd__diode_2 ANTENNA__15634__A1 (.DIODE(net388));
 sky130_fd_sc_hd__diode_2 ANTENNA__15634__A2 (.DIODE(net462));
 sky130_fd_sc_hd__diode_2 ANTENNA__15635__A (.DIODE(net388));
 sky130_fd_sc_hd__diode_2 ANTENNA__15635__B (.DIODE(net462));
 sky130_fd_sc_hd__diode_2 ANTENNA__15637__A1 (.DIODE(net403));
 sky130_fd_sc_hd__diode_2 ANTENNA__15639__A1 (.DIODE(net403));
 sky130_fd_sc_hd__diode_2 ANTENNA__15642__A (.DIODE(_06985_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15642__B (.DIODE(_07119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15643__A (.DIODE(_06985_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15643__B (.DIODE(_07119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15644__A (.DIODE(_07108_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15645__A (.DIODE(_07108_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15646__A (.DIODE(_06983_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15648__A (.DIODE(_06980_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15649__A1 (.DIODE(_06980_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15654__A1 (.DIODE(net497));
 sky130_fd_sc_hd__diode_2 ANTENNA__15655__A (.DIODE(net497));
 sky130_fd_sc_hd__diode_2 ANTENNA__15657__A1 (.DIODE(net369));
 sky130_fd_sc_hd__diode_2 ANTENNA__15658__B (.DIODE(net369));
 sky130_fd_sc_hd__diode_2 ANTENNA__15660__A1 (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 ANTENNA__15660__A2 (.DIODE(net484));
 sky130_fd_sc_hd__diode_2 ANTENNA__15661__A (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 ANTENNA__15661__B (.DIODE(net484));
 sky130_fd_sc_hd__diode_2 ANTENNA__15671__A1 (.DIODE(net378));
 sky130_fd_sc_hd__diode_2 ANTENNA__15671__A2 (.DIODE(net469));
 sky130_fd_sc_hd__diode_2 ANTENNA__15671__B1 (.DIODE(net465));
 sky130_fd_sc_hd__diode_2 ANTENNA__15671__B2 (.DIODE(net384));
 sky130_fd_sc_hd__diode_2 ANTENNA__15673__A (.DIODE(net384));
 sky130_fd_sc_hd__diode_2 ANTENNA__15673__B (.DIODE(net378));
 sky130_fd_sc_hd__diode_2 ANTENNA__15673__C (.DIODE(net468));
 sky130_fd_sc_hd__diode_2 ANTENNA__15673__D (.DIODE(net465));
 sky130_fd_sc_hd__diode_2 ANTENNA__15674__A1_N (.DIODE(net373));
 sky130_fd_sc_hd__diode_2 ANTENNA__15675__C (.DIODE(net372));
 sky130_fd_sc_hd__diode_2 ANTENNA__15677__B (.DIODE(_07148_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15678__A (.DIODE(_07148_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15694__A1 (.DIODE(net514));
 sky130_fd_sc_hd__diode_2 ANTENNA__15694__A2 (.DIODE(net335));
 sky130_fd_sc_hd__diode_2 ANTENNA__15694__B1 (.DIODE(net332));
 sky130_fd_sc_hd__diode_2 ANTENNA__15695__A (.DIODE(net514));
 sky130_fd_sc_hd__diode_2 ANTENNA__15695__C (.DIODE(net335));
 sky130_fd_sc_hd__diode_2 ANTENNA__15695__D (.DIODE(net332));
 sky130_fd_sc_hd__diode_2 ANTENNA__15697__A2 (.DIODE(net329));
 sky130_fd_sc_hd__diode_2 ANTENNA__15698__B (.DIODE(net329));
 sky130_fd_sc_hd__diode_2 ANTENNA__15702__A_N (.DIODE(net533));
 sky130_fd_sc_hd__diode_2 ANTENNA__15702__B (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA__15702__C (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA__15702__D (.DIODE(net528));
 sky130_fd_sc_hd__diode_2 ANTENNA__15704__A1_N (.DIODE(net528));
 sky130_fd_sc_hd__diode_2 ANTENNA__15704__A2_N (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA__15704__B1 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__15704__B2 (.DIODE(net533));
 sky130_fd_sc_hd__diode_2 ANTENNA__15715__B1 (.DIODE(net342));
 sky130_fd_sc_hd__diode_2 ANTENNA__15717__D (.DIODE(net342));
 sky130_fd_sc_hd__diode_2 ANTENNA__15718__A2_N (.DIODE(net338));
 sky130_fd_sc_hd__diode_2 ANTENNA__15719__B (.DIODE(net338));
 sky130_fd_sc_hd__diode_2 ANTENNA__15759__A (.DIODE(_03057_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15760__A1 (.DIODE(net600));
 sky130_fd_sc_hd__diode_2 ANTENNA__15760__B1 (.DIODE(_02703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15760__B2 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__15761__S (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__15762__A (.DIODE(net403));
 sky130_fd_sc_hd__diode_2 ANTENNA__15763__A (.DIODE(net403));
 sky130_fd_sc_hd__diode_2 ANTENNA__15765__A1 (.DIODE(net394));
 sky130_fd_sc_hd__diode_2 ANTENNA__15765__B1 (.DIODE(net453));
 sky130_fd_sc_hd__diode_2 ANTENNA__15765__B2 (.DIODE(net398));
 sky130_fd_sc_hd__diode_2 ANTENNA__15766__A (.DIODE(net398));
 sky130_fd_sc_hd__diode_2 ANTENNA__15766__B (.DIODE(net394));
 sky130_fd_sc_hd__diode_2 ANTENNA__15766__D (.DIODE(net453));
 sky130_fd_sc_hd__diode_2 ANTENNA__15768__A (.DIODE(net389));
 sky130_fd_sc_hd__diode_2 ANTENNA__15774__A (.DIODE(_06985_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15775__A (.DIODE(_06985_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15779__A (.DIODE(_06983_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15780__A (.DIODE(_06983_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15782__A (.DIODE(_06980_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15783__A1 (.DIODE(_06980_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15786__A (.DIODE(net488));
 sky130_fd_sc_hd__diode_2 ANTENNA__15787__A1 (.DIODE(net493));
 sky130_fd_sc_hd__diode_2 ANTENNA__15787__A2 (.DIODE(net349));
 sky130_fd_sc_hd__diode_2 ANTENNA__15788__A (.DIODE(net493));
 sky130_fd_sc_hd__diode_2 ANTENNA__15788__B (.DIODE(net349));
 sky130_fd_sc_hd__diode_2 ANTENNA__15790__A1 (.DIODE(net369));
 sky130_fd_sc_hd__diode_2 ANTENNA__15791__B (.DIODE(net369));
 sky130_fd_sc_hd__diode_2 ANTENNA__15793__A1 (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 ANTENNA__15794__A (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 ANTENNA__15804__A1 (.DIODE(net378));
 sky130_fd_sc_hd__diode_2 ANTENNA__15804__A2 (.DIODE(net465));
 sky130_fd_sc_hd__diode_2 ANTENNA__15804__B1 (.DIODE(net462));
 sky130_fd_sc_hd__diode_2 ANTENNA__15804__B2 (.DIODE(net384));
 sky130_fd_sc_hd__diode_2 ANTENNA__15806__A (.DIODE(net384));
 sky130_fd_sc_hd__diode_2 ANTENNA__15806__B (.DIODE(net378));
 sky130_fd_sc_hd__diode_2 ANTENNA__15806__C (.DIODE(net465));
 sky130_fd_sc_hd__diode_2 ANTENNA__15806__D (.DIODE(net462));
 sky130_fd_sc_hd__diode_2 ANTENNA__15807__A1_N (.DIODE(net372));
 sky130_fd_sc_hd__diode_2 ANTENNA__15807__A2_N (.DIODE(net468));
 sky130_fd_sc_hd__diode_2 ANTENNA__15808__B (.DIODE(net468));
 sky130_fd_sc_hd__diode_2 ANTENNA__15808__C (.DIODE(net372));
 sky130_fd_sc_hd__diode_2 ANTENNA__15828__A2 (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA__15828__B1 (.DIODE(net332));
 sky130_fd_sc_hd__diode_2 ANTENNA__15828__B2 (.DIODE(net514));
 sky130_fd_sc_hd__diode_2 ANTENNA__15829__A (.DIODE(net510));
 sky130_fd_sc_hd__diode_2 ANTENNA__15829__C (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA__15829__D (.DIODE(net332));
 sky130_fd_sc_hd__diode_2 ANTENNA__15831__A2 (.DIODE(net330));
 sky130_fd_sc_hd__diode_2 ANTENNA__15832__B (.DIODE(net330));
 sky130_fd_sc_hd__diode_2 ANTENNA__15838__A_N (.DIODE(net528));
 sky130_fd_sc_hd__diode_2 ANTENNA__15838__B (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA__15838__C (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA__15839__A2_N (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA__15839__B2 (.DIODE(net529));
 sky130_fd_sc_hd__diode_2 ANTENNA__15850__A2 (.DIODE(net347));
 sky130_fd_sc_hd__diode_2 ANTENNA__15850__B1 (.DIODE(net343));
 sky130_fd_sc_hd__diode_2 ANTENNA__15852__C (.DIODE(net347));
 sky130_fd_sc_hd__diode_2 ANTENNA__15852__D (.DIODE(net343));
 sky130_fd_sc_hd__diode_2 ANTENNA__15853__A2_N (.DIODE(net338));
 sky130_fd_sc_hd__diode_2 ANTENNA__15854__B (.DIODE(net338));
 sky130_fd_sc_hd__diode_2 ANTENNA__15889__A1 (.DIODE(net600));
 sky130_fd_sc_hd__diode_2 ANTENNA__15889__B1 (.DIODE(_02711_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15889__B2 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__15890__A1 (.DIODE(_03058_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15890__A2 (.DIODE(_07365_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15891__S (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__15892__A (.DIODE(net398));
 sky130_fd_sc_hd__diode_2 ANTENNA__15892__B (.DIODE(net394));
 sky130_fd_sc_hd__diode_2 ANTENNA__15893__A1 (.DIODE(net398));
 sky130_fd_sc_hd__diode_2 ANTENNA__15893__A2 (.DIODE(net393));
 sky130_fd_sc_hd__diode_2 ANTENNA__15895__A (.DIODE(net388));
 sky130_fd_sc_hd__diode_2 ANTENNA__15895__B (.DIODE(net456));
 sky130_fd_sc_hd__diode_2 ANTENNA__15900__A (.DIODE(_06985_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15901__A (.DIODE(_06985_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15907__A (.DIODE(_06980_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15908__A1 (.DIODE(_06980_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15910__A1 (.DIODE(net484));
 sky130_fd_sc_hd__diode_2 ANTENNA__15912__A1 (.DIODE(net488));
 sky130_fd_sc_hd__diode_2 ANTENNA__15912__A2 (.DIODE(net349));
 sky130_fd_sc_hd__diode_2 ANTENNA__15915__A1 (.DIODE(net368));
 sky130_fd_sc_hd__diode_2 ANTENNA__15915__B1 (.DIODE(net468));
 sky130_fd_sc_hd__diode_2 ANTENNA__15915__B2 (.DIODE(net635));
 sky130_fd_sc_hd__diode_2 ANTENNA__15916__A (.DIODE(net635));
 sky130_fd_sc_hd__diode_2 ANTENNA__15916__B (.DIODE(net369));
 sky130_fd_sc_hd__diode_2 ANTENNA__15916__D (.DIODE(net468));
 sky130_fd_sc_hd__diode_2 ANTENNA__15918__A1 (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 ANTENNA__15919__A (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 ANTENNA__15928__A1 (.DIODE(net388));
 sky130_fd_sc_hd__diode_2 ANTENNA__15929__A1 (.DIODE(net378));
 sky130_fd_sc_hd__diode_2 ANTENNA__15929__A2 (.DIODE(net462));
 sky130_fd_sc_hd__diode_2 ANTENNA__15929__B2 (.DIODE(net384));
 sky130_fd_sc_hd__diode_2 ANTENNA__15931__A (.DIODE(net384));
 sky130_fd_sc_hd__diode_2 ANTENNA__15931__B (.DIODE(net378));
 sky130_fd_sc_hd__diode_2 ANTENNA__15931__C (.DIODE(net462));
 sky130_fd_sc_hd__diode_2 ANTENNA__15932__A1_N (.DIODE(net373));
 sky130_fd_sc_hd__diode_2 ANTENNA__15932__A2_N (.DIODE(net465));
 sky130_fd_sc_hd__diode_2 ANTENNA__15933__B (.DIODE(net465));
 sky130_fd_sc_hd__diode_2 ANTENNA__15933__C (.DIODE(net373));
 sky130_fd_sc_hd__diode_2 ANTENNA__15953__B1 (.DIODE(net331));
 sky130_fd_sc_hd__diode_2 ANTENNA__15953__B2 (.DIODE(net510));
 sky130_fd_sc_hd__diode_2 ANTENNA__15954__B (.DIODE(net510));
 sky130_fd_sc_hd__diode_2 ANTENNA__15954__C (.DIODE(net335));
 sky130_fd_sc_hd__diode_2 ANTENNA__15954__D (.DIODE(net331));
 sky130_fd_sc_hd__diode_2 ANTENNA__15956__A2 (.DIODE(\mul0.b[29] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15957__B (.DIODE(\mul0.b[29] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15961__A_N (.DIODE(net523));
 sky130_fd_sc_hd__diode_2 ANTENNA__15961__C (.DIODE(\mul0.b[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15963__A1_N (.DIODE(net519));
 sky130_fd_sc_hd__diode_2 ANTENNA__15963__B2 (.DIODE(net523));
 sky130_fd_sc_hd__diode_2 ANTENNA__15974__A2 (.DIODE(net347));
 sky130_fd_sc_hd__diode_2 ANTENNA__15974__B1 (.DIODE(net343));
 sky130_fd_sc_hd__diode_2 ANTENNA__15976__C (.DIODE(net347));
 sky130_fd_sc_hd__diode_2 ANTENNA__15976__D (.DIODE(net342));
 sky130_fd_sc_hd__diode_2 ANTENNA__15977__A2_N (.DIODE(net338));
 sky130_fd_sc_hd__diode_2 ANTENNA__15978__B (.DIODE(net338));
 sky130_fd_sc_hd__diode_2 ANTENNA__16024__A (.DIODE(_03057_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16025__A1 (.DIODE(net600));
 sky130_fd_sc_hd__diode_2 ANTENNA__16025__B1 (.DIODE(_02716_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16025__B2 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__16027__A (.DIODE(net388));
 sky130_fd_sc_hd__diode_2 ANTENNA__16030__A (.DIODE(_06985_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16031__A (.DIODE(_06985_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16036__A (.DIODE(_06983_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16037__A1 (.DIODE(_06983_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16037__B1_N (.DIODE(_06980_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16039__A1 (.DIODE(net354));
 sky130_fd_sc_hd__diode_2 ANTENNA__16039__B2 (.DIODE(net359));
 sky130_fd_sc_hd__diode_2 ANTENNA__16040__A (.DIODE(net359));
 sky130_fd_sc_hd__diode_2 ANTENNA__16040__B (.DIODE(net354));
 sky130_fd_sc_hd__diode_2 ANTENNA__16041__A2 (.DIODE(net351));
 sky130_fd_sc_hd__diode_2 ANTENNA__16042__B (.DIODE(net351));
 sky130_fd_sc_hd__diode_2 ANTENNA__16044__A1 (.DIODE(net368));
 sky130_fd_sc_hd__diode_2 ANTENNA__16044__A2 (.DIODE(net468));
 sky130_fd_sc_hd__diode_2 ANTENNA__16044__B1 (.DIODE(\mul0.a[27] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16044__B2 (.DIODE(net635));
 sky130_fd_sc_hd__diode_2 ANTENNA__16045__A (.DIODE(net635));
 sky130_fd_sc_hd__diode_2 ANTENNA__16045__B (.DIODE(net368));
 sky130_fd_sc_hd__diode_2 ANTENNA__16045__C (.DIODE(net468));
 sky130_fd_sc_hd__diode_2 ANTENNA__16045__D (.DIODE(net465));
 sky130_fd_sc_hd__diode_2 ANTENNA__16047__A1 (.DIODE(net363));
 sky130_fd_sc_hd__diode_2 ANTENNA__16048__A (.DIODE(net363));
 sky130_fd_sc_hd__diode_2 ANTENNA__16057__A1 (.DIODE(net388));
 sky130_fd_sc_hd__diode_2 ANTENNA__16058__A1 (.DIODE(net379));
 sky130_fd_sc_hd__diode_2 ANTENNA__16058__B2 (.DIODE(net385));
 sky130_fd_sc_hd__diode_2 ANTENNA__16059__A (.DIODE(net385));
 sky130_fd_sc_hd__diode_2 ANTENNA__16059__B (.DIODE(net379));
 sky130_fd_sc_hd__diode_2 ANTENNA__16061__A1 (.DIODE(net374));
 sky130_fd_sc_hd__diode_2 ANTENNA__16061__A2 (.DIODE(net462));
 sky130_fd_sc_hd__diode_2 ANTENNA__16062__B (.DIODE(net462));
 sky130_fd_sc_hd__diode_2 ANTENNA__16062__C (.DIODE(net374));
 sky130_fd_sc_hd__diode_2 ANTENNA__16083__A2 (.DIODE(net335));
 sky130_fd_sc_hd__diode_2 ANTENNA__16083__B1 (.DIODE(net332));
 sky130_fd_sc_hd__diode_2 ANTENNA__16084__C (.DIODE(net335));
 sky130_fd_sc_hd__diode_2 ANTENNA__16084__D (.DIODE(net332));
 sky130_fd_sc_hd__diode_2 ANTENNA__16086__A2 (.DIODE(net330));
 sky130_fd_sc_hd__diode_2 ANTENNA__16087__B (.DIODE(\mul0.b[29] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16092__A_N (.DIODE(net519));
 sky130_fd_sc_hd__diode_2 ANTENNA__16092__C (.DIODE(\mul0.b[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16093__B1 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__16093__B2 (.DIODE(net519));
 sky130_fd_sc_hd__diode_2 ANTENNA__16103__A2 (.DIODE(net347));
 sky130_fd_sc_hd__diode_2 ANTENNA__16103__B1 (.DIODE(net343));
 sky130_fd_sc_hd__diode_2 ANTENNA__16105__C (.DIODE(net347));
 sky130_fd_sc_hd__diode_2 ANTENNA__16105__D (.DIODE(net343));
 sky130_fd_sc_hd__diode_2 ANTENNA__16106__A2_N (.DIODE(\mul0.b[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16107__B (.DIODE(\mul0.b[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16119__A (.DIODE(_07575_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16121__B1 (.DIODE(_07575_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16145__A (.DIODE(_03057_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16146__A1 (.DIODE(net600));
 sky130_fd_sc_hd__diode_2 ANTENNA__16146__B1 (.DIODE(_02722_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16146__B2 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__16148__A1 (.DIODE(_06983_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16148__B1_N (.DIODE(_06980_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16153__A1 (.DIODE(net354));
 sky130_fd_sc_hd__diode_2 ANTENNA__16153__B1 (.DIODE(net471));
 sky130_fd_sc_hd__diode_2 ANTENNA__16153__B2 (.DIODE(net359));
 sky130_fd_sc_hd__diode_2 ANTENNA__16154__A (.DIODE(net359));
 sky130_fd_sc_hd__diode_2 ANTENNA__16154__B (.DIODE(net354));
 sky130_fd_sc_hd__diode_2 ANTENNA__16154__D (.DIODE(net471));
 sky130_fd_sc_hd__diode_2 ANTENNA__16156__A1 (.DIODE(net479));
 sky130_fd_sc_hd__diode_2 ANTENNA__16156__A2 (.DIODE(net351));
 sky130_fd_sc_hd__diode_2 ANTENNA__16157__A (.DIODE(net479));
 sky130_fd_sc_hd__diode_2 ANTENNA__16157__B (.DIODE(net351));
 sky130_fd_sc_hd__diode_2 ANTENNA__16159__A1 (.DIODE(net368));
 sky130_fd_sc_hd__diode_2 ANTENNA__16159__A2 (.DIODE(net465));
 sky130_fd_sc_hd__diode_2 ANTENNA__16159__B1 (.DIODE(\mul0.a[28] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16159__B2 (.DIODE(net635));
 sky130_fd_sc_hd__diode_2 ANTENNA__16160__A (.DIODE(net635));
 sky130_fd_sc_hd__diode_2 ANTENNA__16160__B (.DIODE(net368));
 sky130_fd_sc_hd__diode_2 ANTENNA__16160__C (.DIODE(\mul0.a[27] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16160__D (.DIODE(net462));
 sky130_fd_sc_hd__diode_2 ANTENNA__16162__A1 (.DIODE(net363));
 sky130_fd_sc_hd__diode_2 ANTENNA__16162__A2 (.DIODE(net469));
 sky130_fd_sc_hd__diode_2 ANTENNA__16163__A (.DIODE(net363));
 sky130_fd_sc_hd__diode_2 ANTENNA__16163__B (.DIODE(net468));
 sky130_fd_sc_hd__diode_2 ANTENNA__16173__A (.DIODE(net385));
 sky130_fd_sc_hd__diode_2 ANTENNA__16173__B (.DIODE(net453));
 sky130_fd_sc_hd__diode_2 ANTENNA__16174__A1 (.DIODE(net379));
 sky130_fd_sc_hd__diode_2 ANTENNA__16175__A (.DIODE(net379));
 sky130_fd_sc_hd__diode_2 ANTENNA__16177__A (.DIODE(net374));
 sky130_fd_sc_hd__diode_2 ANTENNA__16195__A2 (.DIODE(net336));
 sky130_fd_sc_hd__diode_2 ANTENNA__16195__B1 (.DIODE(net333));
 sky130_fd_sc_hd__diode_2 ANTENNA__16196__C (.DIODE(net336));
 sky130_fd_sc_hd__diode_2 ANTENNA__16196__D (.DIODE(net333));
 sky130_fd_sc_hd__diode_2 ANTENNA__16198__A1 (.DIODE(net506));
 sky130_fd_sc_hd__diode_2 ANTENNA__16198__A2 (.DIODE(net330));
 sky130_fd_sc_hd__diode_2 ANTENNA__16199__A (.DIODE(net506));
 sky130_fd_sc_hd__diode_2 ANTENNA__16199__B (.DIODE(net330));
 sky130_fd_sc_hd__diode_2 ANTENNA__16203__A_N (.DIODE(net514));
 sky130_fd_sc_hd__diode_2 ANTENNA__16203__B (.DIODE(net328));
 sky130_fd_sc_hd__diode_2 ANTENNA__16203__C (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA__16203__D (.DIODE(net510));
 sky130_fd_sc_hd__diode_2 ANTENNA__16204__A1_N (.DIODE(net510));
 sky130_fd_sc_hd__diode_2 ANTENNA__16204__A2_N (.DIODE(net328));
 sky130_fd_sc_hd__diode_2 ANTENNA__16204__B1 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__16204__B2 (.DIODE(net514));
 sky130_fd_sc_hd__diode_2 ANTENNA__16214__A1 (.DIODE(net484));
 sky130_fd_sc_hd__diode_2 ANTENNA__16214__A2 (.DIODE(net347));
 sky130_fd_sc_hd__diode_2 ANTENNA__16214__B1 (.DIODE(net343));
 sky130_fd_sc_hd__diode_2 ANTENNA__16214__B2 (.DIODE(net488));
 sky130_fd_sc_hd__diode_2 ANTENNA__16215__A (.DIODE(net488));
 sky130_fd_sc_hd__diode_2 ANTENNA__16215__B (.DIODE(net484));
 sky130_fd_sc_hd__diode_2 ANTENNA__16215__C (.DIODE(net347));
 sky130_fd_sc_hd__diode_2 ANTENNA__16215__D (.DIODE(net343));
 sky130_fd_sc_hd__diode_2 ANTENNA__16217__A1 (.DIODE(net493));
 sky130_fd_sc_hd__diode_2 ANTENNA__16217__A2 (.DIODE(\mul0.b[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16218__A (.DIODE(net493));
 sky130_fd_sc_hd__diode_2 ANTENNA__16218__B (.DIODE(net337));
 sky130_fd_sc_hd__diode_2 ANTENNA__16232__A (.DIODE(_07685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16233__B1 (.DIODE(_07685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16257__A (.DIODE(_03057_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16258__A1 (.DIODE(net600));
 sky130_fd_sc_hd__diode_2 ANTENNA__16258__B1 (.DIODE(_02727_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16258__B2 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__16262__A1 (.DIODE(_06980_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16265__A1 (.DIODE(net354));
 sky130_fd_sc_hd__diode_2 ANTENNA__16265__A2 (.DIODE(net471));
 sky130_fd_sc_hd__diode_2 ANTENNA__16265__B1 (.DIODE(net468));
 sky130_fd_sc_hd__diode_2 ANTENNA__16265__B2 (.DIODE(net359));
 sky130_fd_sc_hd__diode_2 ANTENNA__16266__A (.DIODE(net359));
 sky130_fd_sc_hd__diode_2 ANTENNA__16266__B (.DIODE(net354));
 sky130_fd_sc_hd__diode_2 ANTENNA__16266__C (.DIODE(net471));
 sky130_fd_sc_hd__diode_2 ANTENNA__16267__A1 (.DIODE(net468));
 sky130_fd_sc_hd__diode_2 ANTENNA__16268__A (.DIODE(net351));
 sky130_fd_sc_hd__diode_2 ANTENNA__16270__A1 (.DIODE(net368));
 sky130_fd_sc_hd__diode_2 ANTENNA__16270__A2 (.DIODE(net462));
 sky130_fd_sc_hd__diode_2 ANTENNA__16270__B1 (.DIODE(\mul0.a[29] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16270__B2 (.DIODE(net635));
 sky130_fd_sc_hd__diode_2 ANTENNA__16271__A (.DIODE(net635));
 sky130_fd_sc_hd__diode_2 ANTENNA__16271__B (.DIODE(net368));
 sky130_fd_sc_hd__diode_2 ANTENNA__16271__C (.DIODE(net462));
 sky130_fd_sc_hd__diode_2 ANTENNA__16273__A (.DIODE(net363));
 sky130_fd_sc_hd__diode_2 ANTENNA__16273__B (.DIODE(net465));
 sky130_fd_sc_hd__diode_2 ANTENNA__16282__A1 (.DIODE(net385));
 sky130_fd_sc_hd__diode_2 ANTENNA__16282__A2 (.DIODE(net379));
 sky130_fd_sc_hd__diode_2 ANTENNA__16284__A (.DIODE(net379));
 sky130_fd_sc_hd__diode_2 ANTENNA__16285__A1 (.DIODE(net374));
 sky130_fd_sc_hd__diode_2 ANTENNA__16286__A (.DIODE(net374));
 sky130_fd_sc_hd__diode_2 ANTENNA__16304__A2 (.DIODE(net336));
 sky130_fd_sc_hd__diode_2 ANTENNA__16304__B1 (.DIODE(net333));
 sky130_fd_sc_hd__diode_2 ANTENNA__16304__B2 (.DIODE(net497));
 sky130_fd_sc_hd__diode_2 ANTENNA__16305__A (.DIODE(net497));
 sky130_fd_sc_hd__diode_2 ANTENNA__16305__C (.DIODE(net336));
 sky130_fd_sc_hd__diode_2 ANTENNA__16305__D (.DIODE(net333));
 sky130_fd_sc_hd__diode_2 ANTENNA__16307__B (.DIODE(net330));
 sky130_fd_sc_hd__diode_2 ANTENNA__16313__A1 (.DIODE(net506));
 sky130_fd_sc_hd__diode_2 ANTENNA__16313__A2 (.DIODE(net328));
 sky130_fd_sc_hd__diode_2 ANTENNA__16313__B1 (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA__16314__A (.DIODE(net506));
 sky130_fd_sc_hd__diode_2 ANTENNA__16314__C (.DIODE(net328));
 sky130_fd_sc_hd__diode_2 ANTENNA__16314__D (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA__16325__A1 (.DIODE(net479));
 sky130_fd_sc_hd__diode_2 ANTENNA__16325__A2 (.DIODE(net347));
 sky130_fd_sc_hd__diode_2 ANTENNA__16325__B1 (.DIODE(net343));
 sky130_fd_sc_hd__diode_2 ANTENNA__16325__B2 (.DIODE(net484));
 sky130_fd_sc_hd__diode_2 ANTENNA__16326__A (.DIODE(net484));
 sky130_fd_sc_hd__diode_2 ANTENNA__16326__B (.DIODE(net479));
 sky130_fd_sc_hd__diode_2 ANTENNA__16326__C (.DIODE(net347));
 sky130_fd_sc_hd__diode_2 ANTENNA__16326__D (.DIODE(net343));
 sky130_fd_sc_hd__diode_2 ANTENNA__16328__A (.DIODE(net488));
 sky130_fd_sc_hd__diode_2 ANTENNA__16328__B (.DIODE(net337));
 sky130_fd_sc_hd__diode_2 ANTENNA__16358__A (.DIODE(_07829_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16359__A (.DIODE(_07829_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16363__A (.DIODE(net600));
 sky130_fd_sc_hd__diode_2 ANTENNA__16364__A1 (.DIODE(_02732_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16364__A2 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__16364__B2 (.DIODE(_03058_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16369__A (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 ANTENNA__16369__B (.DIODE(net462));
 sky130_fd_sc_hd__diode_2 ANTENNA__16371__A (.DIODE(net368));
 sky130_fd_sc_hd__diode_2 ANTENNA__16371__B (.DIODE(\mul0.a[29] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16374__A (.DIODE(net506));
 sky130_fd_sc_hd__diode_2 ANTENNA__16374__B (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__16377__A (.DIODE(net351));
 sky130_fd_sc_hd__diode_2 ANTENNA__16380__A (.DIODE(net635));
 sky130_fd_sc_hd__diode_2 ANTENNA__16380__B (.DIODE(net456));
 sky130_fd_sc_hd__diode_2 ANTENNA__16386__A1 (.DIODE(net363));
 sky130_fd_sc_hd__diode_2 ANTENNA__16386__A2 (.DIODE(net465));
 sky130_fd_sc_hd__diode_2 ANTENNA__16387__A (.DIODE(_07857_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16391__A (.DIODE(net359));
 sky130_fd_sc_hd__diode_2 ANTENNA__16391__B (.DIODE(net465));
 sky130_fd_sc_hd__diode_2 ANTENNA__16396__B (.DIODE(net347));
 sky130_fd_sc_hd__diode_2 ANTENNA__16399__B (.DIODE(net336));
 sky130_fd_sc_hd__diode_2 ANTENNA__16401__A1 (.DIODE(net351));
 sky130_fd_sc_hd__diode_2 ANTENNA__16401__B2 (.DIODE(net468));
 sky130_fd_sc_hd__diode_2 ANTENNA__16402__A2 (.DIODE(net330));
 sky130_fd_sc_hd__diode_2 ANTENNA__16404__A (.DIODE(net497));
 sky130_fd_sc_hd__diode_2 ANTENNA__16404__B (.DIODE(net330));
 sky130_fd_sc_hd__diode_2 ANTENNA__16406__B (.DIODE(net328));
 sky130_fd_sc_hd__diode_2 ANTENNA__16409__A (.DIODE(net493));
 sky130_fd_sc_hd__diode_2 ANTENNA__16409__B (.DIODE(net333));
 sky130_fd_sc_hd__diode_2 ANTENNA__16414__A (.DIODE(net354));
 sky130_fd_sc_hd__diode_2 ANTENNA__16414__B (.DIODE(net468));
 sky130_fd_sc_hd__diode_2 ANTENNA__16415__B1 (.DIODE(_06980_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16417__A1 (.DIODE(net488));
 sky130_fd_sc_hd__diode_2 ANTENNA__16417__A2 (.DIODE(\mul0.b[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16418__A (.DIODE(net479));
 sky130_fd_sc_hd__diode_2 ANTENNA__16418__B (.DIODE(net343));
 sky130_fd_sc_hd__diode_2 ANTENNA__16424__B (.DIODE(\mul0.b[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16427__D1 (.DIODE(net374));
 sky130_fd_sc_hd__diode_2 ANTENNA__16428__A1 (.DIODE(net385));
 sky130_fd_sc_hd__diode_2 ANTENNA__16428__A2 (.DIODE(net379));
 sky130_fd_sc_hd__diode_2 ANTENNA__16437__B (.DIODE(_07908_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16438__A1 (.DIODE(net600));
 sky130_fd_sc_hd__diode_2 ANTENNA__16438__B1 (.DIODE(_03058_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16439__A1 (.DIODE(_02735_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16439__A2 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__16441__B (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__16441__C (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__16441__D (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA__16442__A2 (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__16442__B1 (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA__16442__B2 (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__16443__C (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__16443__D (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA__16445__A (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__16445__B (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA__16446__A1 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__16446__A2 (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA__16446__B2 (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA__16447__A (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__16447__B (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA__16448__A1 (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA__16451__A (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__16451__B (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA__16451__D (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA__16452__A (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__16452__B (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA__16453__A1 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__16453__B1 (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA__16453__B2 (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA__16455__A1 (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__16455__A2 (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 ANTENNA__16458__A (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__16458__B (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA__16459__A2 (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA__16459__B1 (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA__16460__C (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA__16461__A1 (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA__16463__C (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA__16463__D (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA__16464__A (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__16464__B (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA__16465__A2 (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA__16465__B1 (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA__16467__A1 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__16467__A2 (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA__16469__A1 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__16469__A2 (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA__16469__B1 (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA__16469__B2 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__16470__A (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__16470__B (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__16470__C (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA__16470__D (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA__16472__A (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__16473__A1 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__16473__A2 (.DIODE(net320));
 sky130_fd_sc_hd__diode_2 ANTENNA__16479__C (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA__16479__D (.DIODE(net309));
 sky130_fd_sc_hd__diode_2 ANTENNA__16480__A (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__16480__B (.DIODE(net314));
 sky130_fd_sc_hd__diode_2 ANTENNA__16481__A2 (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA__16481__B1 (.DIODE(net309));
 sky130_fd_sc_hd__diode_2 ANTENNA__16483__A1 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__16483__A2 (.DIODE(net314));
 sky130_fd_sc_hd__diode_2 ANTENNA__16486__A1 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__16486__A2 (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA__16486__B2 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__16487__A (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__16487__B (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__16487__C (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA__16489__A (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__16489__B (.DIODE(net323));
 sky130_fd_sc_hd__diode_2 ANTENNA__16490__A1 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__16490__A2 (.DIODE(net323));
 sky130_fd_sc_hd__diode_2 ANTENNA__16496__A (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__16496__B (.DIODE(net323));
 sky130_fd_sc_hd__diode_2 ANTENNA__16498__A2 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__16498__B1 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__16498__B2 (.DIODE(net323));
 sky130_fd_sc_hd__diode_2 ANTENNA__16499__B (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__16499__C (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__16499__D (.DIODE(net323));
 sky130_fd_sc_hd__diode_2 ANTENNA__16500__A (.DIODE(net320));
 sky130_fd_sc_hd__diode_2 ANTENNA__16500__B (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__16500__C (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__16500__D (.DIODE(net323));
 sky130_fd_sc_hd__diode_2 ANTENNA__16507__A (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__16507__B (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__16507__C (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA__16507__D (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__16508__A1 (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__16508__A2 (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA__16508__B1 (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__16508__B2 (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__16509__C (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__16509__D (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA__16510__A1 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__16510__A2 (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA__16510__B1 (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA__16510__B2 (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA__16511__A (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__16511__B (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA__16511__C (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA__16511__D (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA__16512__A (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__16512__B (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA__16513__A1 (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__16513__A2 (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA__16515__A1 (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__16515__A2 (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA__16515__B2 (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA__16519__A (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__16519__B (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA__16520__A1 (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA__16520__B2 (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA__16521__A (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA__16521__D (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA__16524__A1 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__16524__A2 (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 ANTENNA__16524__B2 (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA__16527__A (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__16527__B (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA__16528__A1 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__16528__A2 (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 ANTENNA__16528__B1 (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA__16528__B2 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__16529__A (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__16529__B (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__16529__C (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 ANTENNA__16529__D (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA__16539__A1 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__16539__A2 (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA__16540__A (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__16540__B (.DIODE(net323));
 sky130_fd_sc_hd__diode_2 ANTENNA__16541__A (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA__16541__C (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__16541__D (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__16542__A1 (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA__16542__A2 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__16542__B1 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__16554__A (.DIODE(\mul1.b[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16554__B (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__16554__C (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA__16554__D (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA__16555__A (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__16555__B (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__16556__A1 (.DIODE(\mul1.b[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16556__A2 (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA__16556__B1 (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA__16556__B2 (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__16558__A1 (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__16558__A2 (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__16559__A1 (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__16559__A2 (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__16559__B1 (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA__16559__B2 (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA__16560__A (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__16560__B (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA__16560__C (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__16560__D (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA__16561__A (.DIODE(\mul1.b[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16561__B (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA__16562__A1 (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__16562__A2 (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA__16568__A (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__16568__B (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA__16569__A (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA__16569__B (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__16569__C (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__16569__D (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 ANTENNA__16570__A1 (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA__16570__A2 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__16570__B1 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__16570__B2 (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 ANTENNA__16573__A (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA__16573__B (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA__16574__A1 (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA__16574__B2 (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA__16575__A (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__16575__B (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA__16576__A1 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__16576__A2 (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA__16587__A (.DIODE(\mul1.b[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16587__B (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__16587__C (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__16587__D (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA__16588__A1 (.DIODE(\mul1.b[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16588__A2 (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__16588__B1 (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA__16588__B2 (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__16589__C (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__16589__D (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA__16591__A (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__16591__B (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA__16592__A (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA__16592__B (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__16592__C (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA__16592__D (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 ANTENNA__16593__A1 (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA__16593__A2 (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__16593__B1 (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA__16593__B2 (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 ANTENNA__16600__A (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__16600__B (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA__16601__A1 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__16601__A2 (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__16601__B1 (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__16601__B2 (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__16602__A (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__16602__B (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__16602__C (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__16602__D (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__16605__A (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__16605__B (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__16606__A (.DIODE(net625));
 sky130_fd_sc_hd__diode_2 ANTENNA__16606__B (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__16606__C (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__16606__D (.DIODE(net630));
 sky130_fd_sc_hd__diode_2 ANTENNA__16607__A1 (.DIODE(net625));
 sky130_fd_sc_hd__diode_2 ANTENNA__16607__A2 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__16607__B1 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__16607__B2 (.DIODE(net630));
 sky130_fd_sc_hd__diode_2 ANTENNA__16610__A (.DIODE(\mul1.b[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16610__B (.DIODE(\mul1.b[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16610__C (.DIODE(net630));
 sky130_fd_sc_hd__diode_2 ANTENNA__16610__D (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__16611__A (.DIODE(\mul1.b[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16611__B (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__16612__A1 (.DIODE(\mul1.b[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16612__A2 (.DIODE(net630));
 sky130_fd_sc_hd__diode_2 ANTENNA__16612__B1 (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__16612__B2 (.DIODE(\mul1.b[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16619__A (.DIODE(net622));
 sky130_fd_sc_hd__diode_2 ANTENNA__16619__B (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__16619__C (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__16619__D (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__16620__A (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__16620__B (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__16621__A1 (.DIODE(net622));
 sky130_fd_sc_hd__diode_2 ANTENNA__16621__A2 (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__16621__B1 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__16621__B2 (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__16627__A1_N (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__16627__A2_N (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA__16636__A (.DIODE(net622));
 sky130_fd_sc_hd__diode_2 ANTENNA__16636__B (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__16636__C (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__16636__D (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__16637__A (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__16637__B (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA__16638__A1 (.DIODE(net622));
 sky130_fd_sc_hd__diode_2 ANTENNA__16638__A2 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__16638__B1 (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__16638__B2 (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__16659__C (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__16659__D (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA__16660__A (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__16660__B (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA__16661__A2 (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__16661__B1 (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA__16667__A1_N (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__16667__A2_N (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA__16688__C (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA__16688__D (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA__16689__A (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__16689__B (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__16690__A2 (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA__16690__B1 (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA__16696__A1_N (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__16696__A2_N (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA__16724__B (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__16724__C (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA__16724__D (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__16725__A (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__16725__B (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA__16726__A1 (.DIODE(net622));
 sky130_fd_sc_hd__diode_2 ANTENNA__16726__A2 (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA__16726__B1 (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__16726__B2 (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__16732__A (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__16733__B (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__16733__C (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA__16734__B (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__16734__C (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA__16734__D (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA__16735__A2 (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA__16735__B1 (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA__16735__B2 (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__16743__A (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__16743__B (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA__16743__C (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA__16743__D (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA__16744__A (.DIODE(\mul1.b[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16744__B (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA__16745__A1 (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__16745__A2 (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA__16745__B1 (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA__16745__B2 (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA__16747__A1 (.DIODE(\mul1.b[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16747__A2 (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA__16748__A1 (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__16759__C (.DIODE(net309));
 sky130_fd_sc_hd__diode_2 ANTENNA__16759__D (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA__16760__A (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__16761__A2 (.DIODE(net309));
 sky130_fd_sc_hd__diode_2 ANTENNA__16761__B1 (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA__16763__A1 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__16766__A1 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__16766__B1 (.DIODE(net323));
 sky130_fd_sc_hd__diode_2 ANTENNA__16766__B2 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__16768__A (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__16768__B (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__16768__D (.DIODE(net323));
 sky130_fd_sc_hd__diode_2 ANTENNA__16794__C (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__16794__D (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA__16795__A (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__16795__B (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA__16796__A2 (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__16796__B1 (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA__16802__A (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__16802__B (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA__16803__A2 (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA__16803__B2 (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__16812__A (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__16812__B (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA__16812__C (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 ANTENNA__16812__D (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA__16813__A (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__16813__B (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA__16813__C (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 ANTENNA__16813__D (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA__16814__A1 (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__16814__A2 (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 ANTENNA__16814__B1 (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA__16814__B2 (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA__16815__A (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__16815__B (.DIODE(net309));
 sky130_fd_sc_hd__diode_2 ANTENNA__16817__A1 (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__16817__A2 (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA__16829__C (.DIODE(net314));
 sky130_fd_sc_hd__diode_2 ANTENNA__16829__D (.DIODE(net320));
 sky130_fd_sc_hd__diode_2 ANTENNA__16831__A2 (.DIODE(net314));
 sky130_fd_sc_hd__diode_2 ANTENNA__16831__B1 (.DIODE(net320));
 sky130_fd_sc_hd__diode_2 ANTENNA__16832__C (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__16832__D (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA__16835__A (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__16835__B (.DIODE(net323));
 sky130_fd_sc_hd__diode_2 ANTENNA__16860__C (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA__16860__D (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA__16861__A (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__16862__A2 (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA__16862__B1 (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA__16867__A1 (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__16867__B1 (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA__16867__B2 (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__16868__B (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__16869__A1 (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA__16870__A (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__16870__B (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA__16877__A1 (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__16877__A2 (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA__16877__B2 (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA__16878__A1 (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__16878__A2 (.DIODE(net309));
 sky130_fd_sc_hd__diode_2 ANTENNA__16882__A (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__16882__B (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA__16882__C (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA__16883__A (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__16883__B (.DIODE(net313));
 sky130_fd_sc_hd__diode_2 ANTENNA__16884__A1 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__16884__A2 (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA__16884__B1 (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA__16884__B2 (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA__16885__A1 (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA__16886__A1_N (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA__16897__A1 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__16897__A2 (.DIODE(net325));
 sky130_fd_sc_hd__diode_2 ANTENNA__16899__C (.DIODE(net320));
 sky130_fd_sc_hd__diode_2 ANTENNA__16899__D (.DIODE(net325));
 sky130_fd_sc_hd__diode_2 ANTENNA__16917__C (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA__16918__A (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__16918__B (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA__16919__A2 (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA__16924__A1 (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__16924__A2 (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA__16924__B1 (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA__16924__B2 (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__16925__A (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__16925__B (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__16925__C (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA__16925__D (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA__16927__A (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__16927__B (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA__16938__A (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__16938__B (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA__16938__C (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA__16938__D (.DIODE(net313));
 sky130_fd_sc_hd__diode_2 ANTENNA__16939__A (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__16939__B (.DIODE(net318));
 sky130_fd_sc_hd__diode_2 ANTENNA__16940__A1 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__16940__A2 (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA__16940__B1 (.DIODE(net313));
 sky130_fd_sc_hd__diode_2 ANTENNA__16940__B2 (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA__16942__A1 (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__16942__A2 (.DIODE(net318));
 sky130_fd_sc_hd__diode_2 ANTENNA__16968__D (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA__16969__A (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__16969__B (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA__16970__B1 (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA__16974__A1 (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__16974__A2 (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA__16974__B1 (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA__16974__B2 (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__16975__A (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__16975__B (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__16975__C (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA__16975__D (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA__16976__A1_N (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__16976__A2_N (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA__16977__C (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__16977__D (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA__16987__A (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__16987__B (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA__16987__C (.DIODE(net313));
 sky130_fd_sc_hd__diode_2 ANTENNA__16987__D (.DIODE(net318));
 sky130_fd_sc_hd__diode_2 ANTENNA__16988__A1 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__16988__A2 (.DIODE(net313));
 sky130_fd_sc_hd__diode_2 ANTENNA__16988__B1 (.DIODE(net318));
 sky130_fd_sc_hd__diode_2 ANTENNA__16988__B2 (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA__16989__C (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__16989__D (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA__16996__A2 (.DIODE(net320));
 sky130_fd_sc_hd__diode_2 ANTENNA__16996__B1 (.DIODE(net325));
 sky130_fd_sc_hd__diode_2 ANTENNA__17013__A (.DIODE(net622));
 sky130_fd_sc_hd__diode_2 ANTENNA__17013__C (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA__17013__D (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA__17014__A (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__17014__B (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA__17015__A2 (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA__17015__B1 (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA__17019__A (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__17019__B (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__17019__C (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA__17019__D (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA__17020__A1 (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__17020__A2 (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA__17020__B1 (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA__17020__B2 (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__17022__A (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__17022__B (.DIODE(net313));
 sky130_fd_sc_hd__diode_2 ANTENNA__17029__A (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__17029__B (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA__17029__C (.DIODE(net318));
 sky130_fd_sc_hd__diode_2 ANTENNA__17029__D (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA__17031__A1 (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__17031__A2 (.DIODE(net313));
 sky130_fd_sc_hd__diode_2 ANTENNA__17032__A1_N (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__17032__A2_N (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA__17041__B (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA__17052__A (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__17052__B (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__17052__C (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA__17052__D (.DIODE(net313));
 sky130_fd_sc_hd__diode_2 ANTENNA__17053__A1 (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__17053__A2 (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA__17053__B1 (.DIODE(net313));
 sky130_fd_sc_hd__diode_2 ANTENNA__17053__B2 (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__17055__A (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__17055__B (.DIODE(net318));
 sky130_fd_sc_hd__diode_2 ANTENNA__17056__A1 (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__17056__A2 (.DIODE(net318));
 sky130_fd_sc_hd__diode_2 ANTENNA__17057__A1 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__17057__A2 (.DIODE(net318));
 sky130_fd_sc_hd__diode_2 ANTENNA__17057__B1 (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA__17057__B2 (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA__17063__A (.DIODE(net622));
 sky130_fd_sc_hd__diode_2 ANTENNA__17063__B (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__17063__C (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 ANTENNA__17063__D (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA__17064__A (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__17064__B (.DIODE(net309));
 sky130_fd_sc_hd__diode_2 ANTENNA__17065__A1 (.DIODE(net622));
 sky130_fd_sc_hd__diode_2 ANTENNA__17065__A2 (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 ANTENNA__17065__B1 (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA__17065__B2 (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__17086__A (.DIODE(net622));
 sky130_fd_sc_hd__diode_2 ANTENNA__17086__B (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__17086__C (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA__17086__D (.DIODE(net309));
 sky130_fd_sc_hd__diode_2 ANTENNA__17087__A (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__17087__B (.DIODE(net313));
 sky130_fd_sc_hd__diode_2 ANTENNA__17088__A1 (.DIODE(net622));
 sky130_fd_sc_hd__diode_2 ANTENNA__17088__A2 (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA__17088__B1 (.DIODE(net309));
 sky130_fd_sc_hd__diode_2 ANTENNA__17088__B2 (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__17092__A1 (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__17092__A2 (.DIODE(net313));
 sky130_fd_sc_hd__diode_2 ANTENNA__17092__B1 (.DIODE(net318));
 sky130_fd_sc_hd__diode_2 ANTENNA__17092__B2 (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__17093__A (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__17093__B (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__17093__C (.DIODE(net313));
 sky130_fd_sc_hd__diode_2 ANTENNA__17093__D (.DIODE(net318));
 sky130_fd_sc_hd__diode_2 ANTENNA__17095__A (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__17095__B (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA__17096__A (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__17096__B (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA__17102__B1 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__17102__C1 (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA__17103__A1 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__17103__A2 (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA__17123__A (.DIODE(net622));
 sky130_fd_sc_hd__diode_2 ANTENNA__17123__B (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__17123__C (.DIODE(net309));
 sky130_fd_sc_hd__diode_2 ANTENNA__17123__D (.DIODE(net313));
 sky130_fd_sc_hd__diode_2 ANTENNA__17124__A (.DIODE(net622));
 sky130_fd_sc_hd__diode_2 ANTENNA__17124__B (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__17124__C (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA__17124__D (.DIODE(net314));
 sky130_fd_sc_hd__diode_2 ANTENNA__17125__A1 (.DIODE(net622));
 sky130_fd_sc_hd__diode_2 ANTENNA__17125__A2 (.DIODE(net309));
 sky130_fd_sc_hd__diode_2 ANTENNA__17125__B1 (.DIODE(net314));
 sky130_fd_sc_hd__diode_2 ANTENNA__17125__B2 (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__17126__A (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__17126__B (.DIODE(net320));
 sky130_fd_sc_hd__diode_2 ANTENNA__17128__A1 (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__17128__A2 (.DIODE(net318));
 sky130_fd_sc_hd__diode_2 ANTENNA__17128__B1 (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA__17128__B2 (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__17129__A (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__17129__B (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__17129__C (.DIODE(net318));
 sky130_fd_sc_hd__diode_2 ANTENNA__17129__D (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA__17139__A1 (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__17139__A2 (.DIODE(net318));
 sky130_fd_sc_hd__diode_2 ANTENNA__17141__C (.DIODE(net314));
 sky130_fd_sc_hd__diode_2 ANTENNA__17141__D (.DIODE(net320));
 sky130_fd_sc_hd__diode_2 ANTENNA__17142__A2 (.DIODE(net313));
 sky130_fd_sc_hd__diode_2 ANTENNA__17142__B1 (.DIODE(net318));
 sky130_fd_sc_hd__diode_2 ANTENNA__17143__A1 (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__17143__A2 (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA__17144__A (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__17144__B (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA__17145__A (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__17145__B (.DIODE(net313));
 sky130_fd_sc_hd__diode_2 ANTENNA__17146__A (.DIODE(net622));
 sky130_fd_sc_hd__diode_2 ANTENNA__17146__B (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__17146__C (.DIODE(net318));
 sky130_fd_sc_hd__diode_2 ANTENNA__17146__D (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA__17172__A (.DIODE(_03049_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17172__B (.DIODE(_08642_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17173__A (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__17173__B (.DIODE(_03792_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17174__A2 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__17174__B1 (.DIODE(_03056_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17179__A1 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__17179__A2 (.DIODE(net323));
 sky130_fd_sc_hd__diode_2 ANTENNA__17180__A1 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__17180__A2 (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA__17181__A (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA__17181__B (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA__17181__C (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__17181__D (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__17182__A1 (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA__17182__A2 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__17182__B1 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__17182__B2 (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA__17183__B (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__17184__A2 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__17192__A (.DIODE(net323));
 sky130_fd_sc_hd__diode_2 ANTENNA__17192__B (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__17193__A (.DIODE(net323));
 sky130_fd_sc_hd__diode_2 ANTENNA__17193__B (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__17200__A (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA__17200__B (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA__17200__C (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__17200__D (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__17202__A1 (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA__17202__A2 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__17202__B1 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__17202__B2 (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA__17203__C (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 ANTENNA__17203__D (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__17204__A1 (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 ANTENNA__17204__A2 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__17206__A (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA__17206__B (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__17207__A (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA__17207__B (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA__17208__A1 (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA__17208__B2 (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA__17221__A1 (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__17221__A2 (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA__17223__A (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__17223__B (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__17224__A (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA__17224__B (.DIODE(net272));
 sky130_fd_sc_hd__diode_2 ANTENNA__17224__C (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__17224__D (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__17225__A1 (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA__17225__A2 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__17225__B1 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__17225__B2 (.DIODE(net272));
 sky130_fd_sc_hd__diode_2 ANTENNA__17232__A (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__17232__B (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__17233__A1 (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__17233__A2 (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__17233__B1 (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__17233__B2 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__17234__A (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__17234__B (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__17234__C (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__17234__D (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__17237__A (.DIODE(net630));
 sky130_fd_sc_hd__diode_2 ANTENNA__17237__B (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__17238__A (.DIODE(net625));
 sky130_fd_sc_hd__diode_2 ANTENNA__17238__B (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__17238__C (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__17238__D (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA__17239__A1 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__17239__A2 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__17239__B1 (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA__17239__B2 (.DIODE(net625));
 sky130_fd_sc_hd__diode_2 ANTENNA__17272__A1 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__17272__A2 (.DIODE(_03893_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17272__B1 (.DIODE(_08741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17272__B2 (.DIODE(_03049_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17273__A2 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__17276__A2 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__17276__B1 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__17276__B2 (.DIODE(net323));
 sky130_fd_sc_hd__diode_2 ANTENNA__17277__B (.DIODE(net323));
 sky130_fd_sc_hd__diode_2 ANTENNA__17277__C (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__17277__D (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__17280__A1 (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA__17280__A2 (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA__17280__A3 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__17280__A4 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__17282__A (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA__17282__B (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__17283__A (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 ANTENNA__17283__B (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA__17283__C (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__17283__D (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__17284__A1 (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 ANTENNA__17284__A2 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__17284__B1 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__17284__B2 (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA__17300__A (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA__17300__B (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA__17300__C (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__17300__D (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__17302__A1 (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA__17302__A2 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__17302__B1 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__17302__B2 (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA__17303__C (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA__17303__D (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__17304__A1 (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA__17304__A2 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__17306__A (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA__17306__B (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__17307__A (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 ANTENNA__17307__B (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA__17308__A1 (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 ANTENNA__17308__B2 (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA__17311__A1 (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA__17311__A2 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__17321__A1 (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__17321__A2 (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__17323__A (.DIODE(net272));
 sky130_fd_sc_hd__diode_2 ANTENNA__17323__B (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__17324__A (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__17324__B (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA__17324__C (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__17324__D (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__17325__A1 (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__17325__A2 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__17325__B1 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__17325__B2 (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA__17332__A (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__17332__B (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__17333__A1 (.DIODE(net630));
 sky130_fd_sc_hd__diode_2 ANTENNA__17333__A2 (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__17333__B1 (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__17333__B2 (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__17334__A (.DIODE(net630));
 sky130_fd_sc_hd__diode_2 ANTENNA__17334__B (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__17334__C (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__17334__D (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__17337__A (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__17337__B (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__17338__A (.DIODE(net625));
 sky130_fd_sc_hd__diode_2 ANTENNA__17338__B (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__17338__C (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA__17338__D (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA__17339__A1 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__17339__A2 (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA__17339__B1 (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA__17339__B2 (.DIODE(net625));
 sky130_fd_sc_hd__diode_2 ANTENNA__17375__A1 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__17375__A2 (.DIODE(_03993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17375__B1 (.DIODE(_08843_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17375__B2 (.DIODE(_03049_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17376__A2 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__17378__A (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__17378__B (.DIODE(_04100_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17384__A (.DIODE(\mul1.a[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17384__B (.DIODE(net320));
 sky130_fd_sc_hd__diode_2 ANTENNA__17384__C (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__17384__D (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__17385__A1 (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA__17385__A2 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__17385__B1 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__17387__A (.DIODE(net323));
 sky130_fd_sc_hd__diode_2 ANTENNA__17387__B (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__17392__A1 (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA__17392__A2 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__17394__A (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA__17394__B (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__17395__A (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA__17395__B (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 ANTENNA__17395__C (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__17395__D (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__17396__A1 (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA__17396__A2 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__17396__B1 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__17396__B2 (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 ANTENNA__17411__A (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA__17411__B (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA__17411__C (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__17411__D (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__17412__A1 (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA__17412__A2 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__17412__B1 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__17412__B2 (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA__17413__A (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA__17413__B (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__17414__A1 (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA__17414__A2 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__17416__A (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA__17416__B (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__17417__A (.DIODE(net272));
 sky130_fd_sc_hd__diode_2 ANTENNA__17417__B (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 ANTENNA__17418__A1 (.DIODE(net272));
 sky130_fd_sc_hd__diode_2 ANTENNA__17418__B2 (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 ANTENNA__17421__A1 (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA__17421__A2 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__17431__A1 (.DIODE(net272));
 sky130_fd_sc_hd__diode_2 ANTENNA__17431__A2 (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__17433__A (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA__17433__B (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__17434__A (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__17434__B (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__17434__C (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__17434__D (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA__17435__A1 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__17435__A2 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__17435__B1 (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA__17435__B2 (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__17442__A (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__17442__B (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__17443__A (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__17443__B (.DIODE(net630));
 sky130_fd_sc_hd__diode_2 ANTENNA__17443__C (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__17443__D (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__17444__A1 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__17444__B1 (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__17444__B2 (.DIODE(net630));
 sky130_fd_sc_hd__diode_2 ANTENNA__17447__A (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__17447__B (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA__17448__A (.DIODE(net625));
 sky130_fd_sc_hd__diode_2 ANTENNA__17448__B (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__17448__C (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA__17448__D (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA__17449__A1 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__17449__A2 (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA__17449__B1 (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA__17449__B2 (.DIODE(net625));
 sky130_fd_sc_hd__diode_2 ANTENNA__17485__A2 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__17485__B1 (.DIODE(_08952_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17485__B2 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__17490__A (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA__17490__B (.DIODE(\mul1.a[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17490__C (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__17490__D (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__17492__A1 (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA__17492__A2 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__17492__B1 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__17492__B2 (.DIODE(\mul1.a[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17493__A (.DIODE(net320));
 sky130_fd_sc_hd__diode_2 ANTENNA__17493__B (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__17494__A1 (.DIODE(net320));
 sky130_fd_sc_hd__diode_2 ANTENNA__17494__A2 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__17499__A (.DIODE(net325));
 sky130_fd_sc_hd__diode_2 ANTENNA__17499__B (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__17501__A1 (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA__17501__A2 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__17502__A (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA__17502__B (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA__17502__C (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__17502__D (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__17503__A1 (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA__17503__A2 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__17503__B1 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__17503__B2 (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA__17504__C (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 ANTENNA__17504__D (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__17505__A1_N (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 ANTENNA__17505__A2_N (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__17520__A (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA__17520__B (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA__17520__C (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__17520__D (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__17521__A1 (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA__17521__A2 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__17521__B1 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__17521__B2 (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA__17522__A (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA__17522__B (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__17523__A1 (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA__17523__A2 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__17525__A (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 ANTENNA__17525__B (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__17526__A (.DIODE(\mul1.a[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17526__B (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA__17526__C (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__17526__D (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__17527__A1 (.DIODE(\mul1.a[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17527__B2 (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA__17530__A1 (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA__17530__A2 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__17540__A1 (.DIODE(\mul1.a[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17540__A2 (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__17542__A (.DIODE(\mul1.a[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17542__B (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__17543__A (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__17543__B (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__17543__C (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA__17544__A1 (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__17544__A2 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__17544__B1 (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA__17544__B2 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__17545__A1 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__17551__A1 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__17551__B1 (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA__17552__A (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__17552__D (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA__17553__C (.DIODE(net630));
 sky130_fd_sc_hd__diode_2 ANTENNA__17554__A1_N (.DIODE(net630));
 sky130_fd_sc_hd__diode_2 ANTENNA__17556__A (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__17556__B (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA__17557__A (.DIODE(net625));
 sky130_fd_sc_hd__diode_2 ANTENNA__17557__B (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__17557__C (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA__17557__D (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA__17558__A1 (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__17558__A2 (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA__17558__B1 (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA__17596__A (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__17596__B (.DIODE(_04209_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17597__A2 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__17597__B1 (.DIODE(_09062_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17597__B2 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__17597__C1 (.DIODE(_03056_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17599__A (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA__17599__B (.DIODE(_04325_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17600__A1 (.DIODE(net325));
 sky130_fd_sc_hd__diode_2 ANTENNA__17600__A2 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__17604__A1 (.DIODE(net320));
 sky130_fd_sc_hd__diode_2 ANTENNA__17604__A2 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__17604__B1 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__17604__B2 (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA__17606__A (.DIODE(net321));
 sky130_fd_sc_hd__diode_2 ANTENNA__17606__B (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA__17606__C (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__17606__D (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__17608__A (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA__17608__B (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA__17608__C (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__17608__D (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__17610__A1 (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA__17610__A2 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__17610__B1 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__17610__B2 (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA__17611__A (.DIODE(net317));
 sky130_fd_sc_hd__diode_2 ANTENNA__17611__B (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__17612__A1 (.DIODE(net317));
 sky130_fd_sc_hd__diode_2 ANTENNA__17612__A2 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__17619__A (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA__17619__B (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA__17619__C (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__17619__D (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__17620__A1 (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA__17620__A2 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__17620__B1 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__17620__B2 (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA__17621__C (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA__17621__D (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__17622__A1_N (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA__17622__A2_N (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__17636__A (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__17636__B (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__17637__A (.DIODE(net277));
 sky130_fd_sc_hd__diode_2 ANTENNA__17637__B (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA__17637__C (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__17638__A1 (.DIODE(net277));
 sky130_fd_sc_hd__diode_2 ANTENNA__17638__A2 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__17638__B1 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__17638__B2 (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA__17639__A1 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__17641__A (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA__17641__B (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__17642__A (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA__17642__B (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA__17642__C (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__17643__A1 (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA__17643__A2 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__17643__B1 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__17643__B2 (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA__17644__A1 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__17646__A1 (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 ANTENNA__17646__A2 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__17656__A1 (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__17656__A2 (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__17656__B2 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__17657__A (.DIODE(net630));
 sky130_fd_sc_hd__diode_2 ANTENNA__17657__B (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__17657__C (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__17657__D (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA__17658__A1 (.DIODE(net630));
 sky130_fd_sc_hd__diode_2 ANTENNA__17658__A2 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__17658__B1 (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA__17658__B2 (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__17659__A (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__17659__B (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__17660__A1 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__17660__A2 (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__17665__A2 (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA__17665__B1 (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA__17666__A (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__17666__C (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA__17666__D (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA__17667__C (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__17668__A1_N (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__17670__A (.DIODE(\mul1.b[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17670__B (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA__17671__B (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__17671__C (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA__17671__D (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA__17672__A1 (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__17672__A2 (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA__17672__B1 (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA__17711__A2 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__17711__B1 (.DIODE(_09176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17711__B2 (.DIODE(_03050_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17720__A (.DIODE(net317));
 sky130_fd_sc_hd__diode_2 ANTENNA__17720__B (.DIODE(net321));
 sky130_fd_sc_hd__diode_2 ANTENNA__17720__C (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__17720__D (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__17721__A1 (.DIODE(net317));
 sky130_fd_sc_hd__diode_2 ANTENNA__17721__A2 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__17721__B1 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__17721__B2 (.DIODE(net321));
 sky130_fd_sc_hd__diode_2 ANTENNA__17723__C (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA__17723__D (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__17724__A1_N (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA__17724__A2_N (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__17726__A (.DIODE(\mul1.a[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17726__B (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA__17726__C (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__17726__D (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__17727__A1 (.DIODE(\mul1.a[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17727__A2 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__17727__B1 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__17727__B2 (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA__17729__C (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA__17729__D (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__17730__A1_N (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA__17730__A2_N (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__17738__A1 (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__17738__A2 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__17738__B2 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__17739__A (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__17739__B (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA__17739__C (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__17739__D (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__17740__A1 (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__17740__A2 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__17740__B1 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__17740__B2 (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA__17741__A (.DIODE(\mul1.a[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17741__B (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__17742__A1 (.DIODE(\mul1.a[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17742__A2 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__17757__A (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA__17757__B (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__17758__A (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA__17758__B (.DIODE(net277));
 sky130_fd_sc_hd__diode_2 ANTENNA__17758__C (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__17759__A1 (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA__17759__A2 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__17759__B1 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__17759__B2 (.DIODE(net277));
 sky130_fd_sc_hd__diode_2 ANTENNA__17760__A1 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__17762__A (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA__17762__B (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__17763__A (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__17763__B (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA__17763__C (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__17763__D (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__17764__A1 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__17764__A2 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__17764__B1 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__17764__B2 (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA__17767__A1 (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA__17767__A2 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__17767__B2 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__17778__A (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__17778__B (.DIODE(net629));
 sky130_fd_sc_hd__diode_2 ANTENNA__17778__C (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__17778__D (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__17779__A1 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__17779__A2 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__17779__B1 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__17779__B2 (.DIODE(net630));
 sky130_fd_sc_hd__diode_2 ANTENNA__17780__A (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__17780__B (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__17781__A1 (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__17781__A2 (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__17786__B (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA__17787__A2 (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA__17787__B1 (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA__17788__C (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA__17789__A1 (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA__17791__A (.DIODE(\mul1.b[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17791__B (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA__17792__B (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__17792__C (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA__17792__D (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA__17793__A1 (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__17793__A2 (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA__17833__A (.DIODE(_03049_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17833__B (.DIODE(_09297_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17834__A (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA__17834__B (.DIODE(_04449_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17835__A2 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__17835__B1 (.DIODE(_03056_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17836__B1 (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__17843__B1 (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA__17843__C1 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__17844__A1 (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA__17844__A2 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__17854__A (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA__17854__B (.DIODE(net317));
 sky130_fd_sc_hd__diode_2 ANTENNA__17854__C (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__17854__D (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__17856__A1 (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA__17856__A2 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__17856__B1 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__17856__B2 (.DIODE(net317));
 sky130_fd_sc_hd__diode_2 ANTENNA__17857__A (.DIODE(net321));
 sky130_fd_sc_hd__diode_2 ANTENNA__17857__B (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__17858__A1 (.DIODE(net321));
 sky130_fd_sc_hd__diode_2 ANTENNA__17858__A2 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__17860__A (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA__17860__B (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__17861__A (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA__17861__B (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA__17861__C (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__17861__D (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__17862__A1 (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA__17862__A2 (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__17862__B1 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__17862__B2 (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA__17871__A1 (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA__17871__A2 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__17871__B2 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__17872__A (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA__17872__B (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__17872__C (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__17872__D (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__17873__A1 (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA__17873__A2 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__17873__B1 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__17873__B2 (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__17874__A (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA__17874__B (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__17875__A1 (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA__17875__A2 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__17893__A (.DIODE(net277));
 sky130_fd_sc_hd__diode_2 ANTENNA__17893__B (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__17894__A (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA__17894__B (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA__17894__C (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__17895__A1 (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA__17895__A2 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__17895__B1 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__17895__B2 (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA__17896__A1 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__17898__A (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA__17898__B (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__17899__A (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__17899__B (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__17899__C (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__17899__D (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__17900__A1 (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__17900__A2 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__17900__B1 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__17900__B2 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__17914__A2 (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA__17914__B2 (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA__17915__A (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__17915__B (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__17915__C (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__17915__D (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA__17916__A1 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__17916__A2 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__17916__B1 (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA__17916__B2 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__17917__A (.DIODE(net629));
 sky130_fd_sc_hd__diode_2 ANTENNA__17917__B (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__17918__A1 (.DIODE(net629));
 sky130_fd_sc_hd__diode_2 ANTENNA__17918__A2 (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__17924__A (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__17924__B (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA__17925__C (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA__17925__D (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA__17926__A2 (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA__17926__B1 (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA__17929__A (.DIODE(\mul1.b[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17930__B (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__17930__D (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA__17931__A1 (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__17931__B1 (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA__17965__B (.DIODE(_09306_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17966__A (.DIODE(_09306_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17967__A (.DIODE(_09292_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17968__A (.DIODE(_09304_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17969__A (.DIODE(_09304_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17971__A (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__17971__B (.DIODE(_04588_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17972__A2 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__17972__B1 (.DIODE(_09434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17972__B2 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__17973__S (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__17974__A1 (.DIODE(_09292_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17976__A1 (.DIODE(net321));
 sky130_fd_sc_hd__diode_2 ANTENNA__17976__A2 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__17976__B1 (.DIODE(\mul1.b[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17976__B2 (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA__17977__A (.DIODE(\mul1.a[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17977__B (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA__17977__C (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__17977__D (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__17991__A (.DIODE(net306));
 sky130_fd_sc_hd__diode_2 ANTENNA__17991__B (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA__17991__C (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__17991__D (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__17992__A1 (.DIODE(net306));
 sky130_fd_sc_hd__diode_2 ANTENNA__17992__A2 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__17992__B1 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__17992__B2 (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA__17994__A (.DIODE(net316));
 sky130_fd_sc_hd__diode_2 ANTENNA__17994__B (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__17996__A (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA__17996__B (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__17997__A (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA__17997__B (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA__17997__C (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__17997__D (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__17998__A1 (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA__17998__A2 (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__17998__B1 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__17998__B2 (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA__18001__A1 (.DIODE(net306));
 sky130_fd_sc_hd__diode_2 ANTENNA__18001__A2 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__18007__A1 (.DIODE(net277));
 sky130_fd_sc_hd__diode_2 ANTENNA__18007__A2 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__18007__B2 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__18008__A (.DIODE(net277));
 sky130_fd_sc_hd__diode_2 ANTENNA__18008__B (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA__18008__C (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__18008__D (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__18009__A1 (.DIODE(net277));
 sky130_fd_sc_hd__diode_2 ANTENNA__18009__A2 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__18009__B1 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__18009__B2 (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA__18010__A (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__18010__B (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__18011__A1 (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__18011__A2 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__18028__A (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA__18028__B (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__18029__A1 (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA__18029__A2 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__18029__B1 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__18029__B2 (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA__18030__A (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA__18030__B (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA__18030__C (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__18030__D (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__18033__A (.DIODE(net629));
 sky130_fd_sc_hd__diode_2 ANTENNA__18033__B (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__18033__C (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__18033__D (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__18034__A1 (.DIODE(net629));
 sky130_fd_sc_hd__diode_2 ANTENNA__18034__A2 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__18034__B1 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__18034__B2 (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__18035__A (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__18035__B (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__18036__A1 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__18036__A2 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__18049__A1 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__18049__A2 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__18049__B1 (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA__18049__B2 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__18050__A (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__18050__B (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__18050__C (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__18050__D (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA__18051__C (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__18051__D (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__18052__A1_N (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__18052__A2_N (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__18058__A (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__18058__B (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA__18059__C (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA__18060__A2 (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA__18063__A (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__18064__C (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA__18064__D (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__18065__A2 (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA__18065__B1 (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__18102__A (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA__18102__B (.DIODE(_04719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18103__A2 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__18103__B1 (.DIODE(_09564_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18103__B2 (.DIODE(_03050_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18109__A1 (.DIODE(net316));
 sky130_fd_sc_hd__diode_2 ANTENNA__18109__A2 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__18110__A (.DIODE(net316));
 sky130_fd_sc_hd__diode_2 ANTENNA__18110__B (.DIODE(\mul1.a[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__18110__C (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__18110__D (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__18111__A1 (.DIODE(net316));
 sky130_fd_sc_hd__diode_2 ANTENNA__18111__A2 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__18111__B1 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__18111__B2 (.DIODE(\mul1.a[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__18112__C (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA__18112__D (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__18113__A1_N (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA__18113__A2_N (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__18130__A1 (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA__18130__A2 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__18130__B1 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__18130__B2 (.DIODE(net306));
 sky130_fd_sc_hd__diode_2 ANTENNA__18131__A (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA__18131__B (.DIODE(net306));
 sky130_fd_sc_hd__diode_2 ANTENNA__18131__C (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__18132__A1 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__18133__A (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA__18133__B (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__18135__A (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA__18135__B (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA__18135__C (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__18135__D (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__18136__A1 (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA__18136__A2 (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__18136__B1 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__18136__B2 (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA__18137__A (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA__18137__B (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__18138__A1 (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA__18138__A2 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__18146__A (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA__18146__B (.DIODE(net276));
 sky130_fd_sc_hd__diode_2 ANTENNA__18146__C (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__18146__D (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__18147__A1 (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA__18147__A2 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__18147__B1 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__18147__B2 (.DIODE(net276));
 sky130_fd_sc_hd__diode_2 ANTENNA__18148__C (.DIODE(net281));
 sky130_fd_sc_hd__diode_2 ANTENNA__18148__D (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__18149__A1_N (.DIODE(net281));
 sky130_fd_sc_hd__diode_2 ANTENNA__18149__A2_N (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__18165__A1 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__18165__A2 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__18165__B1 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__18165__B2 (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA__18166__A (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__18166__B (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA__18166__C (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__18166__D (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__18167__A (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA__18167__B (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__18168__A1 (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA__18168__A2 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__18170__A1 (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA__18170__A2 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__18170__B1 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__18170__B2 (.DIODE(net626));
 sky130_fd_sc_hd__diode_2 ANTENNA__18171__A (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA__18171__B (.DIODE(net626));
 sky130_fd_sc_hd__diode_2 ANTENNA__18171__C (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__18171__D (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__18172__C (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__18172__D (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__18173__A1_N (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__18173__A2_N (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__18187__A1 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__18187__A2 (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA__18187__B2 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__18188__A (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__18188__B (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__18188__C (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA__18189__C (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__18189__D (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__18190__A1_N (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__18190__A2_N (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__18196__A (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__18196__B (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA__18198__B1 (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA__18201__A (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__18201__B (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA__18202__C (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__18202__D (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__18203__A2 (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__18203__B1 (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__18242__A1 (.DIODE(_09292_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18244__B2 (.DIODE(_09304_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18246__A2_N (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__18246__B1 (.DIODE(_04862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18246__B2 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__18247__A1 (.DIODE(_03049_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18247__A2 (.DIODE(_09707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18248__S (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__18254__A1 (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA__18254__A2 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__18254__B2 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__18255__A1 (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA__18255__A2 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__18255__B1 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__18255__B2 (.DIODE(net316));
 sky130_fd_sc_hd__diode_2 ANTENNA__18256__A (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA__18256__B (.DIODE(net316));
 sky130_fd_sc_hd__diode_2 ANTENNA__18256__C (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__18256__D (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__18257__A1_N (.DIODE(net321));
 sky130_fd_sc_hd__diode_2 ANTENNA__18257__A2_N (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__18258__C (.DIODE(net321));
 sky130_fd_sc_hd__diode_2 ANTENNA__18258__D (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__18271__A (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA__18271__B (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__18278__A1 (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA__18278__A2 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__18278__B1 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__18278__B2 (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA__18279__A (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA__18279__B (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA__18279__C (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__18279__D (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__18280__A1 (.DIODE(net306));
 sky130_fd_sc_hd__diode_2 ANTENNA__18280__A2 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__18281__A (.DIODE(net306));
 sky130_fd_sc_hd__diode_2 ANTENNA__18281__B (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__18283__A (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA__18283__B (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__18284__A1 (.DIODE(net281));
 sky130_fd_sc_hd__diode_2 ANTENNA__18284__A2 (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__18284__B1 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__18284__B2 (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA__18285__A (.DIODE(net281));
 sky130_fd_sc_hd__diode_2 ANTENNA__18285__B (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA__18285__C (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__18285__D (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__18294__A1 (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA__18294__A2 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__18294__B1 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__18294__B2 (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA__18295__A (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA__18295__B (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA__18295__C (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__18295__D (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__18296__A1_N (.DIODE(net276));
 sky130_fd_sc_hd__diode_2 ANTENNA__18296__A2_N (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__18297__C (.DIODE(net276));
 sky130_fd_sc_hd__diode_2 ANTENNA__18297__D (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__18312__A1 (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA__18312__A2 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__18312__B1 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__18312__B2 (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA__18313__A (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA__18313__B (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA__18313__C (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__18313__D (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__18314__A (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__18314__B (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__18315__A1 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__18315__A2 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__18317__A (.DIODE(net626));
 sky130_fd_sc_hd__diode_2 ANTENNA__18317__B (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__18318__A1 (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA__18318__A2 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__18318__B1 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__18318__B2 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__18319__A (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA__18319__B (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__18319__C (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__18319__D (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__18333__A1 (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__18333__A2 (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA__18334__A1 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__18334__B1 (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA__18334__B2 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__18335__A (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__18335__B (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__18335__D (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA__18336__A (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__18336__B (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__18336__D (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA__18337__A1 (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__18337__A2 (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA__18338__A (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__18338__B (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA__18344__A (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__18345__D (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA__18346__A2 (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA__18346__B1 (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA__18349__A (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__18349__B (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__18350__C (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__18351__A2 (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__18391__A (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__18391__B (.DIODE(_05006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18392__A2 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__18392__B1 (.DIODE(_09851_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18392__B2 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__18393__S (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__18397__A1 (.DIODE(_09305_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18399__A1 (.DIODE(\mul1.a[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__18399__A2 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__18399__B1 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__18399__B2 (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA__18400__A (.DIODE(\mul1.a[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__18400__B (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA__18400__C (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__18400__D (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__18403__A1 (.DIODE(net306));
 sky130_fd_sc_hd__diode_2 ANTENNA__18403__A2 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__18403__B1 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__18403__B2 (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA__18404__A (.DIODE(net306));
 sky130_fd_sc_hd__diode_2 ANTENNA__18404__B (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA__18404__C (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__18404__D (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__18405__A1_N (.DIODE(net316));
 sky130_fd_sc_hd__diode_2 ANTENNA__18405__A2_N (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__18406__C (.DIODE(net316));
 sky130_fd_sc_hd__diode_2 ANTENNA__18406__D (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__18426__A1 (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA__18426__A2 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__18426__B1 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__18426__B2 (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA__18427__A (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA__18427__B (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA__18427__C (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__18427__D (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__18428__A1 (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA__18428__A2 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__18429__A (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA__18429__B (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__18431__A1 (.DIODE(net276));
 sky130_fd_sc_hd__diode_2 ANTENNA__18431__A2 (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__18431__B1 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__18431__B2 (.DIODE(net281));
 sky130_fd_sc_hd__diode_2 ANTENNA__18432__A (.DIODE(net276));
 sky130_fd_sc_hd__diode_2 ANTENNA__18432__B (.DIODE(net281));
 sky130_fd_sc_hd__diode_2 ANTENNA__18432__C (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__18432__D (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__18433__A1_N (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA__18433__A2_N (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__18434__C (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA__18434__D (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__18443__A1 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__18443__A2 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__18443__B1 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__18443__B2 (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA__18444__A (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__18444__B (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA__18444__C (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__18444__D (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__18445__A1_N (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA__18445__A2_N (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__18446__C (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA__18446__D (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__18461__A1 (.DIODE(net626));
 sky130_fd_sc_hd__diode_2 ANTENNA__18461__A2 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__18461__B1 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__18461__B2 (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA__18462__A (.DIODE(net626));
 sky130_fd_sc_hd__diode_2 ANTENNA__18462__B (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA__18462__C (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__18462__D (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__18463__A1 (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA__18463__A2 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__18464__A (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA__18464__B (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__18466__A1 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__18466__A2 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__18466__B1 (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA__18466__B2 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__18467__A (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__18467__B (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__18467__C (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__18467__D (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA__18468__A1_N (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA__18468__A2_N (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__18469__C (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA__18469__D (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__18482__A1 (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__18483__A1 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__18483__A2 (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA__18483__B2 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__18484__A (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__18484__B (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__18484__C (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA__18485__A1 (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__18485__A2 (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA__18486__A (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__18486__B (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA__18492__A (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__18493__C (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA__18493__D (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__18494__A2 (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA__18494__B1 (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__18497__A (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__18497__B (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__18499__A1 (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__18538__A (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__18538__B (.DIODE(_05156_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18539__A2 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__18539__B1 (.DIODE(_09997_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18539__B2 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__18544__A1 (.DIODE(net316));
 sky130_fd_sc_hd__diode_2 ANTENNA__18544__A2 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__18544__B1 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__18544__B2 (.DIODE(net321));
 sky130_fd_sc_hd__diode_2 ANTENNA__18545__A (.DIODE(net316));
 sky130_fd_sc_hd__diode_2 ANTENNA__18545__B (.DIODE(net321));
 sky130_fd_sc_hd__diode_2 ANTENNA__18545__C (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__18546__A1 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__18547__A (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA__18547__B (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__18553__A1 (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA__18553__A2 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__18553__B1 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__18553__B2 (.DIODE(net306));
 sky130_fd_sc_hd__diode_2 ANTENNA__18554__A (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA__18554__B (.DIODE(net306));
 sky130_fd_sc_hd__diode_2 ANTENNA__18554__C (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__18554__D (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__18555__A1_N (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA__18555__A2_N (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__18556__C (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA__18556__D (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__18578__A1 (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA__18578__A2 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__18578__B1 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__18578__B2 (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA__18579__A (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA__18579__B (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA__18579__C (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__18579__D (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__18580__A1 (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA__18580__A2 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__18581__A (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA__18581__B (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__18583__A1 (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA__18583__B2 (.DIODE(net276));
 sky130_fd_sc_hd__diode_2 ANTENNA__18584__A (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA__18584__B (.DIODE(net276));
 sky130_fd_sc_hd__diode_2 ANTENNA__18585__A1_N (.DIODE(net281));
 sky130_fd_sc_hd__diode_2 ANTENNA__18585__A2_N (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__18586__C (.DIODE(net281));
 sky130_fd_sc_hd__diode_2 ANTENNA__18586__D (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__18595__A1 (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA__18595__A2 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__18595__B1 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__18595__B2 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__18596__A (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA__18596__B (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__18596__C (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__18596__D (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__18597__A1 (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA__18597__A2 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__18598__A (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA__18598__B (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__18615__A1 (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA__18615__A2 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__18615__B1 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__18615__B2 (.DIODE(net626));
 sky130_fd_sc_hd__diode_2 ANTENNA__18616__A (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA__18616__B (.DIODE(net626));
 sky130_fd_sc_hd__diode_2 ANTENNA__18616__C (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__18616__D (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__18619__A (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA__18619__B (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__18621__A1 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__18621__A2 (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA__18621__B2 (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__18622__A (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__18622__B (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__18622__C (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA__18623__A1 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__18623__A2 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__18624__A (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__18624__B (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__18635__A1 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__18635__A2 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__18635__A3 (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA__18636__A1 (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__18637__A1 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__18637__B2 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__18638__A (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__18638__B (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__18639__A1 (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__18639__A2 (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA__18640__A (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__18640__B (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA__18645__B (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA__18646__A2 (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__18646__B1 (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__18647__C (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__18648__A1 (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__18650__A (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__18651__A1 (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__18651__B1 (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__18652__B (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__18652__D (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__18689__A (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__18689__B (.DIODE(_05305_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18690__A2 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__18690__B1 (.DIODE(_10147_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18690__B2 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__18694__A1 (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA__18694__A2 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__18694__B1 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__18694__B2 (.DIODE(net316));
 sky130_fd_sc_hd__diode_2 ANTENNA__18696__A (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA__18696__B (.DIODE(net316));
 sky130_fd_sc_hd__diode_2 ANTENNA__18696__C (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__18696__D (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__18697__A1_N (.DIODE(net321));
 sky130_fd_sc_hd__diode_2 ANTENNA__18697__A2_N (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__18698__B (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__18698__C (.DIODE(net321));
 sky130_fd_sc_hd__diode_2 ANTENNA__18700__A1 (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA__18700__A2 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__18700__B2 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__18703__A (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA__18703__B (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA__18710__A1 (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA__18710__A2 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__18710__B1 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__18710__B2 (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA__18711__A (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA__18711__B (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA__18711__C (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__18711__D (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__18712__A1 (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA__18712__A2 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__18713__A (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA__18713__B (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__18731__A1 (.DIODE(net281));
 sky130_fd_sc_hd__diode_2 ANTENNA__18731__A2 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__18731__B1 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__18731__B2 (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA__18732__A (.DIODE(net281));
 sky130_fd_sc_hd__diode_2 ANTENNA__18732__B (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA__18732__C (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__18732__D (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__18734__A (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA__18734__B (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__18736__A1 (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA__18736__B2 (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA__18737__A (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA__18737__B (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA__18738__A (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA__18738__B (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA__18738__C (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__18739__A1 (.DIODE(net276));
 sky130_fd_sc_hd__diode_2 ANTENNA__18739__A2 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__18740__A (.DIODE(net276));
 sky130_fd_sc_hd__diode_2 ANTENNA__18740__B (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__18741__A (.DIODE(net276));
 sky130_fd_sc_hd__diode_2 ANTENNA__18741__B (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__18746__A1 (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA__18746__A2 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__18746__A3 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__18746__A4 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__18747__A1 (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA__18747__A2 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__18748__A1 (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA__18748__A2 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__18748__B1 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__18748__B2 (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA__18749__A (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA__18749__B (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA__18749__C (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__18749__D (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__18750__A1 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__18750__A2 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__18751__A (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__18751__B (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__18766__A1 (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA__18766__A2 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__18766__B1 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__18766__B2 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__18767__A (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA__18767__B (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__18767__C (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__18768__A1 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__18769__A (.DIODE(net626));
 sky130_fd_sc_hd__diode_2 ANTENNA__18769__B (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__18771__A1 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__18771__B1 (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA__18771__B2 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__18772__A (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__18772__B (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__18772__D (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA__18773__A (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__18773__B (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA__18785__A2 (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA__18785__B2 (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__18786__A1 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__18786__A2 (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA__18786__B1 (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA__18786__B2 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__18787__A (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__18787__B (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__18787__C (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA__18787__D (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA__18788__A1 (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__18788__A2 (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA__18789__A (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__18789__B (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA__18794__A2 (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__18794__B1 (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__18795__C (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__18795__D (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__18796__C (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__18796__D (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__18797__A1_N (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__18797__A2_N (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__18799__A (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__18800__A1 (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__18800__A2 (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA__18800__B1 (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__18801__B (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__18801__C (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__18801__D (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__18842__A (.DIODE(_03049_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18842__B (.DIODE(_10299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18843__A2 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__18843__B1 (.DIODE(_05457_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18843__B2 (.DIODE(_03052_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18848__A1 (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA__18848__A2 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__18848__B1 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__18848__B2 (.DIODE(net306));
 sky130_fd_sc_hd__diode_2 ANTENNA__18849__A (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA__18849__B (.DIODE(net306));
 sky130_fd_sc_hd__diode_2 ANTENNA__18849__C (.DIODE(\mul1.b[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__18849__D (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__18850__A1_N (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA__18850__A2_N (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__18851__C (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA__18851__D (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__18856__A1 (.DIODE(net316));
 sky130_fd_sc_hd__diode_2 ANTENNA__18856__A2 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__18856__B1 (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA__18856__B2 (.DIODE(net321));
 sky130_fd_sc_hd__diode_2 ANTENNA__18857__A (.DIODE(net316));
 sky130_fd_sc_hd__diode_2 ANTENNA__18857__B (.DIODE(net321));
 sky130_fd_sc_hd__diode_2 ANTENNA__18857__C (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__18857__D (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA__18858__A1 (.DIODE(net325));
 sky130_fd_sc_hd__diode_2 ANTENNA__18858__A2 (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__18859__A (.DIODE(net325));
 sky130_fd_sc_hd__diode_2 ANTENNA__18859__B (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__18868__A1 (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA__18868__A2 (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA__18868__A3 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__18868__A4 (.DIODE(\mul1.b[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__18870__A2 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__18870__B1 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__18870__B2 (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA__18871__B (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA__18871__C (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__18871__D (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__18872__A1 (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA__18872__A2 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__18873__A (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA__18873__B (.DIODE(\mul1.b[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__18891__A1 (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA__18891__A2 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__18891__B1 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__18891__B2 (.DIODE(net276));
 sky130_fd_sc_hd__diode_2 ANTENNA__18892__A (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA__18892__B (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA__18892__C (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__18892__D (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__18893__A1 (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA__18893__A2 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__18894__A (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA__18894__B (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__18896__A1 (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA__18896__A2 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__18896__B2 (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA__18897__A (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA__18897__B (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__18897__C (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__18898__B (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA__18898__C (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__18899__A1 (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA__18900__A (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA__18901__A (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA__18901__B (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__18907__A1 (.DIODE(net626));
 sky130_fd_sc_hd__diode_2 ANTENNA__18907__A2 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__18907__B2 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__18908__A1 (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA__18908__A2 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__18908__B1 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__18908__B2 (.DIODE(net626));
 sky130_fd_sc_hd__diode_2 ANTENNA__18909__A (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA__18909__B (.DIODE(net626));
 sky130_fd_sc_hd__diode_2 ANTENNA__18909__C (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__18909__D (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__18910__A1 (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__18910__A2 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__18911__A (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA__18911__B (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__18927__A (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__18927__B (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__18928__A1 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__18928__A2 (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA__18928__B2 (.DIODE(\mul1.b[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__18929__A (.DIODE(\mul1.b[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__18929__B (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__18930__A1 (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA__18932__A (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__18932__B (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA__18933__A1 (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__18933__B2 (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__18934__A (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__18934__B (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__18948__A1 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__18948__A2 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__18948__B1 (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__18949__B (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__18949__C (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__18949__D (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__18950__A1 (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA__18950__A2 (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA__18951__A (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__18951__B (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA__18956__B (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__18957__B1 (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA__18957__B2 (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__18958__A (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__18958__C (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA__18961__A (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__18961__B (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA__18962__A2 (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__18962__B1 (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__18963__B (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__18963__C (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__19002__A (.DIODE(_03049_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19002__B (.DIODE(_10458_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19003__A2 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__19003__B1 (.DIODE(_05615_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19003__B2 (.DIODE(_03052_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19008__A_N (.DIODE(net321));
 sky130_fd_sc_hd__diode_2 ANTENNA__19008__B (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA__19008__C (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__19008__D (.DIODE(net316));
 sky130_fd_sc_hd__diode_2 ANTENNA__19009__A1_N (.DIODE(net316));
 sky130_fd_sc_hd__diode_2 ANTENNA__19009__A2_N (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA__19009__B1 (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__19009__B2 (.DIODE(net321));
 sky130_fd_sc_hd__diode_2 ANTENNA__19012__A1 (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA__19012__A2 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__19012__B1 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__19012__B2 (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA__19013__A (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA__19013__B (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA__19013__C (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__19014__A1 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__19015__A (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA__19015__B (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__19029__A2 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__19029__B1 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__19030__C (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__19030__D (.DIODE(\mul1.b[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__19031__A1 (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA__19031__A2 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__19032__A (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA__19032__B (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__19050__A1 (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA__19050__A2 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__19050__B1 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__19050__B2 (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA__19051__A (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA__19051__B (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA__19051__C (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__19052__A1 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__19053__A (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA__19053__B (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__19055__B2 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__19056__A (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA__19056__B (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__19056__C (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__19056__D (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__19057__A (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA__19057__B (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__19058__A1 (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA__19058__A2 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__19059__A (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA__19059__B (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__19060__A (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA__19060__B (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__19066__A1 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__19066__A2 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__19066__B2 (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA__19067__A1 (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__19067__A2 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__19067__B1 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__19068__A (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__19068__C (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__19068__D (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__19069__A1 (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__19069__A2 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__19070__A (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__19070__B (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__19086__A1 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__19086__B2 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__19087__A (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__19087__B (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__19087__D (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA__19089__A (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__19089__B (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__19091__A1 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__19091__B2 (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__19092__A (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__19092__B (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__19093__A (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__19093__B (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA__19107__A2 (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__19108__A1 (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA__19108__A2 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__19108__B1 (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__19108__B2 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__19109__A (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__19109__B (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA__19109__C (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__19109__D (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__19110__A1 (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__19110__A2 (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA__19111__A (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__19111__B (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA__19116__B1 (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA__19117__C (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA__19119__B (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__19122__B (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__19123__B (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__19123__C (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__19124__A2 (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__19124__B1_N (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__19125__A (.DIODE(\mul1.b[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__19125__B (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA__19168__A1 (.DIODE(_09305_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19169__B (.DIODE(_10624_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19170__A2 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__19170__B1 (.DIODE(_05784_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19170__B2 (.DIODE(_03052_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19171__A1 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__19171__A2 (.DIODE(_10625_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19173__A2 (.DIODE(_10624_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19178__A1 (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA__19178__A2 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__19178__B1 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__19178__B2 (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA__19179__A (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA__19179__B (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA__19179__C (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__19180__A1 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__19181__A (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA__19181__B (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__19183__A1_N (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__19185__A_N (.DIODE(net317));
 sky130_fd_sc_hd__diode_2 ANTENNA__19185__B (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA__19185__C (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__19185__D (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA__19187__A1_N (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA__19187__A2_N (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA__19187__B1 (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__19187__B2 (.DIODE(net317));
 sky130_fd_sc_hd__diode_2 ANTENNA__19196__A3 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__19196__A4 (.DIODE(\mul1.b[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__19197__A1 (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA__19197__A2 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__19197__B2 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__19198__A1 (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA__19198__A2 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__19198__B1 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__19199__A (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA__19199__C (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__19199__D (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__19200__A2 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__19201__B (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__19220__A1 (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA__19220__A2 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__19220__B1 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__19220__B2 (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA__19221__A (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA__19221__B (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA__19221__C (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__19222__A1 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__19223__A (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA__19223__B (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__19225__A1 (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__19225__A2 (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__19225__B1 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__19226__A (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA__19226__C (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__19226__D (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__19227__A (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__19227__C (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__19227__D (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__19228__A1 (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA__19228__A2 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__19229__A (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA__19229__B (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__19230__A (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA__19230__B (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__19237__A1 (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__19237__A2 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__19237__B2 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__19238__A (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__19238__B (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__19238__C (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__19239__A2 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__19240__B (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__19256__A1 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__19256__A2 (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA__19256__B1 (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA__19256__B2 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__19257__A (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__19257__B (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__19257__C (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA__19257__D (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA__19259__A (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__19261__A1 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__19261__B1 (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA__19261__B2 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__19262__A (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__19262__B (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__19262__D (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA__19263__A1 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__19264__A (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__19277__A2 (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__19278__A1 (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA__19278__A2 (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__19278__B1 (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__19278__B2 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__19279__A (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__19279__B (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA__19279__C (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__19279__D (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__19280__A1 (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__19280__A2 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__19281__A (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__19281__B (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__19286__A2 (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA__19286__B1 (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__19287__A1 (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__19290__S (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__19323__A2_N (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__19323__B1 (.DIODE(_05935_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19323__B2 (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA__19324__A1 (.DIODE(_03049_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19324__A2 (.DIODE(_10777_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19330__A2 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__19330__B1 (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__19330__B2 (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA__19331__A (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA__19331__B (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA__19331__C (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__19332__A1 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__19333__A (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA__19333__B (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__19335__A1_N (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__19337__A_N (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA__19337__B (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__19337__C (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__19337__D (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA__19339__A1_N (.DIODE(net306));
 sky130_fd_sc_hd__diode_2 ANTENNA__19339__A2_N (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__19339__B1 (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__19339__B2 (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA__19349__A1 (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA__19349__A2 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__19349__B2 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__19350__A1 (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA__19350__A2 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__19350__B1 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__19350__B2 (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA__19351__A (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA__19351__B (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA__19351__C (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__19351__D (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__19352__A2 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__19353__B (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__19372__A1 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__19372__A2 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__19372__B1 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__19372__B2 (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA__19373__A (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__19373__B (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA__19373__C (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__19374__A1 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__19375__A (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA__19375__B (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__19377__A2 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__19377__B1 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__19377__B2 (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA__19378__B (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__19378__C (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__19378__D (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__19379__B (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__19379__C (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__19379__D (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__19380__A2 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__19381__B (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__19382__B (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__19389__A1 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__19389__B2 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__19390__A (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__19390__B (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__19391__A1 (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__19391__A2 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__19392__A (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__19392__B (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__19408__A1 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__19408__A2 (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA__19408__B2 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__19409__A (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__19409__B (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__19409__C (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA__19411__A (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__19413__A1 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__19413__A2 (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA__19413__B1 (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__19413__B2 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__19414__A (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__19414__B (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__19414__C (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA__19414__D (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__19416__A1 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__19416__A2 (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA__19417__A (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__19417__B (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA__19428__B2 (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__19429__A1 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__19429__A2 (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__19429__B2 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__19430__A (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__19430__B (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA__19430__C (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__19431__A1 (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__19431__A2 (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__19432__A (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__19432__B (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__19437__A2 (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__19437__B1 (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__19438__C (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA__19438__D (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__19439__B (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA__19445__A (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__19474__C_N (.DIODE(_10624_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19477__A2_N (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__19477__B1 (.DIODE(_06090_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19477__B2 (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA__19478__A1 (.DIODE(_03049_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19478__A2 (.DIODE(_00660_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19486__A1 (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA__19486__A2 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__19486__B1 (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__19486__B2 (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA__19487__A (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA__19487__B (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA__19487__C (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__19488__A1 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__19489__A (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA__19489__B (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__19491__A1_N (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__19493__A_N (.DIODE(net306));
 sky130_fd_sc_hd__diode_2 ANTENNA__19493__B (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__19493__C (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__19493__D (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA__19495__A1_N (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA__19495__A2_N (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__19495__B1 (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__19495__B2 (.DIODE(net306));
 sky130_fd_sc_hd__diode_2 ANTENNA__19505__A1 (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA__19505__A2 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__19505__B2 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__19506__A1 (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA__19506__A2 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__19506__B1 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__19506__B2 (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA__19507__A (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA__19507__B (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA__19507__C (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__19507__D (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__19508__A1 (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA__19508__A2 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__19509__A (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA__19509__B (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__19528__A1 (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA__19528__A2 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__19528__B1 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__19528__B2 (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__19529__A (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA__19529__B (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__19529__C (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__19530__A1 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__19531__A (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA__19531__B (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__19533__A1 (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA__19533__A2 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__19533__B1 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__19533__B2 (.DIODE(net626));
 sky130_fd_sc_hd__diode_2 ANTENNA__19534__A (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA__19534__B (.DIODE(net626));
 sky130_fd_sc_hd__diode_2 ANTENNA__19534__C (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__19534__D (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__19535__A (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA__19535__C (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__19535__D (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__19536__A1 (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA__19536__A2 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__19537__A (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA__19537__B (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__19538__A (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA__19538__B (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__19544__A1 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__19545__A1 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__19545__A2 (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA__19545__B2 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__19546__A (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__19546__B (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__19547__A1 (.DIODE(\mul1.b[17] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__19548__A (.DIODE(\mul1.b[17] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__19565__A1 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__19565__B1 (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA__19565__B2 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__19566__A (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__19566__B (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__19567__A1 (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA__19568__A (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__19568__B (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA__19570__A1 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__19570__A2 (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__19570__B1 (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__19570__B2 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__19571__A (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__19571__B (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__19571__C (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__19571__D (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__19573__A1 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__19573__A2 (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA__19574__A (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__19574__B (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA__19575__A (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__19575__B (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA__19586__C (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__19587__C (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__19588__B1 (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__19589__A2 (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__19590__A (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__19590__B (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA__19600__A1 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__19600__B1 (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA__19600__B2 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__19601__A (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__19601__B (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__19601__D (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__19602__A1 (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__19602__A2 (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__19603__A (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__19636__A (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA__19636__B (.DIODE(_06244_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19637__A2 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__19637__B1 (.DIODE(_00818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19637__B2 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__19638__S (.DIODE(_03055_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19643__A1 (.DIODE(net281));
 sky130_fd_sc_hd__diode_2 ANTENNA__19643__A2 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__19643__B1 (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__19643__B2 (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA__19644__A (.DIODE(net281));
 sky130_fd_sc_hd__diode_2 ANTENNA__19644__C (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__19644__D (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__19646__B (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__19648__A1_N (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__19650__A_N (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA__19650__B (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__19650__C (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__19650__D (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA__19652__A1_N (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA__19652__A2_N (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__19652__B1 (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__19652__B2 (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA__19662__A1 (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA__19662__A2 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__19662__B2 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__19663__A1 (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA__19663__A2 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__19663__B1 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__19663__B2 (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA__19664__A (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA__19664__B (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA__19664__C (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__19664__D (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__19665__A1 (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA__19665__A2 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__19666__A (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA__19666__B (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__19685__A1 (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA__19685__A2 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__19685__B1 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__19685__B2 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__19686__A (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA__19686__B (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA__19686__C (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__19687__A1 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__19688__A (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA__19688__B (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__19690__A2 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__19690__B1 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__19690__B2 (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA__19691__A (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA__19691__C (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__19691__D (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__19692__A (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__19692__C (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__19692__D (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__19693__A1 (.DIODE(net626));
 sky130_fd_sc_hd__diode_2 ANTENNA__19693__A2 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__19694__A (.DIODE(net626));
 sky130_fd_sc_hd__diode_2 ANTENNA__19694__B (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__19695__A (.DIODE(net626));
 sky130_fd_sc_hd__diode_2 ANTENNA__19695__B (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__19701__A1 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__19701__A2 (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA__19701__B2 (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA__19702__A1 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__19702__A2 (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA__19702__B1 (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA__19702__B2 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__19703__A (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__19703__B (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__19703__C (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA__19703__D (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA__19704__A1 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__19705__A (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__19722__A1 (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__19722__A2 (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__19723__A (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__19730__A1 (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__19730__A2 (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA__19731__A1 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__19731__A2 (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA__19731__B1 (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA__19731__B2 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__19732__A (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__19732__B (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__19732__C (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA__19732__D (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__19733__A1 (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__19734__A (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__19745__A1 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__19745__A2 (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA__19745__B1 (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA__19745__B2 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__19746__A (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__19746__B (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__19746__C (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA__19747__A1 (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA__19748__A (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__19750__A1 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__19750__A2 (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__19750__B2 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__19751__A (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__19751__B (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__19751__C (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__19752__A1 (.DIODE(\mul1.b[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__19752__A2 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__19753__A (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__19753__B (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__19790__A1 (.DIODE(_10624_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19793__A (.DIODE(_03049_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19794__A2 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__19794__B1 (.DIODE(_06402_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19794__B2 (.DIODE(_03052_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19801__A1 (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA__19801__A2 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__19801__B1 (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__19801__B2 (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA__19802__A (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA__19802__B (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA__19802__C (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__19802__D (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__19803__A2 (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__19804__B (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__19810__A_N (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA__19810__B (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__19810__C (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__19812__A2_N (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__19812__B1 (.DIODE(_02568_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19812__B2 (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA__19821__A1 (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__19821__A2 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__19821__B2 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__19822__A1 (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA__19822__A2 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__19822__B1 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__19822__B2 (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA__19823__A (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA__19823__B (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA__19823__C (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__19823__D (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__19824__A1 (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA__19824__A2 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__19825__A (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA__19825__B (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__19850__A1 (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__19851__A1 (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA__19851__A2 (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__19851__B1 (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__19851__B2 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__19852__A (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__19852__B (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA__19852__C (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__19852__D (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__19853__A1 (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__19853__A2 (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA__19854__A (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__19854__B (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA__19865__A1 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__19865__A2 (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__19865__B1 (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__19865__B2 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__19866__A (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__19866__B (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__19866__C (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA__19866__D (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__19868__A (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__19868__B (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA__19870__A1 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__19870__B2 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__19871__A (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__19871__B (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__19872__A (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__19872__B (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__19873__A1 (.DIODE(\mul1.b[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__19873__A2 (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__19874__A (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__19874__B (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__19889__A1 (.DIODE(net628));
 sky130_fd_sc_hd__diode_2 ANTENNA__19889__A2 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__19889__B1 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__19889__B2 (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__19890__A (.DIODE(net628));
 sky130_fd_sc_hd__diode_2 ANTENNA__19890__B (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__19890__C (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__19890__D (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__19892__A (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__19892__B (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__19894__A1 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__19894__A2 (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA__19894__B1 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__19894__B2 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__19895__A (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__19895__B (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__19895__C (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA__19895__D (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__19896__A (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA__19896__B (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__19904__A1 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__19904__B2 (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA__19905__A1 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__19905__A2 (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA__19905__B2 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__19906__A (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__19906__B (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__19906__C (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA__19907__A1 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__19908__A (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__19945__B (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__19946__A1 (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA__19946__A2 (.DIODE(_06552_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19946__B2 (.DIODE(_03049_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19951__A (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__19951__B (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA__19951__C (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__19952__A1 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__19952__A2 (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA__19952__B1 (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__19954__A1 (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__19954__A2 (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__19955__A (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__19955__B (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__19966__A1 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__19966__A2 (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__19966__B1 (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__19966__B2 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__19967__A (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__19967__B (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__19967__C (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__19968__A1 (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__19969__A (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__19969__B (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__19971__A1 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__19971__B1 (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__19971__B2 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__19972__A (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__19972__B (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__19972__D (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__19973__A1 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__19973__A2 (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__19974__A (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__19974__B (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__19987__A1 (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA__19987__A2 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__19987__B1 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__19987__B2 (.DIODE(net628));
 sky130_fd_sc_hd__diode_2 ANTENNA__19988__A (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA__19988__B (.DIODE(net628));
 sky130_fd_sc_hd__diode_2 ANTENNA__19988__C (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__19989__A1 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__19990__A (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__19990__B (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__19992__A1 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA__19992__A2 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__19992__B1 (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__19992__B2 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__19993__A (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__19993__B (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA__19993__C (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__19994__A1 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__19994__A2 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__19995__A (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__19995__B (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__20003__A1 (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__20003__A2 (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA__20003__B1 (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA__20003__B2 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__20004__A (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__20004__B (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__20004__C (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA__20004__D (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA__20005__A1_N (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__20005__A2_N (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 ANTENNA__20006__C (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__20006__D (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 ANTENNA__20025__A1 (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA__20025__A2 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__20025__B1 (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__20025__B2 (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA__20026__A (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA__20026__B (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA__20026__C (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__20026__D (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__20027__A1_N (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA__20027__A2_N (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__20028__C (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA__20028__D (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__20032__B (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__20032__C (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__20034__A2_N (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__20034__B1 (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__20034__B2 (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA__20045__A1 (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__20045__A2 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__20045__B1 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__20045__B2 (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__20046__A (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__20046__B (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__20046__C (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__20046__D (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__20047__A1_N (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA__20047__A2_N (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__20048__C (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA__20048__D (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__20084__A1 (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA__20084__A2 (.DIODE(_06691_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20084__B2 (.DIODE(_03049_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20085__A2 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__20088__A (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__20088__B (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__20100__A1 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__20100__A2 (.DIODE(\mul1.a[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__20100__B1 (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__20100__B2 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__20101__A (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__20101__B (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__20101__C (.DIODE(\mul1.a[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__20101__D (.DIODE(\mul1.a[27] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__20102__A1 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__20102__A2 (.DIODE(\mul1.a[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__20103__A (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__20103__B (.DIODE(\mul1.a[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__20105__A1 (.DIODE(\mul1.b[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__20105__A2 (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA__20105__B1 (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__20105__B2 (.DIODE(\mul1.b[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__20106__A (.DIODE(\mul1.b[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__20106__B (.DIODE(\mul1.b[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__20106__C (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA__20106__D (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__20107__A1_N (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__20108__C (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__20127__A1 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__20127__A2 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__20127__B1 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__20127__B2 (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA__20128__A (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA__20128__B (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__20128__C (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__20128__D (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__20129__A1 (.DIODE(net628));
 sky130_fd_sc_hd__diode_2 ANTENNA__20129__A2 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__20130__A (.DIODE(net628));
 sky130_fd_sc_hd__diode_2 ANTENNA__20130__B (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__20132__A1 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__20132__B1 (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA__20132__B2 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__20133__A (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__20133__B (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__20133__D (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA__20135__A1 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA__20135__A2 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__20136__A (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA__20136__B (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__20144__A1_N (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__20145__A1 (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__20145__A2 (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA__20145__B1 (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__20145__B2 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__20146__A (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__20146__B (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__20146__C (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA__20146__D (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__20147__A1_N (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__20147__A2_N (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA__20148__C (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__20148__D (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA__20169__A1 (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA__20169__A2 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__20169__B1 (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__20169__B2 (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA__20170__A (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA__20170__B (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA__20170__C (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__20170__D (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__20172__A1 (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA__20172__A2 (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__20173__A (.DIODE(net276));
 sky130_fd_sc_hd__diode_2 ANTENNA__20173__B (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__20178__B (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__20178__C (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__20178__D (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA__20179__A1_N (.DIODE(net281));
 sky130_fd_sc_hd__diode_2 ANTENNA__20179__A2_N (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__20179__B1 (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__20189__A1 (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__20189__A2 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__20189__B2 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__20190__A1 (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__20190__A2 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__20190__B1 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__20190__B2 (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__20191__A (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__20191__B (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__20191__C (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__20191__D (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__20192__A1_N (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__20192__A2_N (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__20193__C (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__20193__D (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__20229__A (.DIODE(_03049_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20230__A2 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__20230__B1 (.DIODE(_06837_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20230__B2 (.DIODE(_03052_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20241__A1 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__20241__A2 (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__20241__B2 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__20242__A (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__20242__B (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__20242__C (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__20243__A1 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__20243__A2 (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__20244__A (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__20244__B (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__20246__A1 (.DIODE(\mul1.b[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__20246__A2 (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__20246__B1 (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__20246__B2 (.DIODE(\mul1.b[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__20247__A (.DIODE(\mul1.b[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__20247__B (.DIODE(\mul1.b[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__20247__C (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__20247__D (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__20249__A (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__20249__B (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA__20264__A1 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA__20264__A2 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__20264__B1 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__20264__B2 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__20265__A (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__20265__B (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA__20265__C (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__20265__D (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__20266__A1 (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA__20266__A2 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__20267__A (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA__20267__B (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__20269__A1 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__20269__A2 (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA__20269__B1 (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA__20269__B2 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__20270__A (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__20270__B (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__20270__C (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA__20270__D (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA__20272__A2 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__20273__B (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__20283__A1 (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__20283__A2 (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__20283__B1 (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__20283__B2 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__20285__A (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__20285__B (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__20285__C (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__20285__D (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__20286__A1_N (.DIODE(\mul1.b[17] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__20286__A2_N (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA__20287__B (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA__20287__C (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__20308__A1 (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__20308__B2 (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA__20309__A (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__20309__B (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA__20311__A1 (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA__20312__A (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA__20317__A_N (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA__20317__B (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__20317__C (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__20317__D (.DIODE(net276));
 sky130_fd_sc_hd__diode_2 ANTENNA__20319__A1_N (.DIODE(net276));
 sky130_fd_sc_hd__diode_2 ANTENNA__20319__A2_N (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__20319__B1 (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__20319__B2 (.DIODE(net281));
 sky130_fd_sc_hd__diode_2 ANTENNA__20331__A1 (.DIODE(net628));
 sky130_fd_sc_hd__diode_2 ANTENNA__20331__A2 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__20331__B1 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__20331__B2 (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__20333__A (.DIODE(net628));
 sky130_fd_sc_hd__diode_2 ANTENNA__20333__B (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__20333__C (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__20333__D (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__20334__A1_N (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__20334__A2_N (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__20335__B (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__20335__C (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__20377__A (.DIODE(_03049_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20378__A2 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__20378__B1 (.DIODE(_06977_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20378__B2 (.DIODE(_03052_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20387__A1 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__20387__A2 (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__20387__B1 (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__20387__B2 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__20388__A (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__20388__B (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__20388__C (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__20388__D (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__20389__A1 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__20389__A2 (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__20390__A (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__20390__B (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__20392__A1 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__20392__A2 (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA__20393__A (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__20393__B (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA__20394__A (.DIODE(\mul1.b[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__20394__B (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__20394__C (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__20395__A1 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__20395__A2 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__20395__B1 (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__20410__A1 (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__20410__A2 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__20410__B1 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__20410__B2 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA__20411__A (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA__20411__B (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__20411__C (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__20411__D (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__20412__A1 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__20412__A2 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__20413__A (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__20413__B (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__20415__A1 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__20415__A2 (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA__20415__B1 (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA__20415__B2 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__20416__A (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__20416__B (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__20416__C (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA__20416__D (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA__20418__A1 (.DIODE(\mul1.b[20] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__20418__A2 (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA__20419__A (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__20419__B (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 ANTENNA__20429__A1 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__20429__A2 (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__20429__B1 (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__20429__B2 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__20431__A (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__20431__B (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__20431__C (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__20431__D (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__20432__A1_N (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__20432__A2_N (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__20433__B (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA__20433__C (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__20454__A1 (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__20454__B2 (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__20455__A (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__20455__B (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__20457__A1 (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA__20458__A (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA__20462__A_N (.DIODE(net277));
 sky130_fd_sc_hd__diode_2 ANTENNA__20462__B (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__20462__C (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__20462__D (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA__20463__A1_N (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA__20463__A2_N (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__20463__B1 (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__20463__B2 (.DIODE(net277));
 sky130_fd_sc_hd__diode_2 ANTENNA__20474__A1 (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA__20474__A2 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__20474__B1 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__20474__B2 (.DIODE(net628));
 sky130_fd_sc_hd__diode_2 ANTENNA__20476__A (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA__20476__B (.DIODE(net628));
 sky130_fd_sc_hd__diode_2 ANTENNA__20476__C (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__20476__D (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__20477__A1_N (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__20477__A2_N (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__20478__B (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__20478__C (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__20515__A2 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__20515__B1 (.DIODE(_07105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20515__B2 (.DIODE(_03052_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20516__A1 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__20519__A1 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__20519__A2 (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__20519__B1 (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA__20519__B2 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__20520__A (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__20520__B (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__20520__C (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__20520__D (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA__20522__A1 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__20522__A2 (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__20523__A (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__20523__B (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__20525__A1 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__20525__A2 (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__20527__A1 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__20541__A1 (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 ANTENNA__20541__A2 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__20541__B1 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__20541__B2 (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__20542__A (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__20542__B (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 ANTENNA__20542__C (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__20542__D (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__20543__A1 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__20543__A2 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__20544__A (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA__20544__B (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__20546__A1 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__20546__A2 (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA__20546__B1 (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__20546__B2 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__20547__A (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__20547__B (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__20547__C (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA__20547__D (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__20549__A1 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__20549__A2 (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA__20550__A (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__20550__B (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA__20560__A1 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__20560__A2 (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__20560__B1 (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__20560__B2 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__20562__A (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__20562__B (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__20562__C (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__20562__D (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__20563__A1_N (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__20563__A2_N (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__20564__B (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__20564__C (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__20582__A1 (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__20582__B2 (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__20583__A (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__20583__B (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__20585__A1 (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__20586__A (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__20590__A_N (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA__20590__B (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__20590__C (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__20590__D (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA__20592__A1_N (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA__20592__A2_N (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__20592__B1 (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__20592__B2 (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA__20604__A1 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__20604__A2 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__20604__B1 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__20604__B2 (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA__20606__A (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA__20606__B (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__20606__C (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__20606__D (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__20607__A1_N (.DIODE(net629));
 sky130_fd_sc_hd__diode_2 ANTENNA__20607__A2_N (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__20608__B (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__20608__C (.DIODE(net629));
 sky130_fd_sc_hd__diode_2 ANTENNA__20646__A (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__20647__A2 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__20647__B2 (.DIODE(_03050_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20648__S (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__20649__A (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__20650__A (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__20652__A1 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__20652__B1 (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__20652__B2 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__20653__A (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__20653__B (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__20653__D (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__20655__A (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__20655__B (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__20668__A1 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__20668__A2 (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA__20668__B1 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__20668__B2 (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 ANTENNA__20669__A (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 ANTENNA__20669__B (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__20669__C (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA__20669__D (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__20670__A1 (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__20670__A2 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__20671__A (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__20671__B (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__20673__A1 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__20673__A2 (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__20673__B1 (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__20673__B2 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__20674__A (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__20674__B (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__20674__C (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__20674__D (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__20676__A1 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__20676__A2 (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA__20677__A (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__20677__B (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA__20687__A1 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__20687__A2 (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__20687__B1 (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__20687__B2 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__20689__A (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__20689__B (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__20689__C (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__20689__D (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__20690__A1_N (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__20690__A2_N (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__20691__B (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__20691__C (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__20713__A1 (.DIODE(net628));
 sky130_fd_sc_hd__diode_2 ANTENNA__20713__B2 (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__20714__A (.DIODE(net628));
 sky130_fd_sc_hd__diode_2 ANTENNA__20714__B (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__20716__A1 (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__20717__A (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__20721__A_N (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA__20721__B (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__20721__C (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__20721__D (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__20722__A1_N (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__20722__A2_N (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__20722__B1 (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__20722__B2 (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA__20731__A1 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__20731__A2 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__20731__B1 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__20731__B2 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__20733__A (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__20733__B (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__20733__C (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__20733__D (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__20734__A1_N (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA__20734__A2_N (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__20735__B (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__20735__C (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA__20770__B (.DIODE(_03049_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20770__C (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__20771__A1 (.DIODE(_03052_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20771__A2 (.DIODE(_07365_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20771__B2 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__20772__S (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__20774__A (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__20774__B (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__20774__C (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__20775__A1 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__20775__A2 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__20775__B1 (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__20777__A (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__20777__B (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA__20791__A1 (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA__20791__A2 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__20791__B1 (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA__20791__B2 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__20792__A (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__20792__B (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA__20792__C (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__20792__D (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA__20793__A1 (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 ANTENNA__20793__A2 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__20794__A (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 ANTENNA__20794__B (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__20796__A1 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__20796__A2 (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__20796__B1 (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__20796__B2 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__20797__A (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__20797__B (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__20797__C (.DIODE(\mul1.a[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__20797__D (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__20799__A1 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__20799__A2 (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__20800__A (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__20800__B (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__20809__A1 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__20810__A1 (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__20810__A2 (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__20810__B2 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__20812__A (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__20812__B (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__20812__C (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__20813__A1_N (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__20813__A2_N (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__20814__B (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__20814__C (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__20837__A1 (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA__20837__B2 (.DIODE(net628));
 sky130_fd_sc_hd__diode_2 ANTENNA__20838__A (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA__20838__B (.DIODE(net628));
 sky130_fd_sc_hd__diode_2 ANTENNA__20838__C (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__20838__D (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__20840__A1 (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__20841__A (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__20841__B (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__20845__A_N (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__20845__B (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__20845__C (.DIODE(\mul1.b[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__20845__D (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__20847__A1_N (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__20847__A2_N (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__20847__B1 (.DIODE(_02568_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20847__B2 (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__20859__A1 (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__20859__A2 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__20859__B1 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__20859__B2 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__20861__A (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__20861__B (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__20861__C (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__20861__D (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__20862__A1_N (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__20862__A2_N (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__20863__B (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__20863__C (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__20907__A (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__20908__A2 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__20908__B2 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__20909__S (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__20910__A (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__20910__B (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__20921__A1 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__20921__A2 (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA__20921__B1 (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__20921__B2 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__20922__A (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__20922__B (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__20922__C (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA__20922__D (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__20923__A1 (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA__20923__A2 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__20924__A (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA__20924__B (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__20926__A1 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__20926__A2 (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__20926__B1 (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__20926__B2 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__20927__A (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__20927__B (.DIODE(\mul1.b[19] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__20927__C (.DIODE(\mul1.a[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__20927__D (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__20929__A1 (.DIODE(\mul1.b[20] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__20929__A2 (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__20930__A (.DIODE(\mul1.b[20] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__20930__B (.DIODE(\mul1.a[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__20939__A1 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__20939__A2 (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA__20940__A1 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__20940__B2 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__20941__A (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__20941__B (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__20943__A1 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__20943__A2 (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__20944__A (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__20944__B (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__20965__A1 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__20965__B2 (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA__20966__A (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA__20966__B (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__20968__A1 (.DIODE(net628));
 sky130_fd_sc_hd__diode_2 ANTENNA__20969__A (.DIODE(net629));
 sky130_fd_sc_hd__diode_2 ANTENNA__20975__A_N (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__20975__B (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__20975__C (.DIODE(\mul1.b[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__20975__D (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__20976__A1_N (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__20976__A2_N (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__20976__B1 (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__20976__B2 (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__20987__A1 (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 ANTENNA__20987__A2 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__20987__B1 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__20987__B2 (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__20989__A (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__20989__B (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 ANTENNA__20989__C (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__20989__D (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__20990__A1_N (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA__20990__A2_N (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__20991__B (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__20991__C (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__21028__A (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__21029__A2 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__21029__B2 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__21036__A1 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__21036__A2 (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA__21036__B1 (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__21036__B2 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__21037__A (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__21037__B (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__21037__C (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA__21037__D (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__21039__A1 (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA__21039__A2 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__21040__A (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA__21040__B (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__21042__A1 (.DIODE(\mul1.b[19] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__21042__A2 (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__21042__B2 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__21043__A (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__21043__B (.DIODE(\mul1.b[19] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__21043__C (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__21045__A1 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__21045__A2 (.DIODE(\mul1.a[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__21046__A (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__21046__B (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__21056__A (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__21056__B (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__21057__A1 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__21057__A2 (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA__21058__A (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__21058__B (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA__21060__A (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__21079__A1 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA__21079__B2 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__21080__A (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__21080__B (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA__21082__A1 (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA__21083__A (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA__21087__A_N (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__21087__B (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__21087__C (.DIODE(\mul1.b[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__21087__D (.DIODE(net629));
 sky130_fd_sc_hd__diode_2 ANTENNA__21088__A1_N (.DIODE(net629));
 sky130_fd_sc_hd__diode_2 ANTENNA__21088__A2_N (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__21088__B1 (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__21088__B2 (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__21098__A1 (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__21098__A2 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__21098__B1 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__21098__B2 (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 ANTENNA__21099__A (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 ANTENNA__21099__B (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__21099__C (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__21099__D (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__21101__A1 (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__21101__A2 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__21102__A (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__21102__B (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__21142__A (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__21143__A2 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__21143__B2 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__21150__A1 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__21150__A2 (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__21150__B1 (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__21150__B2 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__21151__A (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__21151__B (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__21151__C (.DIODE(\mul1.a[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__21152__A1 (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__21153__A (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__21153__B (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__21155__A1 (.DIODE(\mul1.b[19] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__21155__A2 (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__21155__B1 (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__21155__B2 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__21156__A (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__21156__B (.DIODE(\mul1.b[19] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__21156__C (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__21157__A1 (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__21158__A (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__21158__B (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__21167__A1 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__21167__A2 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__21167__B1 (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__21169__A (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__21170__A1 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__21170__A2 (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA__21171__A (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__21171__B (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA__21189__A1 (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__21189__B2 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA__21190__A (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA__21190__B (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__21192__A (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__21198__A1 (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA__21198__A2 (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__21198__B1 (.DIODE(\mul1.b[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__21199__A (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA__21199__C (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__21199__D (.DIODE(\mul1.b[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__21210__A1 (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA__21210__A2 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__21210__B1 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__21210__B2 (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__21211__A (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__21211__B (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA__21211__C (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__21211__D (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__21213__A (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 ANTENNA__21213__B (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__21249__A1 (.DIODE(_03052_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21249__B1 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__21250__A1 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__21252__A2 (.DIODE(_03056_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21256__A (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__21256__B (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__21258__A (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__21258__B (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__21261__A (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA__21261__B (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__21264__A (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__21264__B (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__21267__A (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__21273__A1 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__21273__A2 (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__21273__B2 (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__21278__A (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__21278__B (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__21283__A (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA__21283__B (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__21286__A (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 ANTENNA__21288__A1 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__21288__A2 (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA__21288__B2 (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__21289__A1 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__21291__A (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA__21293__A (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__21293__B (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__21296__A (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__21301__A (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__21301__B (.DIODE(\mul1.a[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__21304__A1 (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 ANTENNA__21304__A2 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__21305__A (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA__21305__B (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__21311__A (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__21311__B (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__21314__C1 (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__21314__D1 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__21315__A1 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__21315__A2 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__21315__C1 (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__21325__A1 (.DIODE(_03052_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21325__B1 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__21326__A1 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__21328__A2 (.DIODE(_03056_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21329__A1 (.DIODE(net595));
 sky130_fd_sc_hd__diode_2 ANTENNA__21329__A2 (.DIODE(net592));
 sky130_fd_sc_hd__diode_2 ANTENNA__21329__B1 (.DIODE(net645));
 sky130_fd_sc_hd__diode_2 ANTENNA__21330__A1 (.DIODE(net597));
 sky130_fd_sc_hd__diode_2 ANTENNA__21330__A2 (.DIODE(net592));
 sky130_fd_sc_hd__diode_2 ANTENNA__21330__B1 (.DIODE(net638));
 sky130_fd_sc_hd__diode_2 ANTENNA__21331__A (.DIODE(net597));
 sky130_fd_sc_hd__diode_2 ANTENNA__21331__B (.DIODE(_08642_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21332__A1 (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__21332__A2 (.DIODE(_03792_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21332__B1 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__21333__A2 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__21334__A (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__21334__B (.DIODE(_08741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21335__A1 (.DIODE(net597));
 sky130_fd_sc_hd__diode_2 ANTENNA__21335__A2 (.DIODE(_03893_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21335__B1 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__21336__A2 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__21337__A (.DIODE(net597));
 sky130_fd_sc_hd__diode_2 ANTENNA__21337__B (.DIODE(_08843_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21338__A1 (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__21338__A2 (.DIODE(_03993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21338__B1 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__21339__A2 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__21340__A (.DIODE(net597));
 sky130_fd_sc_hd__diode_2 ANTENNA__21340__B (.DIODE(_04100_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21341__A1 (.DIODE(net597));
 sky130_fd_sc_hd__diode_2 ANTENNA__21341__A2 (.DIODE(_08952_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21341__B1 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__21342__A2 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__21343__A (.DIODE(net597));
 sky130_fd_sc_hd__diode_2 ANTENNA__21343__B (.DIODE(_04209_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21344__A1 (.DIODE(net597));
 sky130_fd_sc_hd__diode_2 ANTENNA__21344__A2 (.DIODE(_09062_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21344__B1 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__21345__A2 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__21346__A (.DIODE(net597));
 sky130_fd_sc_hd__diode_2 ANTENNA__21346__B (.DIODE(_09176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21347__A1 (.DIODE(net597));
 sky130_fd_sc_hd__diode_2 ANTENNA__21347__A2 (.DIODE(_04325_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21347__B1 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__21348__A2 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__21349__A (.DIODE(net597));
 sky130_fd_sc_hd__diode_2 ANTENNA__21349__B (.DIODE(_09297_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21350__A1 (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__21350__A2 (.DIODE(_04449_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21352__A (.DIODE(net595));
 sky130_fd_sc_hd__diode_2 ANTENNA__21352__B (.DIODE(_04588_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21353__A1 (.DIODE(net595));
 sky130_fd_sc_hd__diode_2 ANTENNA__21353__A2 (.DIODE(_09434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21353__B1 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__21354__A2 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__21355__A (.DIODE(net596));
 sky130_fd_sc_hd__diode_2 ANTENNA__21355__B (.DIODE(_04719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21356__A1 (.DIODE(net596));
 sky130_fd_sc_hd__diode_2 ANTENNA__21356__A2 (.DIODE(_09564_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21357__A2 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__21358__A (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__21358__B (.DIODE(_09707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21359__A1 (.DIODE(net595));
 sky130_fd_sc_hd__diode_2 ANTENNA__21359__A2 (.DIODE(_04862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21359__B1 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__21360__A2 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__21361__A (.DIODE(net595));
 sky130_fd_sc_hd__diode_2 ANTENNA__21361__B (.DIODE(_05006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21362__A1 (.DIODE(net595));
 sky130_fd_sc_hd__diode_2 ANTENNA__21362__A2 (.DIODE(_09851_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21362__B1 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__21363__A2 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__21364__A (.DIODE(net595));
 sky130_fd_sc_hd__diode_2 ANTENNA__21364__B (.DIODE(_05156_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21365__A1 (.DIODE(net595));
 sky130_fd_sc_hd__diode_2 ANTENNA__21365__A2 (.DIODE(_09997_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21365__B1 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__21366__A2 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__21367__A (.DIODE(net596));
 sky130_fd_sc_hd__diode_2 ANTENNA__21367__B (.DIODE(_10147_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21368__A1 (.DIODE(net595));
 sky130_fd_sc_hd__diode_2 ANTENNA__21368__A2 (.DIODE(_05305_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21368__B1 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__21369__A2 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__21370__A1 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__21370__A2 (.DIODE(_05457_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21370__B1 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__21371__A1 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__21371__A2 (.DIODE(_10299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21372__A2 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__21373__A (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__21373__B (.DIODE(_10458_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21374__A1 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__21374__A2 (.DIODE(_05615_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21375__A2 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__21376__A0 (.DIODE(_05784_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21376__A1 (.DIODE(_10625_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21376__S (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__21378__B (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__21379__A0 (.DIODE(_05935_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21379__A1 (.DIODE(_10777_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21379__S (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__21380__A1 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__21381__B (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__21382__A0 (.DIODE(_06090_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21382__A1 (.DIODE(_00660_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21382__S (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__21383__A1 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__21384__A (.DIODE(net596));
 sky130_fd_sc_hd__diode_2 ANTENNA__21384__B (.DIODE(_00818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21385__A1 (.DIODE(net596));
 sky130_fd_sc_hd__diode_2 ANTENNA__21385__A2 (.DIODE(_06244_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21385__B1 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__21386__A2 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__21387__A (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__21388__A1 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__21388__A2 (.DIODE(_06402_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21389__A2 (.DIODE(_02499_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21390__B (.DIODE(_02499_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21391__A0 (.DIODE(_06552_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21391__S (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__21392__A1 (.DIODE(_02499_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21393__A (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__21394__A1 (.DIODE(net596));
 sky130_fd_sc_hd__diode_2 ANTENNA__21394__A2 (.DIODE(_06691_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21394__B1 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__21395__A2 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__21396__A (.DIODE(net596));
 sky130_fd_sc_hd__diode_2 ANTENNA__21397__A1 (.DIODE(net596));
 sky130_fd_sc_hd__diode_2 ANTENNA__21397__A2 (.DIODE(_06837_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21399__A (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__21399__B (.DIODE(_06977_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21400__A1 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__21400__B1 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__21401__A2 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__21402__A0 (.DIODE(_07105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21402__S (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__21404__A (.DIODE(net595));
 sky130_fd_sc_hd__diode_2 ANTENNA__21405__A1 (.DIODE(net596));
 sky130_fd_sc_hd__diode_2 ANTENNA__21405__B1 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__21406__A2 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__21407__A0 (.DIODE(_07365_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21407__S (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__21408__S (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__21409__A (.DIODE(net595));
 sky130_fd_sc_hd__diode_2 ANTENNA__21410__A1 (.DIODE(net595));
 sky130_fd_sc_hd__diode_2 ANTENNA__21410__B1 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__21411__A2 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__21412__A (.DIODE(net595));
 sky130_fd_sc_hd__diode_2 ANTENNA__21413__A1 (.DIODE(net596));
 sky130_fd_sc_hd__diode_2 ANTENNA__21413__B1 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__21414__A2 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__21415__A (.DIODE(net596));
 sky130_fd_sc_hd__diode_2 ANTENNA__21416__A1 (.DIODE(net595));
 sky130_fd_sc_hd__diode_2 ANTENNA__21416__B1 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__21417__A2 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__21418__S (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__21419__S (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__21420__S (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__21421__S (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__21422__A (.DIODE(net646));
 sky130_fd_sc_hd__diode_2 ANTENNA__21443__S (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__21490__S (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__21519__A0 (.DIODE(net880));
 sky130_fd_sc_hd__diode_2 ANTENNA__21520__A0 (.DIODE(net904));
 sky130_fd_sc_hd__diode_2 ANTENNA__21521__A0 (.DIODE(net885));
 sky130_fd_sc_hd__diode_2 ANTENNA__21522__A0 (.DIODE(net902));
 sky130_fd_sc_hd__diode_2 ANTENNA__21523__A0 (.DIODE(net936));
 sky130_fd_sc_hd__diode_2 ANTENNA__21524__A0 (.DIODE(net893));
 sky130_fd_sc_hd__diode_2 ANTENNA__21525__A0 (.DIODE(net921));
 sky130_fd_sc_hd__diode_2 ANTENNA__21526__A0 (.DIODE(net955));
 sky130_fd_sc_hd__diode_2 ANTENNA__21527__A0 (.DIODE(net932));
 sky130_fd_sc_hd__diode_2 ANTENNA__21528__A0 (.DIODE(net916));
 sky130_fd_sc_hd__diode_2 ANTENNA__21529__A0 (.DIODE(net945));
 sky130_fd_sc_hd__diode_2 ANTENNA__21530__A0 (.DIODE(net934));
 sky130_fd_sc_hd__diode_2 ANTENNA__21531__A0 (.DIODE(net920));
 sky130_fd_sc_hd__diode_2 ANTENNA__21532__A0 (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA__21533__A0 (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA__21534__A0 (.DIODE(net914));
 sky130_fd_sc_hd__diode_2 ANTENNA__21535__A0 (.DIODE(net923));
 sky130_fd_sc_hd__diode_2 ANTENNA__21536__A0 (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA__21569__A1 (.DIODE(_02738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21570__A1 (.DIODE(_02739_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21571__A1 (.DIODE(_02741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21572__A1 (.DIODE(_02743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21573__A1 (.DIODE(_02744_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21574__A1 (.DIODE(_02745_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21575__A1 (.DIODE(_02746_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21576__A1 (.DIODE(_02747_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21577__A1 (.DIODE(_02748_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21578__A1 (.DIODE(_02749_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21579__A1 (.DIODE(_02751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21581__RESET_B (.DIODE(net638));
 sky130_fd_sc_hd__diode_2 ANTENNA__21619__RESET_B (.DIODE(net644));
 sky130_fd_sc_hd__diode_2 ANTENNA__21621__RESET_B (.DIODE(net644));
 sky130_fd_sc_hd__diode_2 ANTENNA__21622__RESET_B (.DIODE(net644));
 sky130_fd_sc_hd__diode_2 ANTENNA__21623__RESET_B (.DIODE(net644));
 sky130_fd_sc_hd__diode_2 ANTENNA__21624__RESET_B (.DIODE(net644));
 sky130_fd_sc_hd__diode_2 ANTENNA__21625__RESET_B (.DIODE(net644));
 sky130_fd_sc_hd__diode_2 ANTENNA__21626__RESET_B (.DIODE(net644));
 sky130_fd_sc_hd__diode_2 ANTENNA__21627__RESET_B (.DIODE(net644));
 sky130_fd_sc_hd__diode_2 ANTENNA__21628__RESET_B (.DIODE(net644));
 sky130_fd_sc_hd__diode_2 ANTENNA__21629__RESET_B (.DIODE(net644));
 sky130_fd_sc_hd__diode_2 ANTENNA__21630__RESET_B (.DIODE(net644));
 sky130_fd_sc_hd__diode_2 ANTENNA__21631__RESET_B (.DIODE(net644));
 sky130_fd_sc_hd__diode_2 ANTENNA__21632__RESET_B (.DIODE(net644));
 sky130_fd_sc_hd__diode_2 ANTENNA__21633__RESET_B (.DIODE(net644));
 sky130_fd_sc_hd__diode_2 ANTENNA__21634__RESET_B (.DIODE(net644));
 sky130_fd_sc_hd__diode_2 ANTENNA__21651__RESET_B (.DIODE(net646));
 sky130_fd_sc_hd__diode_2 ANTENNA__21716__SET_B (.DIODE(net645));
 sky130_fd_sc_hd__diode_2 ANTENNA__21718__D (.DIODE(net587));
 sky130_fd_sc_hd__diode_2 ANTENNA__21718__RESET_B (.DIODE(net646));
 sky130_fd_sc_hd__diode_2 ANTENNA__21719__RESET_B (.DIODE(net646));
 sky130_fd_sc_hd__diode_2 ANTENNA__21720__D (.DIODE(net596));
 sky130_fd_sc_hd__diode_2 ANTENNA__21721__D (.DIODE(_00000_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21721__RESET_B (.DIODE(net646));
 sky130_fd_sc_hd__diode_2 ANTENNA__21722__RESET_B (.DIODE(net644));
 sky130_fd_sc_hd__diode_2 ANTENNA__21723__D (.DIODE(net610));
 sky130_fd_sc_hd__diode_2 ANTENNA__21723__RESET_B (.DIODE(net639));
 sky130_fd_sc_hd__diode_2 ANTENNA__21724__D (.DIODE(net601));
 sky130_fd_sc_hd__diode_2 ANTENNA__21724__RESET_B (.DIODE(net646));
 sky130_fd_sc_hd__diode_2 ANTENNA__21725__D (.DIODE(net599));
 sky130_fd_sc_hd__diode_2 ANTENNA__21725__RESET_B (.DIODE(net645));
 sky130_fd_sc_hd__diode_2 ANTENNA__21776__CLK (.DIODE(clknet_2_0__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__21806__CLK (.DIODE(clknet_2_1__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__21822__CLK (.DIODE(clknet_2_0__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__22064__RESET_B (.DIODE(net639));
 sky130_fd_sc_hd__diode_2 ANTENNA__22065__RESET_B (.DIODE(net639));
 sky130_fd_sc_hd__diode_2 ANTENNA__22066__RESET_B (.DIODE(net639));
 sky130_fd_sc_hd__diode_2 ANTENNA__22067__RESET_B (.DIODE(net639));
 sky130_fd_sc_hd__diode_2 ANTENNA__22068__RESET_B (.DIODE(net639));
 sky130_fd_sc_hd__diode_2 ANTENNA__22069__RESET_B (.DIODE(net639));
 sky130_fd_sc_hd__diode_2 ANTENNA__22070__RESET_B (.DIODE(net639));
 sky130_fd_sc_hd__diode_2 ANTENNA__22071__RESET_B (.DIODE(net639));
 sky130_fd_sc_hd__diode_2 ANTENNA__22072__RESET_B (.DIODE(net639));
 sky130_fd_sc_hd__diode_2 ANTENNA__22073__RESET_B (.DIODE(net639));
 sky130_fd_sc_hd__diode_2 ANTENNA__22074__RESET_B (.DIODE(net639));
 sky130_fd_sc_hd__diode_2 ANTENNA__22092__RESET_B (.DIODE(net638));
 sky130_fd_sc_hd__diode_2 ANTENNA__22102__RESET_B (.DIODE(net638));
 sky130_fd_sc_hd__diode_2 ANTENNA__22105__RESET_B (.DIODE(net638));
 sky130_fd_sc_hd__diode_2 ANTENNA__22106__RESET_B (.DIODE(net638));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_0__f_clk_i_A (.DIODE(clknet_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_1__f_clk_i_A (.DIODE(clknet_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_2__f_clk_i_A (.DIODE(clknet_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_3__f_clk_i_A (.DIODE(clknet_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_0_clk_i_A (.DIODE(clknet_2_0__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_10_clk_i_A (.DIODE(clknet_2_1__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_11_clk_i_A (.DIODE(clknet_2_1__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_12_clk_i_A (.DIODE(clknet_2_1__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_13_clk_i_A (.DIODE(clknet_2_1__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_14_clk_i_A (.DIODE(clknet_2_1__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_15_clk_i_A (.DIODE(clknet_2_1__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_16_clk_i_A (.DIODE(clknet_2_3__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_17_clk_i_A (.DIODE(clknet_2_3__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_18_clk_i_A (.DIODE(clknet_2_3__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_19_clk_i_A (.DIODE(clknet_2_3__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_1_clk_i_A (.DIODE(clknet_2_0__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_20_clk_i_A (.DIODE(clknet_2_3__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_21_clk_i_A (.DIODE(clknet_2_3__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_22_clk_i_A (.DIODE(clknet_2_3__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_23_clk_i_A (.DIODE(clknet_2_3__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_24_clk_i_A (.DIODE(clknet_2_3__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_25_clk_i_A (.DIODE(clknet_2_3__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_26_clk_i_A (.DIODE(clknet_2_3__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_27_clk_i_A (.DIODE(clknet_2_3__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_28_clk_i_A (.DIODE(clknet_2_2__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_29_clk_i_A (.DIODE(clknet_2_2__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_2_clk_i_A (.DIODE(clknet_2_0__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_30_clk_i_A (.DIODE(clknet_2_3__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_31_clk_i_A (.DIODE(clknet_2_2__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_32_clk_i_A (.DIODE(clknet_2_2__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_33_clk_i_A (.DIODE(clknet_2_2__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_34_clk_i_A (.DIODE(clknet_2_2__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_35_clk_i_A (.DIODE(clknet_2_2__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_36_clk_i_A (.DIODE(clknet_2_2__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_37_clk_i_A (.DIODE(clknet_2_2__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_38_clk_i_A (.DIODE(clknet_2_2__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_3_clk_i_A (.DIODE(clknet_2_0__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_40_clk_i_A (.DIODE(clknet_2_0__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_41_clk_i_A (.DIODE(clknet_2_0__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_43_clk_i_A (.DIODE(clknet_2_0__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_44_clk_i_A (.DIODE(clknet_2_0__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_4_clk_i_A (.DIODE(clknet_2_1__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_5_clk_i_A (.DIODE(clknet_2_1__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_6_clk_i_A (.DIODE(clknet_2_1__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_7_clk_i_A (.DIODE(clknet_2_1__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_9_clk_i_A (.DIODE(clknet_2_1__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout100_A (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout101_A (.DIODE(\mul1.b[20] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout102_A (.DIODE(\mul1.b[19] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout103_A (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout104_A (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout105_A (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout106_A (.DIODE(\mul1.b[19] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout107_A (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout108_A (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout109_A (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout10_A (.DIODE(_03050_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout110_A (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout111_A (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout113_A (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout114_A (.DIODE(\mul1.b[17] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout115_A (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout116_A (.DIODE(\mul1.b[17] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout117_A (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout118_A (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout119_A (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout11_A (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout120_A (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout122_A (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout123_A (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout124_A (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout125_A (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout127_A (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout129_A (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout12_A (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout131_A (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout132_A (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout133_A (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout134_A (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout136_A (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout138_A (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout139_A (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout141_A (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout142_A (.DIODE(\mul1.b[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout143_A (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout144_A (.DIODE(\mul1.b[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout146_A (.DIODE(\mul1.b[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout147_A (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout148_A (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout149_A (.DIODE(\mul1.b[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout14_A (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout151_A (.DIODE(\mul1.b[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout152_A (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout153_A (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout154_A (.DIODE(\mul1.b[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout155_A (.DIODE(\mul1.b[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout156_A (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout157_A (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout158_A (.DIODE(\mul1.b[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout159_A (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout15_A (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout160_A (.DIODE(\mul1.b[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout161_A (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout162_A (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout163_A (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout164_A (.DIODE(\mul1.b[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout165_A (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout166_A (.DIODE(\mul1.b[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout167_A (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout168_A (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout169_A (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout170_A (.DIODE(\mul1.b[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout171_A (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout172_A (.DIODE(\mul1.b[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout173_A (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout174_A (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout175_A (.DIODE(\mul1.b[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout176_A (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout177_A (.DIODE(\mul1.b[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout178_A (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout179_A (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout17_A (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout180_A (.DIODE(\mul1.b[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout182_A (.DIODE(\mul1.b[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout183_A (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout184_A (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout185_A (.DIODE(\mul1.b[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout186_A (.DIODE(\mul1.b[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout187_A (.DIODE(\mul1.b[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout188_A (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout189_A (.DIODE(\mul1.b[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout18_A (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout191_A (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout192_A (.DIODE(\mul1.b[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout193_A (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout195_A (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout197_A (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout199_A (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout19_A (.DIODE(_02823_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1_A (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout200_A (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout202_A (.DIODE(\mul1.a[27] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout203_A (.DIODE(\mul1.a[27] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout204_A (.DIODE(\mul1.a[27] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout205_A (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout206_A (.DIODE(\mul1.a[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout207_A (.DIODE(\mul1.a[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout208_A (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout209_A (.DIODE(\mul1.a[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout20_A (.DIODE(_02823_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout210_A (.DIODE(\mul1.a[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout211_A (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout212_A (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout213_A (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout215_A (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout216_A (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout217_A (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout219_A (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout21_A (.DIODE(_02823_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout220_A (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout221_A (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout222_A (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout224_A (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout225_A (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout226_A (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout228_A (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout22_A (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout231_A (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout233_A (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout234_A (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout236_A (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout238_A (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout239_A (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout23_A (.DIODE(_02757_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout241_A (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout243_A (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout244_A (.DIODE(\mul1.a[17] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout245_A (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout246_A (.DIODE(\mul1.a[17] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout247_A (.DIODE(\mul1.a[17] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout248_A (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout249_A (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout24_A (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout250_A (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout251_A (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout253_A (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout254_A (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout255_A (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout256_A (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout258_A (.DIODE(\mul1.a[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout259_A (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout25_A (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout260_A (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout261_A (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout262_A (.DIODE(\mul1.a[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout263_A (.DIODE(\mul1.a[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout264_A (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout265_A (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout266_A (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout267_A (.DIODE(\mul1.a[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout268_A (.DIODE(net272));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout269_A (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout26_A (.DIODE(_02756_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout270_A (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout271_A (.DIODE(net272));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout273_A (.DIODE(\mul1.a[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout274_A (.DIODE(\mul1.a[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout275_A (.DIODE(net276));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout276_A (.DIODE(net277));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout277_A (.DIODE(\mul1.a[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout278_A (.DIODE(\mul1.a[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout279_A (.DIODE(\mul1.a[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout27_A (.DIODE(_02756_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout280_A (.DIODE(net281));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout281_A (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout282_A (.DIODE(\mul1.a[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout283_A (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout284_A (.DIODE(\mul1.a[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout285_A (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout286_A (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout287_A (.DIODE(\mul1.a[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout288_A (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout289_A (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout28_A (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout290_A (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout291_A (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout293_A (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout294_A (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout295_A (.DIODE(\mul1.a[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout296_A (.DIODE(\mul1.a[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout297_A (.DIODE(\mul1.a[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout298_A (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout299_A (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout29_A (.DIODE(_02755_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout2_A (.DIODE(_03055_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout300_A (.DIODE(\mul1.a[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout301_A (.DIODE(\mul1.a[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout302_A (.DIODE(\mul1.a[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout303_A (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout304_A (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout305_A (.DIODE(\mul1.a[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout306_A (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout307_A (.DIODE(\mul1.a[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout308_A (.DIODE(net309));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout309_A (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout310_A (.DIODE(\mul1.a[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout311_A (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout312_A (.DIODE(\mul1.a[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout313_A (.DIODE(net314));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout314_A (.DIODE(\mul1.a[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout315_A (.DIODE(\mul1.a[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout316_A (.DIODE(net317));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout317_A (.DIODE(\mul1.a[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout318_A (.DIODE(net320));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout319_A (.DIODE(net320));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout31_A (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout320_A (.DIODE(\mul1.a[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout321_A (.DIODE(\mul1.a[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout322_A (.DIODE(net325));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout323_A (.DIODE(net325));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout324_A (.DIODE(net325));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout326_A (.DIODE(\mul0.b[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout327_A (.DIODE(net328));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout329_A (.DIODE(net330));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout330_A (.DIODE(\mul0.b[29] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout331_A (.DIODE(net332));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout332_A (.DIODE(net333));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout334_A (.DIODE(net335));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout335_A (.DIODE(net336));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout337_A (.DIODE(\mul0.b[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout338_A (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout339_A (.DIODE(\mul0.b[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout33_A (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout340_A (.DIODE(net341));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout342_A (.DIODE(net343));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout344_A (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout346_A (.DIODE(net347));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout348_A (.DIODE(\mul0.b[23] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout349_A (.DIODE(net351));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout34_A (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout350_A (.DIODE(net351));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout351_A (.DIODE(\mul0.b[23] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout352_A (.DIODE(net354));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout353_A (.DIODE(net354));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout354_A (.DIODE(net355));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout356_A (.DIODE(net360));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout357_A (.DIODE(net359));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout358_A (.DIODE(net359));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout359_A (.DIODE(net360));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout35_A (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout361_A (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout362_A (.DIODE(net363));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout363_A (.DIODE(\mul0.b[20] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout364_A (.DIODE(\mul0.b[20] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout365_A (.DIODE(\mul0.b[19] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout366_A (.DIODE(net367));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout367_A (.DIODE(net369));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout368_A (.DIODE(net369));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout369_A (.DIODE(\mul0.b[19] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout36_A (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout370_A (.DIODE(net371));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout371_A (.DIODE(\mul0.b[17] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout372_A (.DIODE(\mul0.b[17] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout373_A (.DIODE(\mul0.b[17] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout374_A (.DIODE(\mul0.b[17] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout375_A (.DIODE(net380));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout376_A (.DIODE(net380));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout377_A (.DIODE(net380));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout378_A (.DIODE(net379));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout379_A (.DIODE(net380));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout37_A (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout381_A (.DIODE(\mul0.b[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout382_A (.DIODE(\mul0.b[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout383_A (.DIODE(net385));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout384_A (.DIODE(net385));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout385_A (.DIODE(\mul0.b[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout386_A (.DIODE(net389));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout387_A (.DIODE(net389));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout388_A (.DIODE(net389));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout390_A (.DIODE(\mul0.b[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout391_A (.DIODE(\mul0.b[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout392_A (.DIODE(net394));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout393_A (.DIODE(net394));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout394_A (.DIODE(\mul0.b[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout395_A (.DIODE(net396));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout396_A (.DIODE(\mul0.b[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout399_A (.DIODE(\mul0.b[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout39_A (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout3_A (.DIODE(_03055_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout400_A (.DIODE(net401));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout401_A (.DIODE(\mul0.b[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout402_A (.DIODE(net403));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout403_A (.DIODE(\mul0.b[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout404_A (.DIODE(net405));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout405_A (.DIODE(\mul0.b[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout406_A (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout407_A (.DIODE(\mul0.b[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout408_A (.DIODE(net412));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout409_A (.DIODE(net412));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout40_A (.DIODE(_02499_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout410_A (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout411_A (.DIODE(net412));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout413_A (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout414_A (.DIODE(\mul0.b[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout415_A (.DIODE(net416));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout416_A (.DIODE(\mul0.b[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout417_A (.DIODE(net418));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout418_A (.DIODE(\mul0.b[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout419_A (.DIODE(net420));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout420_A (.DIODE(\mul0.b[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout421_A (.DIODE(net422));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout422_A (.DIODE(net425));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout423_A (.DIODE(net424));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout424_A (.DIODE(net425));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout426_A (.DIODE(net427));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout427_A (.DIODE(\mul0.b[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout428_A (.DIODE(net429));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout429_A (.DIODE(\mul0.b[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout430_A (.DIODE(net431));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout431_A (.DIODE(net432));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout432_A (.DIODE(\mul0.b[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout433_A (.DIODE(net434));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout434_A (.DIODE(\mul0.b[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout435_A (.DIODE(net436));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout436_A (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout437_A (.DIODE(\mul0.b[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout438_A (.DIODE(net439));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout439_A (.DIODE(\mul0.b[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout440_A (.DIODE(net442));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout441_A (.DIODE(net442));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout445_A (.DIODE(net446));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout446_A (.DIODE(\mul0.b[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout447_A (.DIODE(\mul0.b[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout450_A (.DIODE(net452));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout451_A (.DIODE(net452));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout453_A (.DIODE(\mul0.a[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout454_A (.DIODE(\mul0.a[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout455_A (.DIODE(net456));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout458_A (.DIODE(\mul0.a[29] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout459_A (.DIODE(\mul0.a[29] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout460_A (.DIODE(net462));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout461_A (.DIODE(net462));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout462_A (.DIODE(\mul0.a[28] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout463_A (.DIODE(\mul0.a[27] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout464_A (.DIODE(\mul0.a[27] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout465_A (.DIODE(\mul0.a[27] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout466_A (.DIODE(net469));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout467_A (.DIODE(net469));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout468_A (.DIODE(net469));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout46_A (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout470_A (.DIODE(net473));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout471_A (.DIODE(net473));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout472_A (.DIODE(net473));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout474_A (.DIODE(net477));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout475_A (.DIODE(net477));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout476_A (.DIODE(net477));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout478_A (.DIODE(net481));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout479_A (.DIODE(net481));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout47_A (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout480_A (.DIODE(net481));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout482_A (.DIODE(\mul0.a[22] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout483_A (.DIODE(\mul0.a[22] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout484_A (.DIODE(\mul0.a[22] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout485_A (.DIODE(\mul0.a[22] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout486_A (.DIODE(\mul0.a[21] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout487_A (.DIODE(\mul0.a[21] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout488_A (.DIODE(\mul0.a[21] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout489_A (.DIODE(\mul0.a[21] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout48_A (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout490_A (.DIODE(\mul0.a[20] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout491_A (.DIODE(\mul0.a[20] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout492_A (.DIODE(net493));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout493_A (.DIODE(\mul0.a[20] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout494_A (.DIODE(\mul0.a[19] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout495_A (.DIODE(\mul0.a[19] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout496_A (.DIODE(net497));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout497_A (.DIODE(\mul0.a[19] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout498_A (.DIODE(net499));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout499_A (.DIODE(\mul0.a[18] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout4_A (.DIODE(_03055_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout502_A (.DIODE(\mul0.a[18] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout503_A (.DIODE(\mul0.a[17] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout504_A (.DIODE(\mul0.a[17] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout505_A (.DIODE(net506));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout506_A (.DIODE(\mul0.a[17] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout507_A (.DIODE(net508));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout508_A (.DIODE(\mul0.a[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout509_A (.DIODE(net510));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout50_A (.DIODE(_02753_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout510_A (.DIODE(\mul0.a[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout511_A (.DIODE(net512));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout512_A (.DIODE(\mul0.a[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout513_A (.DIODE(\mul0.a[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout514_A (.DIODE(\mul0.a[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout515_A (.DIODE(net516));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout516_A (.DIODE(net517));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout517_A (.DIODE(\mul0.a[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout518_A (.DIODE(\mul0.a[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout519_A (.DIODE(\mul0.a[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout51_A (.DIODE(_02753_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout520_A (.DIODE(net521));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout521_A (.DIODE(net524));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout522_A (.DIODE(net523));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout523_A (.DIODE(net524));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout525_A (.DIODE(net527));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout526_A (.DIODE(net527));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout527_A (.DIODE(\mul0.a[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout528_A (.DIODE(net529));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout529_A (.DIODE(\mul0.a[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout531_A (.DIODE(net532));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout532_A (.DIODE(\mul0.a[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout533_A (.DIODE(\mul0.a[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout534_A (.DIODE(\mul0.a[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout535_A (.DIODE(net536));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout536_A (.DIODE(net537));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout537_A (.DIODE(net539));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout538_A (.DIODE(net539));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout540_A (.DIODE(net541));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout541_A (.DIODE(net542));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout542_A (.DIODE(\mul0.a[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout543_A (.DIODE(\mul0.a[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout544_A (.DIODE(net545));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout545_A (.DIODE(\mul0.a[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout546_A (.DIODE(\mul0.a[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout547_A (.DIODE(\mul0.a[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout548_A (.DIODE(net549));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout549_A (.DIODE(net550));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout54_A (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout550_A (.DIODE(\mul0.a[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout551_A (.DIODE(\mul0.a[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout552_A (.DIODE(net553));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout553_A (.DIODE(net554));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout554_A (.DIODE(net556));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout555_A (.DIODE(net556));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout557_A (.DIODE(net558));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout558_A (.DIODE(\mul0.a[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout559_A (.DIODE(net560));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout560_A (.DIODE(\mul0.a[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout561_A (.DIODE(net565));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout562_A (.DIODE(net563));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout563_A (.DIODE(net564));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout564_A (.DIODE(net565));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout566_A (.DIODE(net570));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout567_A (.DIODE(net570));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout568_A (.DIODE(net569));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout569_A (.DIODE(net570));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout56_A (.DIODE(_02568_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout571_A (.DIODE(net575));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout572_A (.DIODE(net575));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout573_A (.DIODE(net574));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout574_A (.DIODE(net575));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout576_A (.DIODE(\mul0.a[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout577_A (.DIODE(net580));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout578_A (.DIODE(net580));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout579_A (.DIODE(net580));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout580_A (.DIODE(\mul0.a[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout581_A (.DIODE(net582));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout582_A (.DIODE(net584));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout583_A (.DIODE(net584));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout585_A (.DIODE(net586));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout586_A (.DIODE(net587));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout587_A (.DIODE(net592));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout588_A (.DIODE(net592));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout589_A (.DIODE(net592));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout58_A (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout590_A (.DIODE(net591));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout591_A (.DIODE(net592));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout593_A (.DIODE(net598));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout594_A (.DIODE(net598));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout595_A (.DIODE(net596));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout596_A (.DIODE(net597));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout597_A (.DIODE(net598));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout599_A (.DIODE(net600));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout59_A (.DIODE(_02561_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout5_A (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout601_A (.DIODE(net606));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout602_A (.DIODE(net606));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout603_A (.DIODE(net606));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout604_A (.DIODE(net606));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout605_A (.DIODE(net606));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout607_A (.DIODE(\state[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout608_A (.DIODE(\state[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout609_A (.DIODE(\state[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout60_A (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout610_A (.DIODE(\state[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout611_A (.DIODE(\state[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout616_A (.DIODE(\state[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout617_A (.DIODE(\state[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout618_A (.DIODE(\state[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout619_A (.DIODE(\state[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout61_A (.DIODE(_02561_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout620_A (.DIODE(\state[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout621_A (.DIODE(net622));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout622_A (.DIODE(\mul1.b[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout623_A (.DIODE(net625));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout624_A (.DIODE(net625));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout625_A (.DIODE(\mul1.b[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout626_A (.DIODE(net629));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout627_A (.DIODE(net629));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout628_A (.DIODE(net629));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout629_A (.DIODE(net630));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout62_A (.DIODE(\mul1.b[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout631_A (.DIODE(\mul0.b[18] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout632_A (.DIODE(\mul0.b[18] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout633_A (.DIODE(\mul0.b[18] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout634_A (.DIODE(net635));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout635_A (.DIODE(\mul0.b[18] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout636_A (.DIODE(net638));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout637_A (.DIODE(net638));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout638_A (.DIODE(net639));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout639_A (.DIODE(net646));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout63_A (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout642_A (.DIODE(net645));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout643_A (.DIODE(net645));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout644_A (.DIODE(net645));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout645_A (.DIODE(net646));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout64_A (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout66_A (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout67_A (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout69_A (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout6_A (.DIODE(_03794_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout70_A (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout72_A (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout73_A (.DIODE(\mul1.b[27] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout74_A (.DIODE(\mul1.b[27] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout75_A (.DIODE(\mul1.b[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout76_A (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout77_A (.DIODE(\mul1.b[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout78_A (.DIODE(\mul1.b[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout79_A (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout7_A (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout80_A (.DIODE(\mul1.b[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout81_A (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout82_A (.DIODE(\mul1.b[24] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout83_A (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout84_A (.DIODE(\mul1.b[24] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout85_A (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout86_A (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout87_A (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout89_A (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout90_A (.DIODE(\mul1.b[22] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout91_A (.DIODE(\mul1.b[22] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout92_A (.DIODE(\mul1.b[22] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout93_A (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout94_A (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout95_A (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout96_A (.DIODE(\mul1.b[21] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout97_A (.DIODE(\mul1.b[21] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout98_A (.DIODE(\mul1.b[20] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout99_A (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout9_A (.DIODE(_03057_));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold234_A (.DIODE(\in_data[96] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold239_A (.DIODE(\in_data[98] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold241_A (.DIODE(\mul0.b[23] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold247_A (.DIODE(\in_data[101] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold256_A (.DIODE(\in_data[99] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold258_A (.DIODE(\in_data[97] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold262_A (.DIODE(\in_data[109] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold268_A (.DIODE(\in_data[111] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold270_A (.DIODE(\in_data[105] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold274_A (.DIODE(\in_data[108] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold275_A (.DIODE(\in_data[102] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold277_A (.DIODE(\in_data[112] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold283_A (.DIODE(\in_data[113] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold286_A (.DIODE(\in_data[104] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold288_A (.DIODE(\in_data[107] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold290_A (.DIODE(\in_data[100] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold299_A (.DIODE(\in_data[106] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold306_A (.DIODE(\in_data[110] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold309_A (.DIODE(\in_data[103] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold313_A (.DIODE(\mul0.a[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold319_A (.DIODE(\mul0.b[31] ));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_1029 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1033 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_1037 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1045 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1061 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_1073 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_1077 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_1086 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_1097 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_1101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_1110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_1114 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_1121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_1158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_1169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_1188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_1192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_1196 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_1200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_1221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_1273 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_173 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_176 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_416 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_488 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_516 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_568 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_626 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_684 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_766 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_780 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_790 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_794 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_848 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_865 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_883 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_929 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_943 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_957 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_960 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_985 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_994 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_1020 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_1041 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_1045 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_1064 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_1074 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_1078 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_1085 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_1093 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_1097 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_1109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_1123 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_1127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_1164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_1168 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_1205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_1209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_1221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_1232 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_1256 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_1270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_1276 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_235 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_244 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_295 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_370 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_392 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_396 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_619 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_642 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_690 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_699 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_921 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_945 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_962 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_997 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_1000 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_1004 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_1034 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_1038 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_1089 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_1118 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_1128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_1132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_1136 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_1141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_1152 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_1156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_1194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_1198 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1213 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_1229 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_1245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_189 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_25 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_294 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_379 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_426 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_482 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_630 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_638 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_647 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_718 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_9 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_936 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_944 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_982 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_986 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_990 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_1011 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_1015 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_1023 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_103 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_1043 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_1047 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_1079 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_1083 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_1097 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_1101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_1128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_1132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_1153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_1157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_1188 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_1192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_1200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_1229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_1254 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_1270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_1276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_171 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_207 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_211 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_548 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_630 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_638 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_652 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_672 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_690 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_821 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_824 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_840 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_864 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_893 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_905 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_920 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_985 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_994 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_1001 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_1019 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_1023 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_1080 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_1084 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_1097 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_1133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_1152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_1156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_1161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_1165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_1169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_1173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_1181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_1185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_1189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_1193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_1231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_1243 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_1268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_1276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_218 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_490 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_515 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_52 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_646 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_657 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_700 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_712 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_738 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_792 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_804 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_823 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_912 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_969 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_973 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_977 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_982 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_1003 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_1035 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_1078 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_1100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_1117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_1126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_1130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_1183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_1187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_1191 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_1221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_1225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_1244 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_1257 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_1272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_1276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_219 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_392 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_403 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_562 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_599 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_630 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_638 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_658 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_664 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_712 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_722 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_786 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_804 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_823 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_827 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_9 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_917 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_973 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_977 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_984 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_1004 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_1025 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_1029 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_1045 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_108 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_1089 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_1133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_1137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_1148 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_1180 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_1184 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_1194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_1242 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_1246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_1263 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_1273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_267 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_294 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_379 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_388 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_453 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_476 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_487 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_520 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_532 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_583 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_621 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_629 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_704 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_712 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_716 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_727 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_749 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_776 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_780 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_790 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_814 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_826 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_921 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_930 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_940 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_950 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_986 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_99 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_1022 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_1030 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_1067 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_1091 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_1104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_1113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_1117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_1125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_1129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_1165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_1175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_1205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_1232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_1242 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_1246 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_1254 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_1270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_1276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_168 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_192 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_392 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_443 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_472 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_508 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_59 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_626 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_632 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_638 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_660 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_676 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_722 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_726 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_735 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_769 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_794 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_818 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_842 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_923 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_933 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_953 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_1087 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1095 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_1119 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_1127 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_1131 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_1135 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_1141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_1153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_1157 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_1165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_1175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_1208 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_1212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_1241 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_347 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_422 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_453 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_523 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_626 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_638 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_650 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_688 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_7 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_760 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_772 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_778 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_792 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_815 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_832 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_929 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_947 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_951 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_969 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_987 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_991 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_1003 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_1042 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_1046 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_1080 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_1084 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_1088 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1173 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_1185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_1200 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_1222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_1232 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_1259 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_1270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_1276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_431 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_541 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_59 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_622 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_630 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_666 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_684 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_688 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_77 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_777 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_828 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_864 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_976 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_1007 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_1040 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_1044 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_1048 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_1052 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_1058 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_1073 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_1175 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_1183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_1228 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_1272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_1276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_135 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_254 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_350 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_453 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_650 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_681 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_720 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_764 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_776 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_791 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_806 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_818 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_966 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_990 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_1004 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_1008 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_1021 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_1025 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_1033 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_1042 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_1046 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_1052 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_1060 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_1064 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_1068 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1072 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_1084 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_1197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_1273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_155 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_219 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_238 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_375 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_492 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_513 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_640 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_658 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_675 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_734 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_775 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_779 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_789 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_802 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_806 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_829 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_849 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_891 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_894 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_899 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_910 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_915 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_932 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_936 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_940 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_95 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_960 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_968 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_976 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_984 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_988 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_1007 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_1025 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_1029 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_1041 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_1056 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1060 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1072 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_1084 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1173 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_1185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_1221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_1232 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_1259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_1270 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_1274 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_192 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_22 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_270 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_283 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_403 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_456 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_603 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_609 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_630 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_636 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_64 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_699 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_724 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_728 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_744 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_748 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_767 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_776 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_793 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_803 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_91 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_937 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_957 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_967 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_985 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_997 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_100 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_1000 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_1169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_1175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_1177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_1185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_1211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_1224 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_1228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_1237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_216 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_28 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_319 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_43 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_568 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_694 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_736 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_782 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_792 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_801 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_96 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_976 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_988 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_1203 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_1209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_1249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_1261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_1273 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_204 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_275 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_288 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_300 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_416 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_528 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_548 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_602 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_607 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_619 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_638 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_651 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_668 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_672 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_678 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_686 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_831 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_843 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_981 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1201 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_1213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_1219 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_254 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_295 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_541 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_569 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_590 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_599 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_633 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_666 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_670 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_686 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_698 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_723 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_736 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_822 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_834 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_102 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_1217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_1221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_1245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_1270 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_1274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_226 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_288 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_292 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_46 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_572 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_58 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_628 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_638 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_652 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_664 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_676 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_716 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_728 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_732 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_770 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_774 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_829 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_917 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_100 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_1169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_1241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_1252 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_182 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_267 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_406 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_581 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_639 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_661 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_680 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_700 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_710 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_735 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_760 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_803 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_807 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_819 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_945 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_1203 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_1211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_1261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_1265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_1269 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_1273 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_132 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_214 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_37 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_416 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_555 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_562 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_651 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_661 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_667 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_742 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_770 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_787 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1077 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_1275 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_173 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_179 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_320 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_324 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_734 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_778 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_819 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1217 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_1229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_1237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_1240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_1253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_1257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_1270 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_1274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_214 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_230 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_336 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_547 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_593 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_664 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_670 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_696 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_762 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_766 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_779 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_95 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_1225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_1231 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_1239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_127 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_1271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_182 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_476 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_482 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_579 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_591 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_595 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_704 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_734 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_738 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_756 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_760 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_764 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_795 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_807 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_819 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_84 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_88 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_92 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_1002 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_1035 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_1041 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_1069 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1073 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1097 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_1109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_1133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_1137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1152 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_1269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_302 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_420 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_541 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_590 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_620 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_656 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_681 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_686 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_70 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_744 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_767 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_800 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_839 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_859 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_878 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_902 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_911 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_922 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_969 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_973 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_976 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_980 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_1085 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1173 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_1203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_1205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_1213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_1242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_1252 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_1256 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_1270 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_1274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_136 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_226 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_238 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_397 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_434 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_60 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_622 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_672 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_692 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_718 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_732 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_736 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_94 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_1189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_1195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_1198 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_1211 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_1215 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_1229 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_1237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_480 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_535 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_556 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_571 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_588 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_591 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_64 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_644 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_679 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_704 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_736 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_744 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_965 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_1217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_1225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_1229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_1240 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_1250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_1256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_1270 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_1274 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_168 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_235 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_468 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_560 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_60 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_692 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_696 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_728 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_732 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_760 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_764 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_773 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_778 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_790 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_802 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_949 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1009 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_1189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_1197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_1223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_1276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_156 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_18 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_241 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_430 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_460 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_495 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_691 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_70 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_704 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_724 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_736 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_758 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_762 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_770 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_794 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_806 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_818 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1049 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_119 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_1217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_1225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_1245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_1254 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_1258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_1270 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_1274 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_145 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_294 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_336 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_518 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_556 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_58 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_602 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_640 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_708 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_763 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_788 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_795 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_80 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_1169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_1225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_1228 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_1260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_1270 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_1274 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_186 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_303 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_422 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_513 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_528 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_535 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_539 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_687 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_736 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_746 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_770 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_774 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_84 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1017 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_102 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_1252 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_1256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_1270 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_1274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_275 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_506 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_579 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_631 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_681 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_720 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_735 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_764 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_768 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_776 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_802 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1089 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_1169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1189 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_1201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_1205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_1208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_1212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_1216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_1220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_1224 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_1228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_1237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_1241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_1268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_1272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_1276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_142 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_347 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_359 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_366 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_426 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_556 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_571 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_579 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_697 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_712 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_718 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_733 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_768 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_788 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_836 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_1085 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1161 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_1203 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_1211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_1214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_1218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_1222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_1226 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_1234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_1245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_1253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_1257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_1270 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_1274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_13 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_17 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_43 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_444 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_459 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_563 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_643 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_699 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_732 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_760 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_764 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_771 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_792 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_804 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1065 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_118 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_1256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_1260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_1264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_1268 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_1272 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_28 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_434 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_458 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_508 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_532 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_554 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_606 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_647 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_734 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_738 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_742 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_767 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_1000 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_1004 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_1008 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_1012 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_1020 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_1042 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_1046 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_1066 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_1070 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_1074 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1078 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_1273 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_152 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_170 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_274 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_320 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_456 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_506 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_575 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_643 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_672 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_681 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_734 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_749 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_760 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_766 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_806 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_846 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_890 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_898 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_91 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_921 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_925 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_933 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_966 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_992 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1117 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_1197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_1200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_1214 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_1218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_1228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_1232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_1236 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_1240 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_1244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_1253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_1257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_1270 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_1274 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_152 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_175 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_23 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_434 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_472 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_485 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_570 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_602 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_7 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_770 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_784 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1089 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1213 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_1229 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_1267 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_1271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_1275 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_174 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_254 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_276 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_366 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_44 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_463 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_569 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_659 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_736 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_744 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_114 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_117 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_1173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_1178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_1189 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_1203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_1205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_1213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_1259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_1270 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_1274 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_370 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_392 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_410 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_472 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_563 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_682 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_790 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_80 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_849 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1077 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1157 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_1169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_1173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_1224 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_1228 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_1241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_1245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_1271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_1275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_204 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_263 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_28 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_288 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_415 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_492 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_529 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_61 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_644 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_648 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_709 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_732 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_977 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1073 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_108 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_114 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_1185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_1193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_1203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_1205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_1215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_1228 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_1232 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_1236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_1254 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_1258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_1270 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_1274 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_239 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_276 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_404 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_472 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_508 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_515 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_526 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_59 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_651 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_774 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_917 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_100 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_1169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1201 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_1251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_174 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_28 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_323 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_426 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_43 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_469 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_513 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_538 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_591 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_646 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_670 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_84 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_877 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_88 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_10 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1073 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_108 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1149 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_1241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_1269 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_1273 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_136_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_136_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_23 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_247 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_284 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_136_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_136_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_136_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_35 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_386 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_392 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_136_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_416 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_428 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_136_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_136_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_136_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_669 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_688 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_726 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_736 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_80 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_136_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_100 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1077 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_1269 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_151 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_288 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_310 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_399 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_462 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_579 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_590 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_663 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_682 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_689 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_717 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_739 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_764 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_77 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_776 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_889 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_1259 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_1261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_1267 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_1270 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_1274 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_192 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_370 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_400 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_416 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_434 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_450 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_459 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_506 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_572 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_698 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_722 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_728 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_736 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_790 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_1251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_1275 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_139_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_252 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_255 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_276 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_382 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_438 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_471 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_139_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_487 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_139_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_540 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_568 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_598 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_139_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_639 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_139_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_736 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_139_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_771 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_778 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1025 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_1046 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_1050 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_1069 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1073 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1097 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_1109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_184 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_196 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_350 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_458 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_532 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_668 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_736 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_744 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_759 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_76 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_794 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_838 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_851 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_873 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_946 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_990 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_994 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_1273 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_292 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_336 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_454 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_485 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_568 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_584 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_652 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_660 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_674 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_789 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_1253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_294 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_350 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_434 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_525 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_565 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_575 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_583 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_660 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_664 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_691 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_756 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_760 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_778 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_142_1273 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_142_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_201 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_142_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_142_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_142_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_312 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_316 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_142_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_142_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_396 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_426 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_438 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_142_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_520 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_142_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_574 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_586 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_619 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_677 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_728 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_778 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_790 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_1269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_327 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_438 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_442 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_570 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_579 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_639 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_687 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_702 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_707 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_726 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_739 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_144_1273 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_144_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_248 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_144_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_144_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_436 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_144_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_507 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_144_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_144_541 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_144_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_581 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_144_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_144_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_144_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_144_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_669 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_678 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_684 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_144_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_719 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_773 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_144_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_1269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_145_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_145_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_145_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_145_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_397 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_407 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_430 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_145_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_145_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_145_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_145_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_520 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_145_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_145_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_145_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_649 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_145_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_145_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_145_683 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_687 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_702 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_145_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_736 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_764 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_776 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146_1273 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_227 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_146_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_146_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_146_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146_369 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_146_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_392 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_448 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_504 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_566 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_586 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_612 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_616 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_146_624 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_146_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_653 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_668 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_1269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_351 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_147_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_435 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_147_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_512 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_147_527 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_639 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_665 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_708 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_742 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_763 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_148_1273 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_148_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_148_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_148_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_300 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_148_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_148_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_336 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_148_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_372 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_384 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_148_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_148_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_506 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_515 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_148_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_148_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_537 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_551 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_596 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_148_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_148_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_640 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_148_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_667 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_674 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_686 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_710 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_148_716 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_148_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_148_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_149_1269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_270 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_149_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_149_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_350 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_149_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_149_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_149_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_149_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_149_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_149_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_149_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_149_580 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_149_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_149_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_665 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_149_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_692 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_149_739 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_778 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_989 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_1040 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_1044 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_1048 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_1067 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_1071 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1075 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_114 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_1273 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_163 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_235 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_374 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_436 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_440 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_522 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_551 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_562 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_628 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_688 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_731 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_735 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_743 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_753 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_792 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_835 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_916 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_948 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_150_1273 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_150_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_150_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_150_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_316 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_150_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_150_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_150_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_150_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_411 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_150_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_436 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_150_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_150_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_459 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_150_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_472 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_150_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_515 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_150_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_540 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_562 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_150_618 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_150_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_678 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_150_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_150_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_711 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_734 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_1269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_260 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_151_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_151_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_360 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_364 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_151_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_434 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_151_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_151_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_151_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_522 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_151_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_151_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_628 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_638 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_648 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_708 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_152_1273 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_152_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_152_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_152_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_400 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_431 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_152_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_536 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_554 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_152_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_572 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_578 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_652 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_152_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_1269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_245 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_153_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_459 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_153_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_153_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_564 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_592 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_640 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_644 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_153_647 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_154_1273 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_154_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_154_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_154_370 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_154_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_414 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_154_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_154_482 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_154_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_627 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_154_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_154_650 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_662 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_155_1269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_155_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_155_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_344 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_155_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_155_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_155_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_155_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_478 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_155_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_155_51 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_534 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_155_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_155_566 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_570 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_583 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_155_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_606 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_629 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_647 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_650 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_654 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_989 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_1089 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_156_1273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_156_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_156_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_156_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_156_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_156_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_605 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_1004 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_1016 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_1025 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_1035 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1050 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_1072 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_1076 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_1080 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1084 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1096 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1257 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_126 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_180 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_320 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_403 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_635 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_68 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_707 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_745 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_832 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_860 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_895 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_94 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_950 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1011 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1023 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_1035 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_1037 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_1043 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_1053 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_1069 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_1273 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_168 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_338 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_409 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_450 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_510 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_526 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_59 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_652 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_656 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_668 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_676 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_685 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_699 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_743 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_754 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_845 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_899 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_917 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_938 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_950 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_976 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_985 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_1075 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_1079 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1083 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1095 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_1269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_151 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_210 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_316 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_524 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_579 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_628 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_634 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_686 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_692 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_695 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_700 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_756 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_760 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_764 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_889 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_914 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_926 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_938 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_944 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_966 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_1004 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1014 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1043 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_1073 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_1077 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_1088 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1097 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_119 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_1273 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_164 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_214 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_259 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_504 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_667 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_674 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_698 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_736 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_78 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_784 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_813 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_852 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_858 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_867 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_900 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_904 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_920 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_929 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_936 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_967 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_979 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_986 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_992 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_996 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_1007 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_1022 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_1026 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_1032 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_1043 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_1055 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_1073 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_1077 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_1081 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_1095 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_1101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_1105 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_1109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_1169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_1269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_412 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_459 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_679 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_683 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_691 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_700 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_711 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_736 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_756 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_764 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_839 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_857 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_860 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_873 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_889 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_90 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_913 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_917 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_950 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_960 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_972 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_1002 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_1006 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_1044 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_1048 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1063 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1073 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_1095 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1119 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_1145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_1172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_1195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_1199 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1215 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_1227 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_1269 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_252 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_512 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_579 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_682 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_689 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_708 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_759 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_763 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_794 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_819 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_850 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_857 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_876 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_880 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_894 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_936 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_940 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_962 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_966 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_970 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_986 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_990 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_994 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_998 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_1006 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_1012 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_1020 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_1030 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_1044 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_1055 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_1059 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_1068 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_1072 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_1080 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_1102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_1106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_1110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1114 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1126 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_119 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_1273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_210 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_232 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_379 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_611 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_630 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_639 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_666 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_674 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_728 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_732 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_736 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_768 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_777 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_846 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_850 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_856 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_860 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_891 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_899 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_903 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_923 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_979 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_987 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_998 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1020 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_1032 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_1042 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_1053 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_1070 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_1079 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_1083 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_1098 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_1102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_1106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_1110 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_1114 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_1251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_426 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_646 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_691 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_695 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_703 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_733 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_766 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_774 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_818 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_826 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_846 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_850 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_859 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_87 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_875 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_879 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_903 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_946 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_953 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_976 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_994 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_1013 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_1017 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_1025 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_103 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_1033 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_1061 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_1071 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_1079 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_1083 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_1096 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_1100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_1108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_1117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_1137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1161 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1229 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_1259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_127 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_1270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_1276 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_381 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_504 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_664 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_682 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_730 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_734 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_742 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_753 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_787 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_824 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_849 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_858 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_862 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_929 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_956 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_96 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_968 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_976 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_998 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_1007 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_1014 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_1028 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_1048 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_1052 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_1071 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_1075 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_1083 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_1087 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_1091 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_1095 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_1110 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_1114 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_1129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_1133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_1137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_1165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_1225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_1231 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_342 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_432 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_500 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_649 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_662 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_760 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_764 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_778 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_805 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_865 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_893 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_902 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_924 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_928 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_932 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_951 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_969 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_1009 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_1032 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_1041 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_1080 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_1084 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_1088 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_1114 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_1127 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_1131 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_119 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_1203 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1218 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_1230 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_1234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_124 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_1270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_1276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_387 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_524 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_604 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_622 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_736 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_74 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_790 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_794 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_798 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_842 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_846 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_850 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_857 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_865 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_875 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_883 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_886 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_890 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_903 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_907 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_925 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_939 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_943 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_955 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_959 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_969 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_991 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_998 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_1000 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_1020 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_1024 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_1028 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_1035 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_1047 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_1061 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_1073 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_1077 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_1085 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_1089 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_1097 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_1110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_1116 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_1124 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_1128 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_1134 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_1143 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1151 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_1226 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_235 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_31 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_455 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_508 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_647 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_655 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_677 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_691 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_753 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_828 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_845 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_857 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_876 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_907 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_911 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_921 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_929 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_949 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_969 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_975 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_982 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1005 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_1027 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_1040 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_1078 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_1083 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_1102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_1106 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_1110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_1116 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_1125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_1156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1160 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1172 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1184 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_1196 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_1221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_1259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_1270 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_1274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_132 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_17 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_242 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_330 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_585 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_607 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_792 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_813 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_830 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_846 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_850 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_857 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_874 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_878 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_923 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_957 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_976 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_1004 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_1025 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_1028 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_1042 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_1075 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_1079 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_1112 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_1125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_1132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_1136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_1140 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_1158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_1162 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_1166 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_1174 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_1185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_1228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_1275 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_148 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_403 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_428 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_490 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_66 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_7 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_70 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_732 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_736 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_759 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_763 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_767 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_791 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_820 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_824 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_836 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_856 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_874 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_892 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_904 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_912 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_928 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_932 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_936 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_940 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_951 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_964 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_971 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_983 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_988 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_1007 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_1026 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_1035 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_1060 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_1070 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_1074 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_1079 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_1084 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_1098 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_1102 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_1117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_112 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_1122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_1126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1154 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1178 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_1190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_1203 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_1211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_1219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_1236 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_1246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_1261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_1265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_1276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_135 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_178 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_182 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_216 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_227 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_339 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_38 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_386 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_394 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_434 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_584 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_608 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_624 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_642 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_666 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_735 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_739 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_809 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_819 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_822 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_826 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_843 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_899 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_903 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_907 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_912 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_916 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_929 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_943 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_979 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_990 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_1014 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_1020 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_1023 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_1027 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_1031 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_1075 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_1079 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_1083 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_1094 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_1103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_1114 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_1118 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_1121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_1136 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_1142 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_1147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_1151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_1155 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1159 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_1175 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_1181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_1206 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_1216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_1224 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_1228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_1237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_1247 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_1251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_182 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_186 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_210 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_276 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_286 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_30 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_431 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_443 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_458 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_500 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_510 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_591 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_610 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_668 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_702 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_738 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_772 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_792 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_796 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_845 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_853 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_873 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_917 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_934 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_938 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_946 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_950 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_972 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_990 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_1022 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_1044 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_1048 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_1067 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_1071 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_1075 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_1079 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_1097 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_1101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_1116 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_1120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_1124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_1147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_1158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_1162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_1166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_1170 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_1178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_1182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_1191 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_1195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1229 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_1273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_329 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_392 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_567 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_626 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_679 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_735 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_845 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_903 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_907 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_922 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_934 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_954 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_964 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_968 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_981 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_10 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_1001 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_1011 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1015 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_1027 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_1032 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_1043 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_1047 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_1068 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_1072 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_1076 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_1084 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_1088 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_1105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_1114 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_1125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_1185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_1198 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_120 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_1270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_1276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_168 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_184 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_188 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_336 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_344 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_516 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_674 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_7 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_728 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_732 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_776 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_780 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_784 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_791 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_943 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_957 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_968 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_977 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_1002 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_1020 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_1024 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_1032 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_1044 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_1052 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_1056 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_1060 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_1069 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_1073 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1096 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_1113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_1189 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_1211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_1217 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_1231 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_263 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_308 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_500 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_555 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_575 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_649 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_668 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_688 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_700 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_708 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_764 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_792 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_807 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_815 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_819 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_822 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_845 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_851 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_888 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_929 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_936 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_945 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_994 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_1018 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_1025 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_1032 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_1042 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_1046 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_1060 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_1064 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_1068 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_1072 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_1086 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_1103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_1107 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_1123 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_1127 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_1146 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1168 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1180 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_1192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_1200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_1229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_1258 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_1270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_1276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_188 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_275 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_37 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_598 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_618 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_630 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_688 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_777 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_788 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_792 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_796 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_823 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_827 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_846 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_850 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_899 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_903 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_907 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_911 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_915 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_923 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_934 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_938 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_961 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_981 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_987 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_995 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_1009 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_1013 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_1023 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_1031 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_1041 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_1062 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_1065 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_1078 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_1091 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_1099 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_1103 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_1119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_1168 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_1210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_1220 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_1229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_1250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_196 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_22 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_294 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_407 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_420 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_596 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_600 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_608 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_630 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_702 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_710 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_763 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_79 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_816 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_822 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_857 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_868 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_87 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_880 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_917 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_925 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_929 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_939 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_943 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_947 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_968 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_987 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_991 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_994 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_1029 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_1041 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_1050 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_1062 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_1069 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1078 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_1117 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_1138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1186 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_1198 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_1205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_1225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_1254 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_127 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_1270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_1276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_146 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_248 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_276 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_630 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_643 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_675 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_735 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_774 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_786 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_80 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_806 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_820 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_824 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_828 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_848 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_878 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_883 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_899 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_908 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_923 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_932 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_946 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_958 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_1014 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_1018 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_1027 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_1041 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_1055 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_1075 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1079 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_1091 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_1106 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_1119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_1166 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_1170 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_1253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_203 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_397 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_546 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_555 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_646 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_662 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_666 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_679 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_691 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_727 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_734 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_738 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_766 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_814 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_818 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_827 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_844 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_848 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_852 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_894 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_934 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_938 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_942 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_959 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_971 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_983 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_991 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_994 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_1000 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_1025 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_1029 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_103 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_1033 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_1044 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_1072 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_1080 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_1084 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_1088 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_1103 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_1114 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_112 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_1123 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_1127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_1134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_1154 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_1158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_1169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_1174 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_1178 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_1186 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_1203 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_1221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_1225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_1249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_1273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_154 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_182 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_486 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_560 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_564 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_660 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_664 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_672 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_775 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_813 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_854 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_865 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_898 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_902 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_906 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_930 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_935 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_943 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_948 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_956 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_968 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_997 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_1002 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_1016 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_1024 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_1028 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_1032 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_1035 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_1072 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_1080 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_1084 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_1088 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_1092 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_1100 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_1114 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_1127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_1133 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_1142 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_1146 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_1160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_1177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_1181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_1189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_1193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_1217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_1221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_1242 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_1246 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_1272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_1276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_135 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_247 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_258 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_354 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_420 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_510 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_520 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_534 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_538 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_585 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_594 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_668 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_692 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_718 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_754 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_770 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_816 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_822 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_826 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_830 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_845 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_853 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_860 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_868 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_879 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_887 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_912 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_926 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_934 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_941 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_951 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_963 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_983 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_987 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_995 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_1003 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_1011 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_1015 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_1041 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_1045 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_1061 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_1084 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_1103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_1115 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_1133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_1136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_1140 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_1144 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_1157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_1173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_1186 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_1194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_1205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_1218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_1237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_1255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_1259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_1261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_1265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_1276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_203 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_224 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_248 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_292 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_494 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_563 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_606 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_619 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_679 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_712 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_716 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_719 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_728 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_740 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_771 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_787 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_790 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_795 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_799 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_807 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_864 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_872 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_905 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_917 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_929 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_941 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_949 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_955 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_963 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_977 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_995 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_1000 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_1004 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_1016 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_1020 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_1029 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_1043 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_1047 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_1060 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_1073 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1081 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_1104 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_1119 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_1128 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_1134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_1137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_1145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_1148 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_1156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_1160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_1168 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_1181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_1224 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_1233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_210 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_264 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_28 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_308 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_328 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_344 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_374 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_487 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_540 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_638 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_664 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_703 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_742 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_771 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_807 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_812 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_845 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_926 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_930 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_938 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_951 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_956 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_964 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_971 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_1029 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_1041 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_1048 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_1056 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_1060 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_1073 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_1077 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_1085 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_1097 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_1101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_1105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_1109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_1113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_1117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_1125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_1133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_1141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_1157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_1161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_1165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_1169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_1173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_1181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_1185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1189 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_126 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_1269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_478 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_526 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_550 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_642 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_669 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_680 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_692 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_738 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_822 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_845 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_862 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_884 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_912 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_945 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_962 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_980 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_984 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_1003 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_1011 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_1051 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_1072 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_1076 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_1080 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_1084 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_1090 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_1100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_1108 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_1116 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_1128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_1133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_1137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_1162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_1170 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_1174 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_1178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_1186 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_1203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_1250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_126 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_1270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_1276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_148 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_23 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_323 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_396 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_507 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_570 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_574 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_594 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_631 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_638 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_674 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_696 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_718 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_730 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_738 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_752 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_767 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_779 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_791 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_795 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_813 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_842 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_858 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_862 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_882 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_886 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_894 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_899 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_908 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_912 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_916 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_932 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_938 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_942 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_977 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_985 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_988 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_999 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_1016 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_1020 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_1024 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_1028 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_1036 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_1040 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_1044 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_1048 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1080 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_1092 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1104 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_1116 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_1168 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_1172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_1193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_1205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_1242 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_173 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_217 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_240 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_322 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_359 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_444 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_458 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_648 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_670 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_704 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_733 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_746 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_790 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_807 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_815 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_822 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_857 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_861 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_877 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_883 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_886 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_906 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_914 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_923 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_935 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_943 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_965 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_973 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_977 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_988 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_996 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_1000 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_1004 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_1015 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_1022 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_1027 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_1041 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_1055 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_1078 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_1082 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_1086 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_1101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1122 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_1216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_1258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_1270 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_1274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_208 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_212 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_226 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_263 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_292 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_346 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_59 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_630 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_737 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_772 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_776 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_784 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_803 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_810 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_827 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_844 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_856 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_867 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_877 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_884 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_893 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_954 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_969 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_973 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_986 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_990 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_996 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_1029 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_1041 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_1045 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_1071 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1075 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1087 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_1119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_1121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_1135 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_1143 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_1148 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_1152 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_1218 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_1241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_1247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_1271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_140 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_323 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_356 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_376 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_412 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_45 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_462 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_626 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_630 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_650 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_670 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_794 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_812 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_823 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_846 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_850 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_854 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_862 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_870 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_876 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_879 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_891 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_894 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_904 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_912 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_933 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_945 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_96 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_973 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_982 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_999 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_1002 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_1010 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_1014 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_1024 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_1041 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_1050 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_1058 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_1071 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_1075 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_1082 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_1091 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_1106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_1114 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_1124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_1133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_115 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_1153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_1170 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_1178 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_1205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_1223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_1229 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_1254 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_1270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_1276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_182 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_230 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_336 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_347 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_351 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_487 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_730 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_743 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_750 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_777 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_782 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_786 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_800 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_804 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_824 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_839 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_857 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_861 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_864 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_884 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_888 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_899 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_906 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_918 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_936 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_944 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_954 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_959 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_978 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_989 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_998 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_1029 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_1037 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_1041 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_1075 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_1079 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_1088 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_1094 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_1102 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_1114 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_1128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_1134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_1138 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_1146 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_1155 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_1189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_1193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1215 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_1231 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_1249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_1253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_142 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_175 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_343 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_410 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_422 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_430 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_510 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_556 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_593 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_621 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_646 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_692 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_714 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_742 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_792 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_848 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_858 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_86 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_866 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_870 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_895 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_924 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_930 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_940 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_957 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_969 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_1001 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_1019 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_1023 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_1027 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_1041 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_1058 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_1076 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1080 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_1125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_1129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_1133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_1136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_1154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_1161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1170 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_1182 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_1186 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_1198 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_1209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_1257 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_126 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_1270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_1276 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_403 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_412 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_458 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_491 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_629 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_643 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_679 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_696 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_715 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_755 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_760 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_79 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_794 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_809 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_826 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_848 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_857 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_873 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_890 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_906 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_951 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_955 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_969 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_985 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_1004 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_1018 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_1027 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_1031 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_1039 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_1043 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_1062 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_1071 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_1075 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1079 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_1091 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_1100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_1106 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_1114 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_1126 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_1136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_1168 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_1172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_1195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_1237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_17 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_247 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_254 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_260 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_328 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_487 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_492 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_584 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_640 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_697 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_762 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_766 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_799 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_814 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_818 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_826 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_866 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_87 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_870 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_878 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_886 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_892 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_907 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_921 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_934 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_939 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_943 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_947 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_972 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_976 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_979 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_989 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_997 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_1030 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_1046 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_1070 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_1074 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_1078 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_1100 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_1113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_1123 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_1127 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_1132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_1141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_1145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_1202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_1214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_1231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_1242 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_1259 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_1270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_1276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_176 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_180 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_226 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_236 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_275 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_341 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_354 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_618 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_640 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_682 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_698 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_754 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_802 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_833 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_852 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_858 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_881 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_885 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_902 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_922 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_933 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_942 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_946 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_954 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_964 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_968 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_985 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_997 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_1025 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_1033 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_1065 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_1075 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_1079 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_1090 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_1098 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_1109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_1115 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_1131 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_1137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_1167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_1181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_1185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_1189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_1193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_1201 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_1233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_1248 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_1274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_145 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_254 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_340 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_492 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_513 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_538 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_650 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_706 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_760 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_773 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_802 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_823 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_833 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_845 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_861 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_873 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_895 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_926 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_958 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_962 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_971 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_978 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_985 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_996 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_1046 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_1070 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_1074 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_1078 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_1082 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_1086 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_1108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_1125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_1172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_1176 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1180 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_1273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_398 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_674 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_74 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_768 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_784 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_788 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_792 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_800 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_820 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_824 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_828 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_846 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_850 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_854 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_873 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_880 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_884 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_929 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_976 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_1010 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_1014 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_1018 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_1077 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_1081 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_1091 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_1099 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_1105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_1118 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_1122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_1164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_1168 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_1173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_1181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_1198 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_1205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_1218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_1244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_1248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_1251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_1270 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_1274 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_204 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_450 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_492 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_507 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_526 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_541 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_562 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_566 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_628 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_675 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_768 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_793 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_822 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_842 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_847 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_855 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_867 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_873 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_891 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_898 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_921 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_930 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_947 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_956 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_960 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_964 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_968 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_976 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_1001 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_1009 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_1013 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_1023 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_1032 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_1040 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_1056 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_1060 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_1069 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_1073 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_1081 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_1098 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_11 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_1107 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_1112 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_1116 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_1133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_1164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_1170 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_1177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_1181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_1208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_1230 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_1242 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_152 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_238 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_276 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_30 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_323 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_406 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_431 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_435 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_460 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_476 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_500 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_639 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_679 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_691 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_782 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_805 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_828 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_871 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_880 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_908 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_917 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_932 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_940 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_966 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_10 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_1009 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_1013 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_1044 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_1048 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_1052 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_1056 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_1060 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_1064 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1068 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_1080 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_1105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_1113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_1117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_1124 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_1128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_1146 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_1157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_1167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_1171 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_1179 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_1183 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_1205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_1209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_1259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_1270 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_1274 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_132 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_168 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_201 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_210 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_547 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_562 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_619 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_630 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_655 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_667 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_694 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_706 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_736 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_764 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_791 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_795 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_821 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_855 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_859 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_867 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_895 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_898 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_902 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_940 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_956 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_960 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_971 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_996 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_1005 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_1018 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_1041 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_1049 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_1061 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_1069 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_1096 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_1100 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_1104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_1109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_1113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_1117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_1125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_1189 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_1245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_142 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_175 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_47 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_496 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_564 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_592 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_715 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_736 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_756 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_760 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_788 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_812 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_816 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_845 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_855 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_872 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_880 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_926 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_958 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_962 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_967 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_1010 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_1051 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_1059 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_1072 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_1080 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_1090 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_1106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_1165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_1205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_1228 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_1232 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_1236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_1248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_1252 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_1255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_1259 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_1270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_1276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_323 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_395 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_443 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_506 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_569 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_606 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_627 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_631 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_652 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_664 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_681 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_718 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_725 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_734 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_747 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_761 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_776 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_788 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_804 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_857 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_917 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_938 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_946 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_954 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_958 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_962 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_966 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_1006 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_1031 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_1043 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1047 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1073 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_1089 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_1097 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_1100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_1107 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_1126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_1130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_1134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_1142 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_1152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_1161 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_1165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_1173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_1177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_1185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_1204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_1221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_1258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_126 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_1268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_1276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_151 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_17 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_196 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_295 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_319 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_350 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_583 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_588 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_599 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_622 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_668 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_678 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_694 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_702 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_770 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_797 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_807 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_815 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_836 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_848 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_855 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_866 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_878 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_894 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_897 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_928 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_932 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_968 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_972 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_986 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_1008 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_1030 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_1034 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_1043 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_1047 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_1055 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_1077 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_1086 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_1100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_1117 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_1126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_1139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_1153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_117 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_1174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_1180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_1213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_1273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_292 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_336 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_384 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_455 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_459 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_484 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_618 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_672 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_676 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_699 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_794 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_813 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_830 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_858 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_915 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_923 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_933 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_957 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_969 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_976 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_1025 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_1029 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_1033 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_1045 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_1053 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_1061 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_1072 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_1080 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_1086 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_1090 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_1094 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_1102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_1133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_1142 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_1146 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_1150 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_1189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_1199 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_1207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_1228 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_123 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_1274 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_323 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_340 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_402 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_438 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_476 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_519 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_572 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_631 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_687 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_736 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_762 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_774 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_807 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_833 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_875 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_880 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_884 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_892 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_902 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_920 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_924 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_932 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_939 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_948 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_953 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_958 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_963 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_967 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_999 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_1014 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_1026 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_1030 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_1048 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_1061 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_1068 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_1078 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_1082 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_1086 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_1090 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_1100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_1146 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_1154 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1158 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_1170 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_1178 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_1196 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_1214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_1270 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_1274 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_313 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_404 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_438 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_44 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_488 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_560 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_619 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_627 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_674 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_678 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_705 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_744 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_845 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_859 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_890 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_900 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_908 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_917 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_92 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_929 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_937 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_941 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_947 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_954 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_958 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_962 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_978 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_997 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1025 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_1058 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_1072 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_1076 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_1085 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_1095 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_1099 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_1119 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_1150 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_1189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_1222 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_1226 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_1237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_243 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_347 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_444 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_49 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_536 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_570 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_700 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_704 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_736 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_740 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_744 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_750 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_756 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_764 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_771 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_779 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_791 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_824 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_828 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_839 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_844 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_850 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_859 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_872 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_879 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_883 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_897 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_911 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_924 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_945 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_953 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_990 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_994 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_998 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_1000 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_1023 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_1027 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_1074 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_1078 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_1097 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_1101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_1132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_1136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_1156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_1165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_1169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_1269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_379 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_406 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_472 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_478 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_555 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_621 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_681 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_801 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_822 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_826 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_846 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_850 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_854 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_868 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_872 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_876 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_880 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_884 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_911 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_927 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_935 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_939 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_943 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_978 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_982 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_992 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_996 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_1005 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_1011 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_1018 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_102 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_1034 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_1047 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_1063 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_1080 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_1106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_1123 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1128 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_1140 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_1173 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_1181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_1230 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_1238 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_1259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_1270 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_1274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_201 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_42 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_528 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_593 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_602 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_622 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_631 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_672 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_707 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_724 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_728 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_767 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_771 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_787 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_796 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_823 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_827 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_847 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_856 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_872 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_876 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_885 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_892 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_898 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_906 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_914 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_930 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_934 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_941 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_956 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_960 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_968 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_1007 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_1019 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_1023 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1030 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_1042 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_1050 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_1069 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_1088 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_1098 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_1102 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_1106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_1112 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_1133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1156 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_1168 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1189 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_1207 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_1239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_1276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_164 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_247 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_308 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_356 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_453 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_478 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_556 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_566 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_570 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_634 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_640 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_700 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_704 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_732 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_736 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_783 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_791 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_796 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_814 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_818 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_826 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_844 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_86 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_867 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_875 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_894 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_907 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_911 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_920 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_941 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_963 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_982 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_986 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_990 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_10 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_1035 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_1050 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_1062 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_1071 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_1079 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_1083 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_1087 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_1097 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_1105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_1111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_1120 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_1136 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_1145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_1152 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_1193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_1201 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_1211 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_1235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_1270 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_1274 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_226 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_350 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_510 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_642 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_730 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_734 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_782 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_786 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_790 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_798 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_818 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_830 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_842 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_850 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_854 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_879 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_883 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_887 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_898 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_906 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_922 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_968 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_976 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_1018 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_1031 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_1052 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_1077 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_1085 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_1092 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_1107 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_1117 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_1126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_1141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_1155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_1163 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1201 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_1213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_1217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_1229 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_1271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_1275 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_469 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_481 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_588 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_646 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_687 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_756 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_768 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_772 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_776 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_807 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_814 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_826 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_848 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_852 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_856 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_871 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_875 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_883 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_887 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_929 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_938 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_942 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_951 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_965 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_969 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_975 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_981 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_995 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_1001 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_1014 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_1026 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_1030 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_1074 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_1084 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_1091 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_1105 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_1109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_1117 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_1145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_1153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_1157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_1161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_1165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_1169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1217 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_1229 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_1270 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_1274 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_224 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_338 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_354 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_444 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_46 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_468 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_572 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_586 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_625 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_662 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_858 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_876 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_880 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_921 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_932 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_936 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_945 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_958 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_962 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_979 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_988 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_1000 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1016 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1028 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_1040 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_1058 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_1094 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_1098 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_1102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_1106 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_1110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_1119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_1142 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_1150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_1154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_1158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_1162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_1166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_1170 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_1253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_211 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_243 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_308 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_415 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_459 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_48 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_52 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_575 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_600 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_625 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_653 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_690 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_705 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_743 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_763 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_767 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_814 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_818 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_830 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_857 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_861 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_914 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_918 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_924 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_938 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_942 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_946 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_980 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_988 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_1025 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_1033 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_1050 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_1064 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_1074 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_1078 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_1097 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_1101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_1105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_1109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_1113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_1142 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_1153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_1157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_1161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_1165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_1169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_1173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_1181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_1185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_1201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_1213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_1270 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_1274 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_369 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_400 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_404 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_582 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_674 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_686 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_731 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_778 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_791 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_795 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_840 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_846 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_873 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_877 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_890 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_898 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_908 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_914 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_945 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_949 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_957 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_974 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_1033 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_1040 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_1056 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_1060 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_1088 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_1092 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_1096 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_1100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_1104 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_1108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_1113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_1117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_1125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_1133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_1137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_1158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_1162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_1166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_1170 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_1193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_1197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_1242 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_1246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_1275 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_198 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_252 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_256 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_275 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_424 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_463 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_470 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_567 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_585 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_646 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_660 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_703 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_720 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_780 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_801 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_808 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_846 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_850 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_854 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_858 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_873 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_904 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_908 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_935 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_939 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_943 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_953 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_959 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_969 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_984 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_1003 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_1018 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_1025 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_1058 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_1066 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_1070 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_1087 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_1096 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_1103 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_1107 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_1126 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_1130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_1165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_1169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_1173 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_1193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_1203 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_1257 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_1270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_1276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_257 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_410 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_428 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_507 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_511 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_562 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_612 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_670 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_674 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_752 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_768 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_780 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_784 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_802 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_850 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_929 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_950 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_959 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_978 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_99 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_997 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_10 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_1012 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_1020 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_1024 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_1044 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_1048 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_1053 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_1061 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_1085 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_1089 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_1114 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_1140 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_1166 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_1210 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_1214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_1220 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_1223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_490 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_567 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_574 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_662 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_700 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_704 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_710 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_739 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_763 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_792 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_796 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_808 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_812 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_816 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_819 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_845 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_86 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_872 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_882 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_893 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_908 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_917 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_929 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_978 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_984 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_995 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_1003 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_1019 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_1023 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_1027 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_1041 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_1076 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_1080 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_1084 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_1088 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_1097 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_1101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_1109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_1132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_1136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_1140 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_1144 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1171 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1183 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_1195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1229 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_1273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_176 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_275 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_462 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_564 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_675 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_794 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_810 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_821 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_855 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_863 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_875 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_890 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_902 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_935 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_939 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_943 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_952 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_976 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_987 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_995 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_1002 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_1016 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_1025 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_1031 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_1052 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_1056 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_1060 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_1074 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_1078 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_1082 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_1117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_1140 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_1144 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_1157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_1169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_1173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_1185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_1195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_1210 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_1221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_1255 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_1270 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_1274 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_188 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_201 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_204 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_608 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_618 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_664 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_668 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_719 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_728 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_794 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_817 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_823 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_840 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_844 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_851 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_875 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_920 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_952 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_956 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_979 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_981 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_1007 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_1013 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_1020 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_1030 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_1041 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_1058 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_1073 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_1077 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_1081 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_1085 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_1090 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_1105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_1116 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_1127 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_1133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_1142 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_1150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_1154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_1164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_1180 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_1184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_1192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_1202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_1206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_1231 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_1238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_1251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_1276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_202 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_372 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_376 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_633 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_654 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_676 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_683 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_708 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_792 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_796 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_822 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_851 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_855 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_859 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_878 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_887 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_895 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_905 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_911 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_920 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_924 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_956 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_977 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_1002 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_1006 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_1010 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_1014 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_1017 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_1032 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_1043 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_1047 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_1051 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_1075 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_1085 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_1093 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_1100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_1109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_1126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_1130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_1197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_1205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_1209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_1213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_1217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_1232 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_1236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_1270 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_1274 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_215 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_386 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_425 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_454 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_480 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_504 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_584 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_616 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_620 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_628 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_638 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_658 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_676 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_683 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_70 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_717 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_734 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_764 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_780 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_784 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_794 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_834 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_842 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_848 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_852 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_858 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_942 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_954 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_958 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_976 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_995 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_1002 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_1013 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_1033 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_1053 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_1094 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_1098 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_1102 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_1119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_1124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_1128 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_1132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_1154 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_1204 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_1230 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_1252 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_276 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_30 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_435 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_492 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_588 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_628 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_655 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_691 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_703 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_758 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_762 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_768 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_795 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_808 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_812 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_820 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_824 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_886 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_907 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_915 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_932 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_944 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_974 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_980 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_10 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_1001 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_1013 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_1019 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_1032 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_1042 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_1046 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_1056 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_1093 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_1128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_1160 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_1164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_1202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_1253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_1257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_1270 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_1274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_202 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_291 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_40 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_500 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_562 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_579 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_625 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_629 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_669 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_738 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_764 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_768 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_787 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_796 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_818 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_822 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_834 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_838 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_847 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_853 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_911 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_923 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_945 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_955 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_959 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_994 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_1029 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_1038 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_1042 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_1056 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_1065 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_1118 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_1154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_1199 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_1203 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_1207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_1253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_182 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_202 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_354 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_366 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_591 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_599 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_630 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_652 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_664 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_682 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_692 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_704 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_715 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_770 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_798 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_828 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_849 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_883 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_938 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_965 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_969 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_993 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_997 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_1013 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_1017 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_1037 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_1044 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_1073 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_1091 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_1104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_1205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_1209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_1254 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_1258 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_1270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_1276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_171 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_44 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_596 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_618 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_683 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_710 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_765 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_834 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_845 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_853 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_866 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_877 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_902 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_956 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_969 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_984 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_996 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_1009 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_1029 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_1048 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_1058 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_1079 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_1083 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_1087 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_1099 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_1119 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_1174 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_1185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1191 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_1220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_1237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_1270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_1276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_207 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_30 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_48 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_52 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_602 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_629 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_637 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_647 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_656 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_694 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_750 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_754 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_759 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_792 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_796 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_807 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_844 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_895 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_935 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_939 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_946 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_975 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_979 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_983 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_1012 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_1041 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_1064 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_1068 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_1072 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_1079 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_1083 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_1090 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_1142 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1184 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_1196 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_1250 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_1270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_1276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_324 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_392 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_555 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_564 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_596 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_608 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_628 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_654 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_662 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_672 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_748 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_764 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_787 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_791 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_795 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_811 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_824 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_831 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_840 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_864 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_893 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_929 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_933 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_962 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_966 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_986 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_995 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_1022 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_1030 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_1038 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_1042 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_1046 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_1055 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_108 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_1103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_1111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_1114 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_1145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_1149 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_1153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_1253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_142 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_162 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_295 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_367 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_379 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_588 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_714 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_726 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_736 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_740 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_766 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_795 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_805 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_812 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_845 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_857 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_889 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_923 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_936 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_968 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_1000 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_1014 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_1018 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_1024 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_1028 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_1034 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_1073 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_1077 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_1085 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_1097 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_1105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_1108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_1112 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_1116 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_1128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_1132 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_1136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_1159 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1213 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_1269 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_423 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_476 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_644 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_739 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_762 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_776 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_791 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_795 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_801 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_820 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_836 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_86 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_873 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_894 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_90 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_904 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_926 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_932 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_936 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_958 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_962 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_985 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_989 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_1027 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_1041 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_1045 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_1130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_1134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_1138 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_1142 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_1257 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_1270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_1276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_285 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_394 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_472 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_661 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_678 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_705 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_736 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_767 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_786 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_790 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_802 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_808 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_821 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_828 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_857 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_879 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_888 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_943 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_984 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_988 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_1004 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_1017 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_1023 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_1083 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_1087 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_1095 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_1103 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_1107 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1150 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1189 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_1218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_1222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_1226 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_124 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_1242 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_1271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_136 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_163 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_457 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_551 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_566 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_626 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_695 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_758 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_762 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_766 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_805 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_838 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_849 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_87 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_905 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_922 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_936 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_957 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_978 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_987 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_104 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_1066 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_1070 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_1076 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_1107 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_1111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_1115 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1131 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_1143 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1186 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_119 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_1198 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_1205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_1218 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_1243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_1270 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_1274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_23 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_328 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_516 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_560 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_572 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_655 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_674 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_731 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_735 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_754 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_765 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_768 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_776 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_808 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_845 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_857 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_874 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_929 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_933 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_947 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_951 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_955 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_963 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_966 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_971 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_1001 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_1016 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_1020 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_1047 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_1116 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_1121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_1129 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_1134 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_1140 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_1145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_1149 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_1153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_1158 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_1245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_1276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_190 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_239 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_248 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_252 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_30 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_310 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_328 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_40 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_576 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_588 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_644 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_648 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_666 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_686 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_698 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_706 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_722 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_736 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_759 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_778 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_808 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_816 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_861 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_870 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_900 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_912 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_916 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_920 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_930 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_945 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_965 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_971 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_985 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_997 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_1015 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_1032 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_1040 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_1044 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_1101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_1105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_1109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_1113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_1117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_1132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_1157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_1166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_1170 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1174 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_1186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_1194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_1221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_1238 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_1258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_1270 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_1274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_145 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_163 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_244 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_444 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_448 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_544 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_620 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_642 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_663 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_675 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_687 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_695 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_720 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_738 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_762 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_767 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_771 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_781 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_789 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_842 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_850 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_874 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_878 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_896 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_900 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_912 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_936 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_952 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_956 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_1068 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_1097 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_1119 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_1125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_1128 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_1132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_1153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_1163 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_1192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_1212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_1242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_247 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_286 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_316 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_328 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_364 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_534 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_575 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_586 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_604 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_650 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_670 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_677 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_706 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_759 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_80 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_819 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_845 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_870 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_874 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_882 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_888 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_903 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_912 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_930 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_934 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_957 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_980 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_997 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_1014 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_1046 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_1072 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_1124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_1128 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_1132 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_1137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_1144 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_1158 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_1191 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_1205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_1235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_1246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_1256 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_1270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_1276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_168 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_264 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_327 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_564 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_578 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_614 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_655 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_663 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_682 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_686 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_716 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_761 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_782 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_843 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_852 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_856 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_860 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_864 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_886 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_890 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_896 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_899 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_969 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_1020 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_1046 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_1073 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1077 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_1133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_1137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_1169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_1173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_1186 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_1202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_1226 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_1230 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_160 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_20 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_32 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_403 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_491 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_564 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_574 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_590 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_594 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_622 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_659 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_666 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_688 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_756 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_780 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_79 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_827 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_845 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_855 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_870 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_874 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_880 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_884 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_911 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_915 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_927 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_942 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_946 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_957 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_980 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_1014 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_1041 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_1073 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_1089 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_1125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_1133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_1146 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_1160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_1185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_1214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_1227 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_1270 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_1274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_151 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_192 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_227 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_25 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_352 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_392 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_462 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_482 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_56 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_565 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_606 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_626 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_688 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_706 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_731 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_766 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_774 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_778 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_790 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_800 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_808 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_816 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_824 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_839 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_842 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_877 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_882 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_898 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_936 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_940 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_952 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_959 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_1007 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_1025 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_1029 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_1033 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_1041 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_1073 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_1077 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_1103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_1125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_1129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_1172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_1185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_1189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_119 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_1193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_1231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_1243 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_319 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_323 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_622 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_626 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_66 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_688 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_710 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_715 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_736 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_759 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_80 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_817 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_854 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_872 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_876 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_880 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_913 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_930 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_939 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_957 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_992 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_1002 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_1024 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_1056 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_1060 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_1064 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_1068 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_1072 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1076 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_1273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_220 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_226 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_403 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_519 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_527 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_579 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_690 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_721 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_746 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_810 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_820 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_840 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_844 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_848 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_852 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_856 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_876 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_880 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_891 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_929 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_952 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_956 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_965 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_986 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_990 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_994 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_998 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_1004 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_1023 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_1027 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_1048 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_1052 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_1086 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_1093 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_1106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_1114 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_1118 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_1123 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_1142 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_1196 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_1200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_1236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_1256 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_1270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_1276 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_238 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_257 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_319 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_379 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_392 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_410 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_427 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_470 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_540 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_574 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_580 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_599 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_619 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_663 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_667 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_708 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_712 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_773 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_791 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_800 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_804 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_860 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_878 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_887 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_891 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_911 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_929 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_946 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_954 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_958 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_962 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_966 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_981 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_985 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_1006 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_1031 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_1036 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_1040 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_1061 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_1073 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_1116 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_1125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_1129 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_1141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_1152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_1202 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_1210 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_1229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_1251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_1275 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_231 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_32 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_386 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_420 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_52 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_567 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_584 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_592 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_606 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_610 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_62 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_738 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_760 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_764 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_839 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_84 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_857 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_861 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_895 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_907 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_916 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_920 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_930 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_940 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_948 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_968 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_976 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_980 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_984 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_988 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_992 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_1008 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_1032 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_1052 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_1069 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_1090 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_1109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_1127 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_1131 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_1139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_1145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_1157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_1166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_1180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_1191 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_1195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_1209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_1213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_1216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_1220 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_1244 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_1258 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_1270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_1276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_186 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_226 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_230 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_275 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_291 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_303 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_562 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_576 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_611 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_621 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_675 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_695 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_732 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_736 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_754 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_762 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_771 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_786 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_791 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_795 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_799 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_844 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_848 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_851 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_866 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_9 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_943 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_947 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_954 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_963 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_978 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_1005 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_1023 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_1036 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_1041 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_1053 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_1092 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_1124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_1128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_1132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_1151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_1155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_1163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_1167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_1173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_1186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_1190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_1194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_1198 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_120 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_1229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_1242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_154 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_191 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_272 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_311 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_351 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_378 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_404 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_434 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_456 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_472 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_496 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_532 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_588 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_600 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_613 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_622 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_653 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_700 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_735 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_766 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_795 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_803 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_816 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_830 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_845 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_865 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_875 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_885 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_889 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_907 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_920 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_935 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_939 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_946 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_992 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_1006 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_1012 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_1023 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_1075 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_1083 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_1097 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_1101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_1106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_1111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_1115 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_1119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_1123 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_1144 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_1158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_1193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_1197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_1201 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_1243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_1247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_1251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_1270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_1276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_207 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_259 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_504 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_662 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_679 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_683 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_730 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_734 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_738 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_746 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_762 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_777 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_789 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_809 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_833 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_840 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_881 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_890 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_898 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_920 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_936 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_958 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_962 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_1005 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_1042 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_1060 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_1085 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_1092 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_1103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_1108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_1121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_1125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_1132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_1151 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1196 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_1224 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_1241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_1276 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_142 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_22 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_341 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_364 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_412 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_457 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_481 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_554 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_591 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_647 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_668 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_678 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_756 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_760 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_764 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_782 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_815 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_839 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_863 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_875 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_897 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_918 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_934 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_944 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_990 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_999 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_1002 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_1025 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_1088 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_1117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_1128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_1135 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_1144 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_1157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_1161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_1190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_1194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_1198 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_1202 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_1228 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_1242 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_1259 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_1270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_1276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_235 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_273 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_336 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_370 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_507 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_560 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_585 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_634 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_638 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_672 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_686 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_697 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_764 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_768 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_806 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_832 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_844 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_905 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_909 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_917 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_932 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_936 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_967 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_994 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_1018 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_1022 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_1030 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_1038 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_1053 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_1085 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_1089 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_1101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_1162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_1166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_1170 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_1184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_1188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_1192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_1196 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_1216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_1226 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_1253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_132 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_229 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_375 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_399 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_420 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_556 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_566 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_684 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_792 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_804 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_816 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_820 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_828 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_909 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_96 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_1023 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_1027 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_1041 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_1077 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_1097 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_1139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_1154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_1158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_1162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_1166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_1194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_1205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_1215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_1242 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_1259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_1270 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_1274 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_220 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_295 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_338 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_416 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_431 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_512 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_516 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_638 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_735 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_773 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_994 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_1007 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_1040 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_1044 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_1048 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_1052 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_1056 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_1060 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_1096 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_1100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_1104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_1133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_1137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_1150 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_1154 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_1165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_1194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_1198 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_1202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_1206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_207 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_216 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_22 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_235 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_343 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_471 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_487 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_566 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_648 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_761 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_930 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_953 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_1005 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_1025 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_1029 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_1033 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_1044 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_1052 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_1056 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_1060 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1069 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1081 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_1117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_1129 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_1142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_117 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_1170 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_1269 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_143 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_155 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_214 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_319 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_364 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_368 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_476 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_500 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_647 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_658 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_662 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_679 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_727 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_756 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_760 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_764 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_768 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_793 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_806 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_845 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_857 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_863 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_870 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_874 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_878 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_883 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_887 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_917 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_929 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_946 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_957 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_965 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_969 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_978 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_982 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_988 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_992 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_996 ();
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_148 ();
 sky130_fd_sc_hd__decap_3 PHY_149 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_150 ();
 sky130_fd_sc_hd__decap_3 PHY_151 ();
 sky130_fd_sc_hd__decap_3 PHY_152 ();
 sky130_fd_sc_hd__decap_3 PHY_153 ();
 sky130_fd_sc_hd__decap_3 PHY_154 ();
 sky130_fd_sc_hd__decap_3 PHY_155 ();
 sky130_fd_sc_hd__decap_3 PHY_156 ();
 sky130_fd_sc_hd__decap_3 PHY_157 ();
 sky130_fd_sc_hd__decap_3 PHY_158 ();
 sky130_fd_sc_hd__decap_3 PHY_159 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_160 ();
 sky130_fd_sc_hd__decap_3 PHY_161 ();
 sky130_fd_sc_hd__decap_3 PHY_162 ();
 sky130_fd_sc_hd__decap_3 PHY_163 ();
 sky130_fd_sc_hd__decap_3 PHY_164 ();
 sky130_fd_sc_hd__decap_3 PHY_165 ();
 sky130_fd_sc_hd__decap_3 PHY_166 ();
 sky130_fd_sc_hd__decap_3 PHY_167 ();
 sky130_fd_sc_hd__decap_3 PHY_168 ();
 sky130_fd_sc_hd__decap_3 PHY_169 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_170 ();
 sky130_fd_sc_hd__decap_3 PHY_171 ();
 sky130_fd_sc_hd__decap_3 PHY_172 ();
 sky130_fd_sc_hd__decap_3 PHY_173 ();
 sky130_fd_sc_hd__decap_3 PHY_174 ();
 sky130_fd_sc_hd__decap_3 PHY_175 ();
 sky130_fd_sc_hd__decap_3 PHY_176 ();
 sky130_fd_sc_hd__decap_3 PHY_177 ();
 sky130_fd_sc_hd__decap_3 PHY_178 ();
 sky130_fd_sc_hd__decap_3 PHY_179 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_180 ();
 sky130_fd_sc_hd__decap_3 PHY_181 ();
 sky130_fd_sc_hd__decap_3 PHY_182 ();
 sky130_fd_sc_hd__decap_3 PHY_183 ();
 sky130_fd_sc_hd__decap_3 PHY_184 ();
 sky130_fd_sc_hd__decap_3 PHY_185 ();
 sky130_fd_sc_hd__decap_3 PHY_186 ();
 sky130_fd_sc_hd__decap_3 PHY_187 ();
 sky130_fd_sc_hd__decap_3 PHY_188 ();
 sky130_fd_sc_hd__decap_3 PHY_189 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_190 ();
 sky130_fd_sc_hd__decap_3 PHY_191 ();
 sky130_fd_sc_hd__decap_3 PHY_192 ();
 sky130_fd_sc_hd__decap_3 PHY_193 ();
 sky130_fd_sc_hd__decap_3 PHY_194 ();
 sky130_fd_sc_hd__decap_3 PHY_195 ();
 sky130_fd_sc_hd__decap_3 PHY_196 ();
 sky130_fd_sc_hd__decap_3 PHY_197 ();
 sky130_fd_sc_hd__decap_3 PHY_198 ();
 sky130_fd_sc_hd__decap_3 PHY_199 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_200 ();
 sky130_fd_sc_hd__decap_3 PHY_201 ();
 sky130_fd_sc_hd__decap_3 PHY_202 ();
 sky130_fd_sc_hd__decap_3 PHY_203 ();
 sky130_fd_sc_hd__decap_3 PHY_204 ();
 sky130_fd_sc_hd__decap_3 PHY_205 ();
 sky130_fd_sc_hd__decap_3 PHY_206 ();
 sky130_fd_sc_hd__decap_3 PHY_207 ();
 sky130_fd_sc_hd__decap_3 PHY_208 ();
 sky130_fd_sc_hd__decap_3 PHY_209 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_210 ();
 sky130_fd_sc_hd__decap_3 PHY_211 ();
 sky130_fd_sc_hd__decap_3 PHY_212 ();
 sky130_fd_sc_hd__decap_3 PHY_213 ();
 sky130_fd_sc_hd__decap_3 PHY_214 ();
 sky130_fd_sc_hd__decap_3 PHY_215 ();
 sky130_fd_sc_hd__decap_3 PHY_216 ();
 sky130_fd_sc_hd__decap_3 PHY_217 ();
 sky130_fd_sc_hd__decap_3 PHY_218 ();
 sky130_fd_sc_hd__decap_3 PHY_219 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_220 ();
 sky130_fd_sc_hd__decap_3 PHY_221 ();
 sky130_fd_sc_hd__decap_3 PHY_222 ();
 sky130_fd_sc_hd__decap_3 PHY_223 ();
 sky130_fd_sc_hd__decap_3 PHY_224 ();
 sky130_fd_sc_hd__decap_3 PHY_225 ();
 sky130_fd_sc_hd__decap_3 PHY_226 ();
 sky130_fd_sc_hd__decap_3 PHY_227 ();
 sky130_fd_sc_hd__decap_3 PHY_228 ();
 sky130_fd_sc_hd__decap_3 PHY_229 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_230 ();
 sky130_fd_sc_hd__decap_3 PHY_231 ();
 sky130_fd_sc_hd__decap_3 PHY_232 ();
 sky130_fd_sc_hd__decap_3 PHY_233 ();
 sky130_fd_sc_hd__decap_3 PHY_234 ();
 sky130_fd_sc_hd__decap_3 PHY_235 ();
 sky130_fd_sc_hd__decap_3 PHY_236 ();
 sky130_fd_sc_hd__decap_3 PHY_237 ();
 sky130_fd_sc_hd__decap_3 PHY_238 ();
 sky130_fd_sc_hd__decap_3 PHY_239 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_240 ();
 sky130_fd_sc_hd__decap_3 PHY_241 ();
 sky130_fd_sc_hd__decap_3 PHY_242 ();
 sky130_fd_sc_hd__decap_3 PHY_243 ();
 sky130_fd_sc_hd__decap_3 PHY_244 ();
 sky130_fd_sc_hd__decap_3 PHY_245 ();
 sky130_fd_sc_hd__decap_3 PHY_246 ();
 sky130_fd_sc_hd__decap_3 PHY_247 ();
 sky130_fd_sc_hd__decap_3 PHY_248 ();
 sky130_fd_sc_hd__decap_3 PHY_249 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_250 ();
 sky130_fd_sc_hd__decap_3 PHY_251 ();
 sky130_fd_sc_hd__decap_3 PHY_252 ();
 sky130_fd_sc_hd__decap_3 PHY_253 ();
 sky130_fd_sc_hd__decap_3 PHY_254 ();
 sky130_fd_sc_hd__decap_3 PHY_255 ();
 sky130_fd_sc_hd__decap_3 PHY_256 ();
 sky130_fd_sc_hd__decap_3 PHY_257 ();
 sky130_fd_sc_hd__decap_3 PHY_258 ();
 sky130_fd_sc_hd__decap_3 PHY_259 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_260 ();
 sky130_fd_sc_hd__decap_3 PHY_261 ();
 sky130_fd_sc_hd__decap_3 PHY_262 ();
 sky130_fd_sc_hd__decap_3 PHY_263 ();
 sky130_fd_sc_hd__decap_3 PHY_264 ();
 sky130_fd_sc_hd__decap_3 PHY_265 ();
 sky130_fd_sc_hd__decap_3 PHY_266 ();
 sky130_fd_sc_hd__decap_3 PHY_267 ();
 sky130_fd_sc_hd__decap_3 PHY_268 ();
 sky130_fd_sc_hd__decap_3 PHY_269 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_270 ();
 sky130_fd_sc_hd__decap_3 PHY_271 ();
 sky130_fd_sc_hd__decap_3 PHY_272 ();
 sky130_fd_sc_hd__decap_3 PHY_273 ();
 sky130_fd_sc_hd__decap_3 PHY_274 ();
 sky130_fd_sc_hd__decap_3 PHY_275 ();
 sky130_fd_sc_hd__decap_3 PHY_276 ();
 sky130_fd_sc_hd__decap_3 PHY_277 ();
 sky130_fd_sc_hd__decap_3 PHY_278 ();
 sky130_fd_sc_hd__decap_3 PHY_279 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_280 ();
 sky130_fd_sc_hd__decap_3 PHY_281 ();
 sky130_fd_sc_hd__decap_3 PHY_282 ();
 sky130_fd_sc_hd__decap_3 PHY_283 ();
 sky130_fd_sc_hd__decap_3 PHY_284 ();
 sky130_fd_sc_hd__decap_3 PHY_285 ();
 sky130_fd_sc_hd__decap_3 PHY_286 ();
 sky130_fd_sc_hd__decap_3 PHY_287 ();
 sky130_fd_sc_hd__decap_3 PHY_288 ();
 sky130_fd_sc_hd__decap_3 PHY_289 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_290 ();
 sky130_fd_sc_hd__decap_3 PHY_291 ();
 sky130_fd_sc_hd__decap_3 PHY_292 ();
 sky130_fd_sc_hd__decap_3 PHY_293 ();
 sky130_fd_sc_hd__decap_3 PHY_294 ();
 sky130_fd_sc_hd__decap_3 PHY_295 ();
 sky130_fd_sc_hd__decap_3 PHY_296 ();
 sky130_fd_sc_hd__decap_3 PHY_297 ();
 sky130_fd_sc_hd__decap_3 PHY_298 ();
 sky130_fd_sc_hd__decap_3 PHY_299 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_300 ();
 sky130_fd_sc_hd__decap_3 PHY_301 ();
 sky130_fd_sc_hd__decap_3 PHY_302 ();
 sky130_fd_sc_hd__decap_3 PHY_303 ();
 sky130_fd_sc_hd__decap_3 PHY_304 ();
 sky130_fd_sc_hd__decap_3 PHY_305 ();
 sky130_fd_sc_hd__decap_3 PHY_306 ();
 sky130_fd_sc_hd__decap_3 PHY_307 ();
 sky130_fd_sc_hd__decap_3 PHY_308 ();
 sky130_fd_sc_hd__decap_3 PHY_309 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_310 ();
 sky130_fd_sc_hd__decap_3 PHY_311 ();
 sky130_fd_sc_hd__decap_3 PHY_312 ();
 sky130_fd_sc_hd__decap_3 PHY_313 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_999 ();
 sky130_fd_sc_hd__inv_2 _10790_ (.A(mstream_i),
    .Y(_02560_));
 sky130_fd_sc_hd__inv_2 _10791_ (.A(net598),
    .Y(_02561_));
 sky130_fd_sc_hd__clkinv_4 _10792_ (.A(sstream_i[114]),
    .Y(_02562_));
 sky130_fd_sc_hd__inv_2 _10793_ (.A(net510),
    .Y(_02563_));
 sky130_fd_sc_hd__inv_2 _10794_ (.A(net374),
    .Y(_02564_));
 sky130_fd_sc_hd__inv_2 _10795_ (.A(net628),
    .Y(_02565_));
 sky130_fd_sc_hd__inv_2 _10796_ (.A(net113),
    .Y(_02566_));
 sky130_fd_sc_hd__inv_2 _10797_ (.A(net326),
    .Y(_02567_));
 sky130_fd_sc_hd__inv_2 _10798_ (.A(net62),
    .Y(_02568_));
 sky130_fd_sc_hd__a21o_1 _10799_ (.A1(mstream_o[114]),
    .A2(_02560_),
    .B1(net619),
    .X(_00002_));
 sky130_fd_sc_hd__a22o_1 _10800_ (.A1(mstream_o[114]),
    .A2(mstream_i),
    .B1(sstream_o),
    .B2(_02562_),
    .X(_00001_));
 sky130_fd_sc_hd__and2_2 _10801_ (.A(sstream_o),
    .B(sstream_i[114]),
    .X(_00000_));
 sky130_fd_sc_hd__or2_1 _10802_ (.A(\add0.a_i[11] ),
    .B(\add0.b_i[11] ),
    .X(_02569_));
 sky130_fd_sc_hd__nand2_1 _10803_ (.A(\add0.a_i[11] ),
    .B(\add0.b_i[11] ),
    .Y(_02570_));
 sky130_fd_sc_hd__nand2_1 _10804_ (.A(\add0.a_i[10] ),
    .B(\add0.b_i[10] ),
    .Y(_02571_));
 sky130_fd_sc_hd__inv_2 _10805_ (.A(_02571_),
    .Y(_02572_));
 sky130_fd_sc_hd__or2_1 _10806_ (.A(\add0.a_i[10] ),
    .B(\add0.b_i[10] ),
    .X(_02573_));
 sky130_fd_sc_hd__nand2_1 _10807_ (.A(_02571_),
    .B(_02573_),
    .Y(_02574_));
 sky130_fd_sc_hd__nand2_1 _10808_ (.A(\add0.a_i[8] ),
    .B(\add0.b_i[8] ),
    .Y(_02575_));
 sky130_fd_sc_hd__or2_1 _10809_ (.A(\add0.a_i[8] ),
    .B(\add0.b_i[8] ),
    .X(_02576_));
 sky130_fd_sc_hd__nand2_2 _10810_ (.A(_02575_),
    .B(_02576_),
    .Y(_02577_));
 sky130_fd_sc_hd__nand2_1 _10811_ (.A(\add0.a_i[7] ),
    .B(\add0.b_i[7] ),
    .Y(_02578_));
 sky130_fd_sc_hd__or2_1 _10812_ (.A(\add0.a_i[7] ),
    .B(\add0.b_i[7] ),
    .X(_02579_));
 sky130_fd_sc_hd__nand2_1 _10813_ (.A(\add0.a_i[6] ),
    .B(\add0.b_i[6] ),
    .Y(_02580_));
 sky130_fd_sc_hd__or2_1 _10814_ (.A(\add0.a_i[6] ),
    .B(\add0.b_i[6] ),
    .X(_02581_));
 sky130_fd_sc_hd__nand2_2 _10815_ (.A(_02580_),
    .B(_02581_),
    .Y(_02582_));
 sky130_fd_sc_hd__and2_1 _10816_ (.A(\add0.a_i[5] ),
    .B(\add0.b_i[5] ),
    .X(_02583_));
 sky130_fd_sc_hd__nand2_1 _10817_ (.A(\add0.a_i[5] ),
    .B(\add0.b_i[5] ),
    .Y(_02584_));
 sky130_fd_sc_hd__nor2_2 _10818_ (.A(\add0.a_i[5] ),
    .B(\add0.b_i[5] ),
    .Y(_02585_));
 sky130_fd_sc_hd__nand2_1 _10819_ (.A(\add0.a_i[4] ),
    .B(\add0.b_i[4] ),
    .Y(_02586_));
 sky130_fd_sc_hd__or2_1 _10820_ (.A(\add0.a_i[4] ),
    .B(\add0.b_i[4] ),
    .X(_02587_));
 sky130_fd_sc_hd__nand2_2 _10821_ (.A(_02586_),
    .B(_02587_),
    .Y(_02588_));
 sky130_fd_sc_hd__and2_1 _10822_ (.A(\add0.a_i[3] ),
    .B(\add0.b_i[3] ),
    .X(_02589_));
 sky130_fd_sc_hd__nor2_1 _10823_ (.A(\add0.a_i[3] ),
    .B(\add0.b_i[3] ),
    .Y(_02590_));
 sky130_fd_sc_hd__and2_1 _10824_ (.A(\add0.a_i[2] ),
    .B(\add0.b_i[2] ),
    .X(_02591_));
 sky130_fd_sc_hd__nor2_1 _10825_ (.A(\add0.a_i[2] ),
    .B(\add0.b_i[2] ),
    .Y(_02592_));
 sky130_fd_sc_hd__nand2_1 _10826_ (.A(\add0.a_i[1] ),
    .B(\add0.b_i[1] ),
    .Y(_02593_));
 sky130_fd_sc_hd__nand2_2 _10827_ (.A(\add0.a_i[0] ),
    .B(\add0.b_i[0] ),
    .Y(_02594_));
 sky130_fd_sc_hd__nor2_1 _10828_ (.A(\add0.a_i[1] ),
    .B(\add0.b_i[1] ),
    .Y(_02595_));
 sky130_fd_sc_hd__or2_1 _10829_ (.A(\add0.a_i[1] ),
    .B(\add0.b_i[1] ),
    .X(_02596_));
 sky130_fd_sc_hd__nand2_2 _10830_ (.A(_02593_),
    .B(_02596_),
    .Y(_02597_));
 sky130_fd_sc_hd__o21a_2 _10831_ (.A1(_02594_),
    .A2(_02595_),
    .B1(_02593_),
    .X(_02598_));
 sky130_fd_sc_hd__o21ba_2 _10832_ (.A1(_02592_),
    .A2(_02598_),
    .B1_N(_02591_),
    .X(_02599_));
 sky130_fd_sc_hd__o21ba_2 _10833_ (.A1(_02590_),
    .A2(_02599_),
    .B1_N(_02589_),
    .X(_02600_));
 sky130_fd_sc_hd__o21a_2 _10834_ (.A1(_02588_),
    .A2(_02600_),
    .B1(_02586_),
    .X(_02601_));
 sky130_fd_sc_hd__nand3b_1 _10835_ (.A_N(_02585_),
    .B(\add0.b_i[4] ),
    .C(\add0.a_i[4] ),
    .Y(_02602_));
 sky130_fd_sc_hd__nor2_2 _10836_ (.A(_02583_),
    .B(_02585_),
    .Y(_02603_));
 sky130_fd_sc_hd__or3b_1 _10837_ (.A(_02588_),
    .B(_02600_),
    .C_N(_02603_),
    .X(_02604_));
 sky130_fd_sc_hd__o21ai_4 _10838_ (.A1(_02585_),
    .A2(_02601_),
    .B1(_02584_),
    .Y(_02605_));
 sky130_fd_sc_hd__a21bo_1 _10839_ (.A1(_02581_),
    .A2(_02605_),
    .B1_N(_02580_),
    .X(_02606_));
 sky130_fd_sc_hd__nand3_1 _10840_ (.A(\add0.a_i[6] ),
    .B(\add0.b_i[6] ),
    .C(_02579_),
    .Y(_02607_));
 sky130_fd_sc_hd__nand2_2 _10841_ (.A(_02578_),
    .B(_02579_),
    .Y(_02608_));
 sky130_fd_sc_hd__a311o_1 _10842_ (.A1(_02584_),
    .A2(_02602_),
    .A3(_02604_),
    .B1(_02608_),
    .C1(_02582_),
    .X(_02609_));
 sky130_fd_sc_hd__and3_2 _10843_ (.A(_02578_),
    .B(_02607_),
    .C(_02609_),
    .X(_02610_));
 sky130_fd_sc_hd__o21a_2 _10844_ (.A1(_02577_),
    .A2(_02610_),
    .B1(_02575_),
    .X(_02611_));
 sky130_fd_sc_hd__o211a_1 _10845_ (.A1(\add0.a_i[9] ),
    .A2(\add0.b_i[9] ),
    .B1(\add0.a_i[8] ),
    .C1(\add0.b_i[8] ),
    .X(_02612_));
 sky130_fd_sc_hd__a21oi_1 _10846_ (.A1(\add0.a_i[9] ),
    .A2(\add0.b_i[9] ),
    .B1(_02612_),
    .Y(_02613_));
 sky130_fd_sc_hd__xnor2_2 _10847_ (.A(\add0.a_i[9] ),
    .B(\add0.b_i[9] ),
    .Y(_02614_));
 sky130_fd_sc_hd__a311o_1 _10848_ (.A1(_02578_),
    .A2(_02607_),
    .A3(_02609_),
    .B1(_02614_),
    .C1(_02577_),
    .X(_02615_));
 sky130_fd_sc_hd__a21oi_2 _10849_ (.A1(_02613_),
    .A2(_02615_),
    .B1(_02574_),
    .Y(_02616_));
 sky130_fd_sc_hd__o211ai_2 _10850_ (.A1(_02572_),
    .A2(_02616_),
    .B1(_02569_),
    .C1(_02570_),
    .Y(_02617_));
 sky130_fd_sc_hd__a211o_1 _10851_ (.A1(_02569_),
    .A2(_02570_),
    .B1(_02572_),
    .C1(_02616_),
    .X(_02618_));
 sky130_fd_sc_hd__and2_2 _10852_ (.A(_02617_),
    .B(_02618_),
    .X(_02619_));
 sky130_fd_sc_hd__mux2_1 _10853_ (.A0(mstream_o[43]),
    .A1(_02619_),
    .S(net614),
    .X(_00003_));
 sky130_fd_sc_hd__or2_1 _10854_ (.A(\add0.a_i[12] ),
    .B(\add0.b_i[12] ),
    .X(_02620_));
 sky130_fd_sc_hd__nand2_1 _10855_ (.A(\add0.a_i[12] ),
    .B(\add0.b_i[12] ),
    .Y(_02621_));
 sky130_fd_sc_hd__inv_2 _10856_ (.A(_02621_),
    .Y(_02622_));
 sky130_fd_sc_hd__nand2_1 _10857_ (.A(_02620_),
    .B(_02621_),
    .Y(_02623_));
 sky130_fd_sc_hd__a21oi_2 _10858_ (.A1(_02570_),
    .A2(_02617_),
    .B1(_02623_),
    .Y(_02624_));
 sky130_fd_sc_hd__and3_1 _10859_ (.A(_02570_),
    .B(_02617_),
    .C(_02623_),
    .X(_02625_));
 sky130_fd_sc_hd__nor2_2 _10860_ (.A(_02624_),
    .B(_02625_),
    .Y(_02626_));
 sky130_fd_sc_hd__mux2_1 _10861_ (.A0(mstream_o[44]),
    .A1(_02626_),
    .S(net615),
    .X(_00004_));
 sky130_fd_sc_hd__or2_1 _10862_ (.A(\add0.a_i[13] ),
    .B(\add0.b_i[13] ),
    .X(_02627_));
 sky130_fd_sc_hd__nand2_1 _10863_ (.A(\add0.a_i[13] ),
    .B(\add0.b_i[13] ),
    .Y(_02628_));
 sky130_fd_sc_hd__nand2_1 _10864_ (.A(_02627_),
    .B(_02628_),
    .Y(_02629_));
 sky130_fd_sc_hd__o21bai_2 _10865_ (.A1(_02622_),
    .A2(_02624_),
    .B1_N(_02629_),
    .Y(_02630_));
 sky130_fd_sc_hd__or3b_1 _10866_ (.A(_02622_),
    .B(_02624_),
    .C_N(_02629_),
    .X(_02631_));
 sky130_fd_sc_hd__and2_2 _10867_ (.A(_02630_),
    .B(_02631_),
    .X(_02632_));
 sky130_fd_sc_hd__mux2_1 _10868_ (.A0(mstream_o[45]),
    .A1(_02632_),
    .S(net615),
    .X(_00005_));
 sky130_fd_sc_hd__nor2_1 _10869_ (.A(\add0.a_i[14] ),
    .B(\add0.b_i[14] ),
    .Y(_02633_));
 sky130_fd_sc_hd__and2_1 _10870_ (.A(\add0.a_i[14] ),
    .B(\add0.b_i[14] ),
    .X(_02634_));
 sky130_fd_sc_hd__or2_1 _10871_ (.A(_02633_),
    .B(_02634_),
    .X(_02635_));
 sky130_fd_sc_hd__a21oi_2 _10872_ (.A1(_02628_),
    .A2(_02630_),
    .B1(_02635_),
    .Y(_02636_));
 sky130_fd_sc_hd__and3_1 _10873_ (.A(_02628_),
    .B(_02630_),
    .C(_02635_),
    .X(_02637_));
 sky130_fd_sc_hd__nor2_4 _10874_ (.A(_02636_),
    .B(_02637_),
    .Y(_02638_));
 sky130_fd_sc_hd__mux2_1 _10875_ (.A0(mstream_o[46]),
    .A1(_02638_),
    .S(net615),
    .X(_00006_));
 sky130_fd_sc_hd__or2_1 _10876_ (.A(\add0.a_i[15] ),
    .B(\add0.b_i[15] ),
    .X(_02639_));
 sky130_fd_sc_hd__nand2_1 _10877_ (.A(\add0.a_i[15] ),
    .B(\add0.b_i[15] ),
    .Y(_02640_));
 sky130_fd_sc_hd__nand2_1 _10878_ (.A(_02639_),
    .B(_02640_),
    .Y(_02641_));
 sky130_fd_sc_hd__o21bai_2 _10879_ (.A1(_02634_),
    .A2(_02636_),
    .B1_N(_02641_),
    .Y(_02642_));
 sky130_fd_sc_hd__or3b_1 _10880_ (.A(_02634_),
    .B(_02636_),
    .C_N(_02641_),
    .X(_02643_));
 sky130_fd_sc_hd__and2_2 _10881_ (.A(_02642_),
    .B(_02643_),
    .X(_02644_));
 sky130_fd_sc_hd__mux2_1 _10882_ (.A0(mstream_o[47]),
    .A1(_02644_),
    .S(net615),
    .X(_00007_));
 sky130_fd_sc_hd__xnor2_1 _10883_ (.A(\add0.a_i[16] ),
    .B(\add0.b_i[16] ),
    .Y(_02645_));
 sky130_fd_sc_hd__a21oi_1 _10884_ (.A1(_02640_),
    .A2(_02642_),
    .B1(_02645_),
    .Y(_02646_));
 sky130_fd_sc_hd__and3_1 _10885_ (.A(_02640_),
    .B(_02642_),
    .C(_02645_),
    .X(_02647_));
 sky130_fd_sc_hd__nor2_2 _10886_ (.A(_02646_),
    .B(_02647_),
    .Y(_02648_));
 sky130_fd_sc_hd__mux2_1 _10887_ (.A0(mstream_o[48]),
    .A1(_02648_),
    .S(net615),
    .X(_00008_));
 sky130_fd_sc_hd__nor2_1 _10888_ (.A(\add0.a_i[17] ),
    .B(\add0.b_i[17] ),
    .Y(_02649_));
 sky130_fd_sc_hd__and2_1 _10889_ (.A(\add0.a_i[17] ),
    .B(\add0.b_i[17] ),
    .X(_02650_));
 sky130_fd_sc_hd__or2_2 _10890_ (.A(_02649_),
    .B(_02650_),
    .X(_02651_));
 sky130_fd_sc_hd__a21o_1 _10891_ (.A1(\add0.a_i[16] ),
    .A2(\add0.b_i[16] ),
    .B1(_02646_),
    .X(_02652_));
 sky130_fd_sc_hd__xnor2_4 _10892_ (.A(_02651_),
    .B(_02652_),
    .Y(_02653_));
 sky130_fd_sc_hd__mux2_1 _10893_ (.A0(mstream_o[49]),
    .A1(_02653_),
    .S(net615),
    .X(_00009_));
 sky130_fd_sc_hd__or2_1 _10894_ (.A(\add0.a_i[18] ),
    .B(\add0.b_i[18] ),
    .X(_02654_));
 sky130_fd_sc_hd__nand2_1 _10895_ (.A(\add0.a_i[18] ),
    .B(\add0.b_i[18] ),
    .Y(_02655_));
 sky130_fd_sc_hd__inv_2 _10896_ (.A(_02655_),
    .Y(_02656_));
 sky130_fd_sc_hd__nand2_1 _10897_ (.A(_02654_),
    .B(_02655_),
    .Y(_02657_));
 sky130_fd_sc_hd__o211a_1 _10898_ (.A1(\add0.a_i[17] ),
    .A2(\add0.b_i[17] ),
    .B1(\add0.a_i[16] ),
    .C1(\add0.b_i[16] ),
    .X(_02658_));
 sky130_fd_sc_hd__nor2_1 _10899_ (.A(_02650_),
    .B(_02658_),
    .Y(_02659_));
 sky130_fd_sc_hd__a211o_1 _10900_ (.A1(_02640_),
    .A2(_02642_),
    .B1(_02645_),
    .C1(_02651_),
    .X(_02660_));
 sky130_fd_sc_hd__a21oi_1 _10901_ (.A1(_02659_),
    .A2(_02660_),
    .B1(_02657_),
    .Y(_02661_));
 sky130_fd_sc_hd__and3_1 _10902_ (.A(_02657_),
    .B(_02659_),
    .C(_02660_),
    .X(_02662_));
 sky130_fd_sc_hd__nor2_2 _10903_ (.A(_02661_),
    .B(_02662_),
    .Y(_02663_));
 sky130_fd_sc_hd__mux2_1 _10904_ (.A0(mstream_o[50]),
    .A1(_02663_),
    .S(net615),
    .X(_00010_));
 sky130_fd_sc_hd__or2_1 _10905_ (.A(\add0.a_i[19] ),
    .B(\add0.b_i[19] ),
    .X(_02664_));
 sky130_fd_sc_hd__nand2_1 _10906_ (.A(\add0.a_i[19] ),
    .B(\add0.b_i[19] ),
    .Y(_02665_));
 sky130_fd_sc_hd__inv_2 _10907_ (.A(_02665_),
    .Y(_02666_));
 sky130_fd_sc_hd__nand2_1 _10908_ (.A(_02664_),
    .B(_02665_),
    .Y(_02667_));
 sky130_fd_sc_hd__inv_2 _10909_ (.A(_02667_),
    .Y(_02668_));
 sky130_fd_sc_hd__o21a_1 _10910_ (.A1(_02656_),
    .A2(_02661_),
    .B1(_02668_),
    .X(_02669_));
 sky130_fd_sc_hd__or3_1 _10911_ (.A(_02656_),
    .B(_02661_),
    .C(_02668_),
    .X(_02670_));
 sky130_fd_sc_hd__and2b_2 _10912_ (.A_N(_02669_),
    .B(_02670_),
    .X(_02671_));
 sky130_fd_sc_hd__mux2_1 _10913_ (.A0(mstream_o[51]),
    .A1(_02671_),
    .S(net615),
    .X(_00011_));
 sky130_fd_sc_hd__nor2_1 _10914_ (.A(\add0.a_i[20] ),
    .B(\add0.b_i[20] ),
    .Y(_02672_));
 sky130_fd_sc_hd__and2_1 _10915_ (.A(\add0.a_i[20] ),
    .B(\add0.b_i[20] ),
    .X(_02673_));
 sky130_fd_sc_hd__or2_2 _10916_ (.A(_02672_),
    .B(_02673_),
    .X(_02674_));
 sky130_fd_sc_hd__nor2_2 _10917_ (.A(_02666_),
    .B(_02669_),
    .Y(_02675_));
 sky130_fd_sc_hd__o21ba_1 _10918_ (.A1(_02666_),
    .A2(_02669_),
    .B1_N(_02674_),
    .X(_02676_));
 sky130_fd_sc_hd__xor2_4 _10919_ (.A(_02674_),
    .B(_02675_),
    .X(_02677_));
 sky130_fd_sc_hd__mux2_1 _10920_ (.A0(mstream_o[52]),
    .A1(_02677_),
    .S(net615),
    .X(_00012_));
 sky130_fd_sc_hd__or2_1 _10921_ (.A(\add0.a_i[21] ),
    .B(\add0.b_i[21] ),
    .X(_02678_));
 sky130_fd_sc_hd__nand2_1 _10922_ (.A(\add0.a_i[21] ),
    .B(\add0.b_i[21] ),
    .Y(_02679_));
 sky130_fd_sc_hd__nand2_2 _10923_ (.A(_02678_),
    .B(_02679_),
    .Y(_02680_));
 sky130_fd_sc_hd__nor2_2 _10924_ (.A(_02673_),
    .B(_02676_),
    .Y(_02681_));
 sky130_fd_sc_hd__o21bai_1 _10925_ (.A1(_02673_),
    .A2(_02676_),
    .B1_N(_02680_),
    .Y(_02682_));
 sky130_fd_sc_hd__xor2_4 _10926_ (.A(_02680_),
    .B(_02681_),
    .X(_02683_));
 sky130_fd_sc_hd__mux2_1 _10927_ (.A0(mstream_o[53]),
    .A1(_02683_),
    .S(net615),
    .X(_00013_));
 sky130_fd_sc_hd__or2_1 _10928_ (.A(\add0.a_i[22] ),
    .B(\add0.b_i[22] ),
    .X(_02684_));
 sky130_fd_sc_hd__nand2_1 _10929_ (.A(\add0.a_i[22] ),
    .B(\add0.b_i[22] ),
    .Y(_02685_));
 sky130_fd_sc_hd__inv_2 _10930_ (.A(_02685_),
    .Y(_02686_));
 sky130_fd_sc_hd__nand2_1 _10931_ (.A(_02684_),
    .B(_02685_),
    .Y(_02687_));
 sky130_fd_sc_hd__a21oi_2 _10932_ (.A1(_02679_),
    .A2(_02682_),
    .B1(_02687_),
    .Y(_02688_));
 sky130_fd_sc_hd__o211a_1 _10933_ (.A1(_02680_),
    .A2(_02681_),
    .B1(_02687_),
    .C1(_02679_),
    .X(_02689_));
 sky130_fd_sc_hd__nor2_2 _10934_ (.A(_02688_),
    .B(_02689_),
    .Y(_02690_));
 sky130_fd_sc_hd__mux2_1 _10935_ (.A0(mstream_o[54]),
    .A1(_02690_),
    .S(net615),
    .X(_00014_));
 sky130_fd_sc_hd__or2_1 _10936_ (.A(\add0.a_i[23] ),
    .B(\add0.b_i[23] ),
    .X(_02691_));
 sky130_fd_sc_hd__nand2_1 _10937_ (.A(\add0.a_i[23] ),
    .B(\add0.b_i[23] ),
    .Y(_02692_));
 sky130_fd_sc_hd__nand2_1 _10938_ (.A(_02691_),
    .B(_02692_),
    .Y(_02693_));
 sky130_fd_sc_hd__o21bai_2 _10939_ (.A1(_02686_),
    .A2(_02688_),
    .B1_N(_02693_),
    .Y(_02694_));
 sky130_fd_sc_hd__or3b_1 _10940_ (.A(_02686_),
    .B(_02688_),
    .C_N(_02693_),
    .X(_02695_));
 sky130_fd_sc_hd__and2_2 _10941_ (.A(_02694_),
    .B(_02695_),
    .X(_02696_));
 sky130_fd_sc_hd__mux2_1 _10942_ (.A0(mstream_o[55]),
    .A1(_02696_),
    .S(net615),
    .X(_00015_));
 sky130_fd_sc_hd__xnor2_1 _10943_ (.A(\add0.a_i[24] ),
    .B(\add0.b_i[24] ),
    .Y(_02697_));
 sky130_fd_sc_hd__a21oi_1 _10944_ (.A1(_02692_),
    .A2(_02694_),
    .B1(_02697_),
    .Y(_02698_));
 sky130_fd_sc_hd__and3_1 _10945_ (.A(_02692_),
    .B(_02694_),
    .C(_02697_),
    .X(_02699_));
 sky130_fd_sc_hd__nor2_2 _10946_ (.A(_02698_),
    .B(_02699_),
    .Y(_02700_));
 sky130_fd_sc_hd__mux2_1 _10947_ (.A0(mstream_o[56]),
    .A1(_02700_),
    .S(net616),
    .X(_00016_));
 sky130_fd_sc_hd__xnor2_4 _10948_ (.A(\add0.a_i[25] ),
    .B(\add0.b_i[25] ),
    .Y(_02701_));
 sky130_fd_sc_hd__a21o_1 _10949_ (.A1(\add0.a_i[24] ),
    .A2(\add0.b_i[24] ),
    .B1(_02698_),
    .X(_02702_));
 sky130_fd_sc_hd__xnor2_4 _10950_ (.A(_02701_),
    .B(_02702_),
    .Y(_02703_));
 sky130_fd_sc_hd__mux2_1 _10951_ (.A0(mstream_o[57]),
    .A1(_02703_),
    .S(net615),
    .X(_00017_));
 sky130_fd_sc_hd__o211a_1 _10952_ (.A1(\add0.a_i[25] ),
    .A2(\add0.b_i[25] ),
    .B1(\add0.a_i[24] ),
    .C1(\add0.b_i[24] ),
    .X(_02704_));
 sky130_fd_sc_hd__a211oi_1 _10953_ (.A1(_02692_),
    .A2(_02694_),
    .B1(_02697_),
    .C1(_02701_),
    .Y(_02705_));
 sky130_fd_sc_hd__a211o_2 _10954_ (.A1(\add0.a_i[25] ),
    .A2(\add0.b_i[25] ),
    .B1(_02704_),
    .C1(_02705_),
    .X(_02706_));
 sky130_fd_sc_hd__and2_1 _10955_ (.A(\add0.a_i[26] ),
    .B(\add0.b_i[26] ),
    .X(_02707_));
 sky130_fd_sc_hd__nor2_1 _10956_ (.A(\add0.a_i[26] ),
    .B(\add0.b_i[26] ),
    .Y(_02708_));
 sky130_fd_sc_hd__or2_2 _10957_ (.A(_02707_),
    .B(_02708_),
    .X(_02709_));
 sky130_fd_sc_hd__inv_2 _10958_ (.A(_02709_),
    .Y(_02710_));
 sky130_fd_sc_hd__xnor2_4 _10959_ (.A(_02706_),
    .B(_02709_),
    .Y(_02711_));
 sky130_fd_sc_hd__mux2_1 _10960_ (.A0(mstream_o[58]),
    .A1(_02711_),
    .S(net615),
    .X(_00018_));
 sky130_fd_sc_hd__and2_1 _10961_ (.A(\add0.a_i[27] ),
    .B(\add0.b_i[27] ),
    .X(_02712_));
 sky130_fd_sc_hd__or2_1 _10962_ (.A(\add0.a_i[27] ),
    .B(\add0.b_i[27] ),
    .X(_02713_));
 sky130_fd_sc_hd__and2b_1 _10963_ (.A_N(_02712_),
    .B(_02713_),
    .X(_02714_));
 sky130_fd_sc_hd__a21oi_2 _10964_ (.A1(_02706_),
    .A2(_02710_),
    .B1(_02707_),
    .Y(_02715_));
 sky130_fd_sc_hd__xnor2_4 _10965_ (.A(_02714_),
    .B(_02715_),
    .Y(_02716_));
 sky130_fd_sc_hd__mux2_1 _10966_ (.A0(mstream_o[59]),
    .A1(_02716_),
    .S(net617),
    .X(_00019_));
 sky130_fd_sc_hd__and3_1 _10967_ (.A(\add0.a_i[26] ),
    .B(\add0.b_i[26] ),
    .C(_02713_),
    .X(_02717_));
 sky130_fd_sc_hd__a311o_2 _10968_ (.A1(_02706_),
    .A2(_02710_),
    .A3(_02713_),
    .B1(_02717_),
    .C1(_02712_),
    .X(_02718_));
 sky130_fd_sc_hd__or2_1 _10969_ (.A(\add0.a_i[28] ),
    .B(\add0.b_i[28] ),
    .X(_02719_));
 sky130_fd_sc_hd__nand2_1 _10970_ (.A(\add0.a_i[28] ),
    .B(\add0.b_i[28] ),
    .Y(_02720_));
 sky130_fd_sc_hd__nand2_2 _10971_ (.A(_02719_),
    .B(_02720_),
    .Y(_02721_));
 sky130_fd_sc_hd__xnor2_4 _10972_ (.A(_02718_),
    .B(_02721_),
    .Y(_02722_));
 sky130_fd_sc_hd__mux2_1 _10973_ (.A0(mstream_o[60]),
    .A1(_02722_),
    .S(net617),
    .X(_00020_));
 sky130_fd_sc_hd__a21bo_2 _10974_ (.A1(_02718_),
    .A2(_02719_),
    .B1_N(_02720_),
    .X(_02723_));
 sky130_fd_sc_hd__or2_1 _10975_ (.A(\add0.a_i[29] ),
    .B(\add0.b_i[29] ),
    .X(_02724_));
 sky130_fd_sc_hd__nand2_1 _10976_ (.A(\add0.a_i[29] ),
    .B(\add0.b_i[29] ),
    .Y(_02725_));
 sky130_fd_sc_hd__nand2_2 _10977_ (.A(_02724_),
    .B(_02725_),
    .Y(_02726_));
 sky130_fd_sc_hd__xnor2_4 _10978_ (.A(_02723_),
    .B(_02726_),
    .Y(_02727_));
 sky130_fd_sc_hd__mux2_1 _10979_ (.A0(mstream_o[61]),
    .A1(_02727_),
    .S(net617),
    .X(_00021_));
 sky130_fd_sc_hd__or2_1 _10980_ (.A(\add0.a_i[30] ),
    .B(\add0.b_i[30] ),
    .X(_02728_));
 sky130_fd_sc_hd__nand2_1 _10981_ (.A(\add0.a_i[30] ),
    .B(\add0.b_i[30] ),
    .Y(_02729_));
 sky130_fd_sc_hd__nand2_2 _10982_ (.A(_02728_),
    .B(_02729_),
    .Y(_02730_));
 sky130_fd_sc_hd__a21bo_2 _10983_ (.A1(_02723_),
    .A2(_02724_),
    .B1_N(_02725_),
    .X(_02731_));
 sky130_fd_sc_hd__xnor2_4 _10984_ (.A(_02730_),
    .B(_02731_),
    .Y(_02732_));
 sky130_fd_sc_hd__mux2_1 _10985_ (.A0(mstream_o[62]),
    .A1(_02732_),
    .S(net617),
    .X(_00022_));
 sky130_fd_sc_hd__a21bo_1 _10986_ (.A1(_02728_),
    .A2(_02731_),
    .B1_N(_02729_),
    .X(_02733_));
 sky130_fd_sc_hd__xnor2_2 _10987_ (.A(\add0.a_i[31] ),
    .B(\add0.b_i[31] ),
    .Y(_02734_));
 sky130_fd_sc_hd__xnor2_4 _10988_ (.A(_02733_),
    .B(_02734_),
    .Y(_02735_));
 sky130_fd_sc_hd__mux2_1 _10989_ (.A0(mstream_o[63]),
    .A1(_02735_),
    .S(net617),
    .X(_00023_));
 sky130_fd_sc_hd__mux2_1 _10990_ (.A0(mstream_o[64]),
    .A1(net705),
    .S(net615),
    .X(_00024_));
 sky130_fd_sc_hd__mux2_1 _10991_ (.A0(mstream_o[65]),
    .A1(net718),
    .S(net616),
    .X(_00025_));
 sky130_fd_sc_hd__mux2_1 _10992_ (.A0(mstream_o[66]),
    .A1(net789),
    .S(net615),
    .X(_00026_));
 sky130_fd_sc_hd__mux2_1 _10993_ (.A0(mstream_o[67]),
    .A1(net657),
    .S(net617),
    .X(_00027_));
 sky130_fd_sc_hd__mux2_1 _10994_ (.A0(mstream_o[68]),
    .A1(net732),
    .S(net617),
    .X(_00028_));
 sky130_fd_sc_hd__mux2_1 _10995_ (.A0(mstream_o[69]),
    .A1(net711),
    .S(net617),
    .X(_00029_));
 sky130_fd_sc_hd__mux2_1 _10996_ (.A0(mstream_o[70]),
    .A1(net688),
    .S(net617),
    .X(_00030_));
 sky130_fd_sc_hd__mux2_1 _10997_ (.A0(mstream_o[71]),
    .A1(net712),
    .S(net617),
    .X(_00031_));
 sky130_fd_sc_hd__mux2_1 _10998_ (.A0(mstream_o[72]),
    .A1(net686),
    .S(net617),
    .X(_00032_));
 sky130_fd_sc_hd__mux2_1 _10999_ (.A0(mstream_o[73]),
    .A1(net671),
    .S(net617),
    .X(_00033_));
 sky130_fd_sc_hd__mux2_1 _11000_ (.A0(mstream_o[74]),
    .A1(net727),
    .S(net617),
    .X(_00034_));
 sky130_fd_sc_hd__mux2_1 _11001_ (.A0(mstream_o[75]),
    .A1(net673),
    .S(net618),
    .X(_00035_));
 sky130_fd_sc_hd__mux2_1 _11002_ (.A0(mstream_o[76]),
    .A1(net701),
    .S(net618),
    .X(_00036_));
 sky130_fd_sc_hd__mux2_1 _11003_ (.A0(mstream_o[77]),
    .A1(net745),
    .S(net617),
    .X(_00037_));
 sky130_fd_sc_hd__mux2_1 _11004_ (.A0(mstream_o[78]),
    .A1(net656),
    .S(net617),
    .X(_00038_));
 sky130_fd_sc_hd__mux2_1 _11005_ (.A0(mstream_o[79]),
    .A1(net670),
    .S(net617),
    .X(_00039_));
 sky130_fd_sc_hd__mux2_1 _11006_ (.A0(mstream_o[80]),
    .A1(net714),
    .S(net618),
    .X(_00040_));
 sky130_fd_sc_hd__mux2_1 _11007_ (.A0(mstream_o[81]),
    .A1(net694),
    .S(net618),
    .X(_00041_));
 sky130_fd_sc_hd__mux2_1 _11008_ (.A0(mstream_o[82]),
    .A1(net716),
    .S(net618),
    .X(_00042_));
 sky130_fd_sc_hd__mux2_1 _11009_ (.A0(mstream_o[83]),
    .A1(net715),
    .S(net618),
    .X(_00043_));
 sky130_fd_sc_hd__mux2_1 _11010_ (.A0(mstream_o[84]),
    .A1(net660),
    .S(net618),
    .X(_00044_));
 sky130_fd_sc_hd__mux2_1 _11011_ (.A0(mstream_o[85]),
    .A1(net698),
    .S(net618),
    .X(_00045_));
 sky130_fd_sc_hd__mux2_1 _11012_ (.A0(mstream_o[86]),
    .A1(net664),
    .S(net618),
    .X(_00046_));
 sky130_fd_sc_hd__mux2_1 _11013_ (.A0(mstream_o[87]),
    .A1(net653),
    .S(net619),
    .X(_00047_));
 sky130_fd_sc_hd__mux2_1 _11014_ (.A0(mstream_o[88]),
    .A1(net717),
    .S(net619),
    .X(_00048_));
 sky130_fd_sc_hd__mux2_1 _11015_ (.A0(mstream_o[89]),
    .A1(net708),
    .S(net619),
    .X(_00049_));
 sky130_fd_sc_hd__mux2_1 _11016_ (.A0(mstream_o[90]),
    .A1(net649),
    .S(net619),
    .X(_00050_));
 sky130_fd_sc_hd__mux2_1 _11017_ (.A0(mstream_o[91]),
    .A1(net702),
    .S(net619),
    .X(_00051_));
 sky130_fd_sc_hd__mux2_1 _11018_ (.A0(mstream_o[92]),
    .A1(net690),
    .S(net619),
    .X(_00052_));
 sky130_fd_sc_hd__mux2_1 _11019_ (.A0(mstream_o[93]),
    .A1(net687),
    .S(net619),
    .X(_00053_));
 sky130_fd_sc_hd__mux2_1 _11020_ (.A0(mstream_o[94]),
    .A1(net692),
    .S(net619),
    .X(_00054_));
 sky130_fd_sc_hd__mux2_1 _11021_ (.A0(mstream_o[95]),
    .A1(net652),
    .S(net619),
    .X(_00055_));
 sky130_fd_sc_hd__mux2_1 _11022_ (.A0(mstream_o[96]),
    .A1(net880),
    .S(net619),
    .X(_00056_));
 sky130_fd_sc_hd__mux2_1 _11023_ (.A0(mstream_o[97]),
    .A1(net904),
    .S(net619),
    .X(_00057_));
 sky130_fd_sc_hd__mux2_1 _11024_ (.A0(mstream_o[98]),
    .A1(net885),
    .S(net619),
    .X(_00058_));
 sky130_fd_sc_hd__mux2_1 _11025_ (.A0(mstream_o[99]),
    .A1(net902),
    .S(net619),
    .X(_00059_));
 sky130_fd_sc_hd__mux2_1 _11026_ (.A0(mstream_o[100]),
    .A1(net936),
    .S(net619),
    .X(_00060_));
 sky130_fd_sc_hd__mux2_1 _11027_ (.A0(mstream_o[101]),
    .A1(net893),
    .S(net619),
    .X(_00061_));
 sky130_fd_sc_hd__mux2_1 _11028_ (.A0(mstream_o[102]),
    .A1(net921),
    .S(net620),
    .X(_00062_));
 sky130_fd_sc_hd__mux2_1 _11029_ (.A0(mstream_o[103]),
    .A1(net955),
    .S(net620),
    .X(_00063_));
 sky130_fd_sc_hd__mux2_1 _11030_ (.A0(mstream_o[104]),
    .A1(net932),
    .S(net620),
    .X(_00064_));
 sky130_fd_sc_hd__mux2_1 _11031_ (.A0(mstream_o[105]),
    .A1(net916),
    .S(net620),
    .X(_00065_));
 sky130_fd_sc_hd__mux2_1 _11032_ (.A0(mstream_o[106]),
    .A1(net945),
    .S(net620),
    .X(_00066_));
 sky130_fd_sc_hd__mux2_1 _11033_ (.A0(mstream_o[107]),
    .A1(net934),
    .S(net620),
    .X(_00067_));
 sky130_fd_sc_hd__mux2_1 _11034_ (.A0(mstream_o[108]),
    .A1(net920),
    .S(net620),
    .X(_00068_));
 sky130_fd_sc_hd__mux2_1 _11035_ (.A0(mstream_o[109]),
    .A1(net908),
    .S(net620),
    .X(_00069_));
 sky130_fd_sc_hd__mux2_1 _11036_ (.A0(mstream_o[110]),
    .A1(net952),
    .S(net620),
    .X(_00070_));
 sky130_fd_sc_hd__mux2_1 _11037_ (.A0(mstream_o[111]),
    .A1(net914),
    .S(net620),
    .X(_00071_));
 sky130_fd_sc_hd__mux2_1 _11038_ (.A0(mstream_o[112]),
    .A1(net923),
    .S(net620),
    .X(_00072_));
 sky130_fd_sc_hd__mux2_1 _11039_ (.A0(mstream_o[113]),
    .A1(net929),
    .S(net620),
    .X(_00073_));
 sky130_fd_sc_hd__mux2_1 _11040_ (.A0(mstream_o[115]),
    .A1(sstream_i[115]),
    .S(_00000_),
    .X(_00074_));
 sky130_fd_sc_hd__nand2_2 _11041_ (.A(net642),
    .B(net599),
    .Y(_02736_));
 sky130_fd_sc_hd__or2_1 _11042_ (.A(\add0.a_i[0] ),
    .B(\add0.b_i[0] ),
    .X(_02737_));
 sky130_fd_sc_hd__and2_2 _11043_ (.A(_02594_),
    .B(_02737_),
    .X(_02738_));
 sky130_fd_sc_hd__mux2_1 _11044_ (.A0(_02738_),
    .A1(net705),
    .S(net55),
    .X(_00075_));
 sky130_fd_sc_hd__xor2_4 _11045_ (.A(_02594_),
    .B(_02597_),
    .X(_02739_));
 sky130_fd_sc_hd__mux2_1 _11046_ (.A0(_02739_),
    .A1(net718),
    .S(net55),
    .X(_00076_));
 sky130_fd_sc_hd__nor2_2 _11047_ (.A(_02591_),
    .B(_02592_),
    .Y(_02740_));
 sky130_fd_sc_hd__xnor2_4 _11048_ (.A(_02598_),
    .B(_02740_),
    .Y(_02741_));
 sky130_fd_sc_hd__mux2_1 _11049_ (.A0(_02741_),
    .A1(net789),
    .S(net55),
    .X(_00077_));
 sky130_fd_sc_hd__nor2_2 _11050_ (.A(_02589_),
    .B(_02590_),
    .Y(_02742_));
 sky130_fd_sc_hd__xnor2_4 _11051_ (.A(_02599_),
    .B(_02742_),
    .Y(_02743_));
 sky130_fd_sc_hd__mux2_1 _11052_ (.A0(_02743_),
    .A1(net657),
    .S(net55),
    .X(_00078_));
 sky130_fd_sc_hd__xor2_4 _11053_ (.A(_02588_),
    .B(_02600_),
    .X(_02744_));
 sky130_fd_sc_hd__mux2_1 _11054_ (.A0(_02744_),
    .A1(net732),
    .S(net55),
    .X(_00079_));
 sky130_fd_sc_hd__xnor2_4 _11055_ (.A(_02601_),
    .B(_02603_),
    .Y(_02745_));
 sky130_fd_sc_hd__mux2_1 _11056_ (.A0(_02745_),
    .A1(net711),
    .S(net55),
    .X(_00080_));
 sky130_fd_sc_hd__xnor2_4 _11057_ (.A(_02582_),
    .B(_02605_),
    .Y(_02746_));
 sky130_fd_sc_hd__mux2_1 _11058_ (.A0(_02746_),
    .A1(net688),
    .S(net55),
    .X(_00081_));
 sky130_fd_sc_hd__xnor2_4 _11059_ (.A(_02606_),
    .B(_02608_),
    .Y(_02747_));
 sky130_fd_sc_hd__mux2_1 _11060_ (.A0(_02747_),
    .A1(net712),
    .S(net55),
    .X(_00082_));
 sky130_fd_sc_hd__xor2_4 _11061_ (.A(_02577_),
    .B(_02610_),
    .X(_02748_));
 sky130_fd_sc_hd__mux2_1 _11062_ (.A0(_02748_),
    .A1(net686),
    .S(net55),
    .X(_00083_));
 sky130_fd_sc_hd__xor2_4 _11063_ (.A(_02611_),
    .B(_02614_),
    .X(_02749_));
 sky130_fd_sc_hd__mux2_1 _11064_ (.A0(_02749_),
    .A1(net671),
    .S(net55),
    .X(_00084_));
 sky130_fd_sc_hd__and3_1 _11065_ (.A(_02574_),
    .B(_02613_),
    .C(_02615_),
    .X(_02750_));
 sky130_fd_sc_hd__nor2_4 _11066_ (.A(_02616_),
    .B(_02750_),
    .Y(_02751_));
 sky130_fd_sc_hd__mux2_1 _11067_ (.A0(_02751_),
    .A1(net727),
    .S(net55),
    .X(_00085_));
 sky130_fd_sc_hd__mux2_1 _11068_ (.A0(_02619_),
    .A1(net673),
    .S(net54),
    .X(_00086_));
 sky130_fd_sc_hd__mux2_1 _11069_ (.A0(_02626_),
    .A1(net701),
    .S(net54),
    .X(_00087_));
 sky130_fd_sc_hd__mux2_1 _11070_ (.A0(_02632_),
    .A1(net745),
    .S(net54),
    .X(_00088_));
 sky130_fd_sc_hd__mux2_1 _11071_ (.A0(_02638_),
    .A1(net656),
    .S(net54),
    .X(_00089_));
 sky130_fd_sc_hd__mux2_1 _11072_ (.A0(_02644_),
    .A1(net670),
    .S(net54),
    .X(_00090_));
 sky130_fd_sc_hd__mux2_1 _11073_ (.A0(_02648_),
    .A1(net714),
    .S(net54),
    .X(_00091_));
 sky130_fd_sc_hd__mux2_1 _11074_ (.A0(_02653_),
    .A1(net694),
    .S(net54),
    .X(_00092_));
 sky130_fd_sc_hd__mux2_1 _11075_ (.A0(_02663_),
    .A1(net716),
    .S(net54),
    .X(_00093_));
 sky130_fd_sc_hd__mux2_1 _11076_ (.A0(_02671_),
    .A1(net715),
    .S(net54),
    .X(_00094_));
 sky130_fd_sc_hd__mux2_1 _11077_ (.A0(_02677_),
    .A1(net660),
    .S(net54),
    .X(_00095_));
 sky130_fd_sc_hd__mux2_1 _11078_ (.A0(_02683_),
    .A1(net698),
    .S(net55),
    .X(_00096_));
 sky130_fd_sc_hd__mux2_1 _11079_ (.A0(_02690_),
    .A1(net664),
    .S(net54),
    .X(_00097_));
 sky130_fd_sc_hd__mux2_1 _11080_ (.A0(_02696_),
    .A1(net653),
    .S(net54),
    .X(_00098_));
 sky130_fd_sc_hd__mux2_1 _11081_ (.A0(_02700_),
    .A1(net717),
    .S(net54),
    .X(_00099_));
 sky130_fd_sc_hd__mux2_1 _11082_ (.A0(_02703_),
    .A1(net708),
    .S(net54),
    .X(_00100_));
 sky130_fd_sc_hd__mux2_1 _11083_ (.A0(_02711_),
    .A1(net649),
    .S(net54),
    .X(_00101_));
 sky130_fd_sc_hd__mux2_1 _11084_ (.A0(_02716_),
    .A1(net702),
    .S(_02736_),
    .X(_00102_));
 sky130_fd_sc_hd__mux2_1 _11085_ (.A0(_02722_),
    .A1(net690),
    .S(net55),
    .X(_00103_));
 sky130_fd_sc_hd__mux2_1 _11086_ (.A0(_02727_),
    .A1(net687),
    .S(net55),
    .X(_00104_));
 sky130_fd_sc_hd__mux2_1 _11087_ (.A0(_02732_),
    .A1(net692),
    .S(net55),
    .X(_00105_));
 sky130_fd_sc_hd__mux2_1 _11088_ (.A0(_02735_),
    .A1(net652),
    .S(net54),
    .X(_00106_));
 sky130_fd_sc_hd__nand2_1 _11089_ (.A(net638),
    .B(net611),
    .Y(_02752_));
 sky130_fd_sc_hd__mux2_1 _11090_ (.A0(_02738_),
    .A1(net659),
    .S(net52),
    .X(_00107_));
 sky130_fd_sc_hd__mux2_1 _11091_ (.A0(_02739_),
    .A1(net655),
    .S(net52),
    .X(_00108_));
 sky130_fd_sc_hd__mux2_1 _11092_ (.A0(_02741_),
    .A1(net731),
    .S(net52),
    .X(_00109_));
 sky130_fd_sc_hd__mux2_1 _11093_ (.A0(_02743_),
    .A1(net667),
    .S(net52),
    .X(_00110_));
 sky130_fd_sc_hd__mux2_1 _11094_ (.A0(_02744_),
    .A1(net650),
    .S(net52),
    .X(_00111_));
 sky130_fd_sc_hd__mux2_1 _11095_ (.A0(_02745_),
    .A1(net661),
    .S(net52),
    .X(_00112_));
 sky130_fd_sc_hd__mux2_1 _11096_ (.A0(_02746_),
    .A1(net662),
    .S(net52),
    .X(_00113_));
 sky130_fd_sc_hd__mux2_1 _11097_ (.A0(_02747_),
    .A1(net665),
    .S(net52),
    .X(_00114_));
 sky130_fd_sc_hd__mux2_1 _11098_ (.A0(_02748_),
    .A1(net679),
    .S(net52),
    .X(_00115_));
 sky130_fd_sc_hd__mux2_1 _11099_ (.A0(_02749_),
    .A1(net819),
    .S(net52),
    .X(_00116_));
 sky130_fd_sc_hd__mux2_1 _11100_ (.A0(_02751_),
    .A1(net728),
    .S(net52),
    .X(_00117_));
 sky130_fd_sc_hd__mux2_1 _11101_ (.A0(_02619_),
    .A1(net695),
    .S(net52),
    .X(_00118_));
 sky130_fd_sc_hd__mux2_1 _11102_ (.A0(_02626_),
    .A1(net798),
    .S(net52),
    .X(_00119_));
 sky130_fd_sc_hd__mux2_1 _11103_ (.A0(_02632_),
    .A1(net677),
    .S(net52),
    .X(_00120_));
 sky130_fd_sc_hd__mux2_1 _11104_ (.A0(_02638_),
    .A1(net654),
    .S(net53),
    .X(_00121_));
 sky130_fd_sc_hd__mux2_1 _11105_ (.A0(_02644_),
    .A1(net752),
    .S(net53),
    .X(_00122_));
 sky130_fd_sc_hd__mux2_1 _11106_ (.A0(_02648_),
    .A1(net719),
    .S(net53),
    .X(_00123_));
 sky130_fd_sc_hd__mux2_1 _11107_ (.A0(_02653_),
    .A1(net678),
    .S(net52),
    .X(_00124_));
 sky130_fd_sc_hd__mux2_1 _11108_ (.A0(_02663_),
    .A1(net663),
    .S(net52),
    .X(_00125_));
 sky130_fd_sc_hd__mux2_1 _11109_ (.A0(_02671_),
    .A1(net790),
    .S(net53),
    .X(_00126_));
 sky130_fd_sc_hd__mux2_1 _11110_ (.A0(_02677_),
    .A1(net710),
    .S(net53),
    .X(_00127_));
 sky130_fd_sc_hd__mux2_1 _11111_ (.A0(_02683_),
    .A1(net672),
    .S(net53),
    .X(_00128_));
 sky130_fd_sc_hd__mux2_1 _11112_ (.A0(_02690_),
    .A1(net814),
    .S(_02752_),
    .X(_00129_));
 sky130_fd_sc_hd__mux2_1 _11113_ (.A0(_02696_),
    .A1(net700),
    .S(net53),
    .X(_00130_));
 sky130_fd_sc_hd__mux2_1 _11114_ (.A0(_02700_),
    .A1(net689),
    .S(net53),
    .X(_00131_));
 sky130_fd_sc_hd__mux2_1 _11115_ (.A0(_02703_),
    .A1(net674),
    .S(net53),
    .X(_00132_));
 sky130_fd_sc_hd__mux2_1 _11116_ (.A0(_02711_),
    .A1(net658),
    .S(net53),
    .X(_00133_));
 sky130_fd_sc_hd__mux2_1 _11117_ (.A0(_02716_),
    .A1(net691),
    .S(net53),
    .X(_00134_));
 sky130_fd_sc_hd__mux2_1 _11118_ (.A0(_02722_),
    .A1(net651),
    .S(net53),
    .X(_00135_));
 sky130_fd_sc_hd__mux2_1 _11119_ (.A0(_02727_),
    .A1(net707),
    .S(net53),
    .X(_00136_));
 sky130_fd_sc_hd__mux2_1 _11120_ (.A0(_02732_),
    .A1(net699),
    .S(net53),
    .X(_00137_));
 sky130_fd_sc_hd__mux2_1 _11121_ (.A0(_02735_),
    .A1(net713),
    .S(net53),
    .X(_00138_));
 sky130_fd_sc_hd__or2_2 _11122_ (.A(net598),
    .B(net601),
    .X(_02753_));
 sky130_fd_sc_hd__or2_1 _11123_ (.A(net607),
    .B(\state[5] ),
    .X(_02754_));
 sky130_fd_sc_hd__nor2_2 _11124_ (.A(net585),
    .B(net46),
    .Y(_02755_));
 sky130_fd_sc_hd__o31a_4 _11125_ (.A1(net585),
    .A2(net50),
    .A3(net46),
    .B1(net646),
    .X(_02756_));
 sky130_fd_sc_hd__nor2_2 _11126_ (.A(net50),
    .B(net46),
    .Y(_02757_));
 sky130_fd_sc_hd__a22o_1 _11127_ (.A1(net871),
    .A2(net50),
    .B1(net46),
    .B2(net846),
    .X(_02758_));
 sky130_fd_sc_hd__a21o_1 _11128_ (.A1(net806),
    .A2(net23),
    .B1(_02758_),
    .X(_02759_));
 sky130_fd_sc_hd__mux2_1 _11129_ (.A0(net582),
    .A1(_02759_),
    .S(net25),
    .X(_00139_));
 sky130_fd_sc_hd__a22o_1 _11130_ (.A1(net870),
    .A2(net50),
    .B1(net46),
    .B2(net843),
    .X(_02760_));
 sky130_fd_sc_hd__a21o_1 _11131_ (.A1(net859),
    .A2(net23),
    .B1(_02760_),
    .X(_02761_));
 sky130_fd_sc_hd__mux2_1 _11132_ (.A0(net576),
    .A1(_02761_),
    .S(net25),
    .X(_00140_));
 sky130_fd_sc_hd__a22o_1 _11133_ (.A1(net868),
    .A2(net50),
    .B1(net46),
    .B2(net822),
    .X(_02762_));
 sky130_fd_sc_hd__a21o_1 _11134_ (.A1(net855),
    .A2(net23),
    .B1(_02762_),
    .X(_02763_));
 sky130_fd_sc_hd__mux2_1 _11135_ (.A0(net571),
    .A1(_02763_),
    .S(net25),
    .X(_00141_));
 sky130_fd_sc_hd__a22o_1 _11136_ (.A1(net963),
    .A2(net50),
    .B1(net46),
    .B2(net838),
    .X(_02764_));
 sky130_fd_sc_hd__a21o_1 _11137_ (.A1(net842),
    .A2(net23),
    .B1(_02764_),
    .X(_02765_));
 sky130_fd_sc_hd__mux2_1 _11138_ (.A0(net566),
    .A1(_02765_),
    .S(net25),
    .X(_00142_));
 sky130_fd_sc_hd__a22o_1 _11139_ (.A1(\in_data[4] ),
    .A2(net50),
    .B1(net45),
    .B2(net811),
    .X(_02766_));
 sky130_fd_sc_hd__a21o_1 _11140_ (.A1(net823),
    .A2(net23),
    .B1(_02766_),
    .X(_02767_));
 sky130_fd_sc_hd__mux2_1 _11141_ (.A0(net561),
    .A1(_02767_),
    .S(net25),
    .X(_00143_));
 sky130_fd_sc_hd__a22o_1 _11142_ (.A1(net901),
    .A2(net50),
    .B1(net45),
    .B2(net832),
    .X(_02768_));
 sky130_fd_sc_hd__a21o_1 _11143_ (.A1(net785),
    .A2(net23),
    .B1(_02768_),
    .X(_02769_));
 sky130_fd_sc_hd__mux2_1 _11144_ (.A0(net557),
    .A1(_02769_),
    .S(net25),
    .X(_00144_));
 sky130_fd_sc_hd__a22o_1 _11145_ (.A1(net877),
    .A2(_02753_),
    .B1(net45),
    .B2(net825),
    .X(_02770_));
 sky130_fd_sc_hd__a21o_1 _11146_ (.A1(net850),
    .A2(net23),
    .B1(_02770_),
    .X(_02771_));
 sky130_fd_sc_hd__mux2_1 _11147_ (.A0(net553),
    .A1(_02771_),
    .S(net24),
    .X(_00145_));
 sky130_fd_sc_hd__a22o_1 _11148_ (.A1(net906),
    .A2(net50),
    .B1(net46),
    .B2(net795),
    .X(_02772_));
 sky130_fd_sc_hd__a21o_1 _11149_ (.A1(net828),
    .A2(net23),
    .B1(_02772_),
    .X(_02773_));
 sky130_fd_sc_hd__mux2_1 _11150_ (.A0(net549),
    .A1(_02773_),
    .S(net24),
    .X(_00146_));
 sky130_fd_sc_hd__a22o_1 _11151_ (.A1(net894),
    .A2(net50),
    .B1(net45),
    .B2(\in_data[72] ),
    .X(_02774_));
 sky130_fd_sc_hd__a21o_1 _11152_ (.A1(net829),
    .A2(net23),
    .B1(_02774_),
    .X(_02775_));
 sky130_fd_sc_hd__mux2_1 _11153_ (.A0(net544),
    .A1(_02775_),
    .S(net24),
    .X(_00147_));
 sky130_fd_sc_hd__a22o_1 _11154_ (.A1(net960),
    .A2(net50),
    .B1(net45),
    .B2(\in_data[73] ),
    .X(_02776_));
 sky130_fd_sc_hd__a21o_1 _11155_ (.A1(net845),
    .A2(net23),
    .B1(_02776_),
    .X(_02777_));
 sky130_fd_sc_hd__mux2_1 _11156_ (.A0(net540),
    .A1(_02777_),
    .S(net25),
    .X(_00148_));
 sky130_fd_sc_hd__a22o_1 _11157_ (.A1(net924),
    .A2(net50),
    .B1(net45),
    .B2(\in_data[74] ),
    .X(_02778_));
 sky130_fd_sc_hd__a21o_1 _11158_ (.A1(net856),
    .A2(net23),
    .B1(_02778_),
    .X(_02779_));
 sky130_fd_sc_hd__mux2_1 _11159_ (.A0(net535),
    .A1(_02779_),
    .S(net24),
    .X(_00149_));
 sky130_fd_sc_hd__a22o_1 _11160_ (.A1(net964),
    .A2(net50),
    .B1(net45),
    .B2(\in_data[75] ),
    .X(_02780_));
 sky130_fd_sc_hd__a21o_1 _11161_ (.A1(net857),
    .A2(net23),
    .B1(_02780_),
    .X(_02781_));
 sky130_fd_sc_hd__mux2_1 _11162_ (.A0(net530),
    .A1(_02781_),
    .S(net24),
    .X(_00150_));
 sky130_fd_sc_hd__a22o_1 _11163_ (.A1(net896),
    .A2(net50),
    .B1(net45),
    .B2(\in_data[76] ),
    .X(_02782_));
 sky130_fd_sc_hd__a21o_1 _11164_ (.A1(net769),
    .A2(net23),
    .B1(_02782_),
    .X(_02783_));
 sky130_fd_sc_hd__mux2_1 _11165_ (.A0(net525),
    .A1(_02783_),
    .S(net24),
    .X(_00151_));
 sky130_fd_sc_hd__a22o_1 _11166_ (.A1(net900),
    .A2(net50),
    .B1(net47),
    .B2(net958),
    .X(_02784_));
 sky130_fd_sc_hd__a21o_1 _11167_ (.A1(net816),
    .A2(net23),
    .B1(_02784_),
    .X(_02785_));
 sky130_fd_sc_hd__mux2_1 _11168_ (.A0(net520),
    .A1(_02785_),
    .S(net24),
    .X(_00152_));
 sky130_fd_sc_hd__a22o_1 _11169_ (.A1(net912),
    .A2(net51),
    .B1(net49),
    .B2(\in_data[78] ),
    .X(_02786_));
 sky130_fd_sc_hd__a21o_1 _11170_ (.A1(net844),
    .A2(net22),
    .B1(_02786_),
    .X(_02787_));
 sky130_fd_sc_hd__mux2_1 _11171_ (.A0(net515),
    .A1(_02787_),
    .S(net24),
    .X(_00153_));
 sky130_fd_sc_hd__a22o_1 _11172_ (.A1(net911),
    .A2(net50),
    .B1(net47),
    .B2(\in_data[79] ),
    .X(_02788_));
 sky130_fd_sc_hd__a21o_1 _11173_ (.A1(net799),
    .A2(net23),
    .B1(_02788_),
    .X(_02789_));
 sky130_fd_sc_hd__mux2_1 _11174_ (.A0(net511),
    .A1(_02789_),
    .S(net24),
    .X(_00154_));
 sky130_fd_sc_hd__a22o_1 _11175_ (.A1(net928),
    .A2(net51),
    .B1(net47),
    .B2(\in_data[80] ),
    .X(_02790_));
 sky130_fd_sc_hd__a21o_1 _11176_ (.A1(net800),
    .A2(net22),
    .B1(_02790_),
    .X(_02791_));
 sky130_fd_sc_hd__mux2_1 _11177_ (.A0(net507),
    .A1(_02791_),
    .S(net24),
    .X(_00155_));
 sky130_fd_sc_hd__a22o_1 _11178_ (.A1(net925),
    .A2(net51),
    .B1(net47),
    .B2(\in_data[81] ),
    .X(_02792_));
 sky130_fd_sc_hd__a21o_1 _11179_ (.A1(net830),
    .A2(net22),
    .B1(_02792_),
    .X(_02793_));
 sky130_fd_sc_hd__mux2_1 _11180_ (.A0(net503),
    .A1(_02793_),
    .S(net24),
    .X(_00156_));
 sky130_fd_sc_hd__a22o_1 _11181_ (.A1(net941),
    .A2(net51),
    .B1(net47),
    .B2(\in_data[82] ),
    .X(_02794_));
 sky130_fd_sc_hd__a21o_1 _11182_ (.A1(net808),
    .A2(net22),
    .B1(_02794_),
    .X(_02795_));
 sky130_fd_sc_hd__mux2_1 _11183_ (.A0(net498),
    .A1(_02795_),
    .S(net24),
    .X(_00157_));
 sky130_fd_sc_hd__a22o_1 _11184_ (.A1(net947),
    .A2(net51),
    .B1(net47),
    .B2(\in_data[83] ),
    .X(_02796_));
 sky130_fd_sc_hd__a21o_1 _11185_ (.A1(net788),
    .A2(net22),
    .B1(_02796_),
    .X(_02797_));
 sky130_fd_sc_hd__mux2_1 _11186_ (.A0(net494),
    .A1(_02797_),
    .S(net24),
    .X(_00158_));
 sky130_fd_sc_hd__a22o_1 _11187_ (.A1(net913),
    .A2(net51),
    .B1(net47),
    .B2(\in_data[84] ),
    .X(_02798_));
 sky130_fd_sc_hd__a21o_1 _11188_ (.A1(net812),
    .A2(net22),
    .B1(_02798_),
    .X(_02799_));
 sky130_fd_sc_hd__mux2_1 _11189_ (.A0(net490),
    .A1(_02799_),
    .S(net24),
    .X(_00159_));
 sky130_fd_sc_hd__a22o_1 _11190_ (.A1(net948),
    .A2(net51),
    .B1(net47),
    .B2(net926),
    .X(_02800_));
 sky130_fd_sc_hd__a21o_1 _11191_ (.A1(net777),
    .A2(net22),
    .B1(_02800_),
    .X(_02801_));
 sky130_fd_sc_hd__mux2_1 _11192_ (.A0(net486),
    .A1(_02801_),
    .S(net24),
    .X(_00160_));
 sky130_fd_sc_hd__a22o_1 _11193_ (.A1(net943),
    .A2(net51),
    .B1(net47),
    .B2(\in_data[86] ),
    .X(_02802_));
 sky130_fd_sc_hd__a21o_1 _11194_ (.A1(net762),
    .A2(net22),
    .B1(_02802_),
    .X(_02803_));
 sky130_fd_sc_hd__mux2_1 _11195_ (.A0(net482),
    .A1(_02803_),
    .S(net24),
    .X(_00161_));
 sky130_fd_sc_hd__a22o_1 _11196_ (.A1(net937),
    .A2(net51),
    .B1(net48),
    .B2(net879),
    .X(_02804_));
 sky130_fd_sc_hd__a21o_1 _11197_ (.A1(net810),
    .A2(net22),
    .B1(_02804_),
    .X(_02805_));
 sky130_fd_sc_hd__mux2_1 _11198_ (.A0(net478),
    .A1(_02805_),
    .S(net26),
    .X(_00162_));
 sky130_fd_sc_hd__a22o_1 _11199_ (.A1(net942),
    .A2(net51),
    .B1(net48),
    .B2(\in_data[88] ),
    .X(_02806_));
 sky130_fd_sc_hd__a21o_1 _11200_ (.A1(net776),
    .A2(net22),
    .B1(_02806_),
    .X(_02807_));
 sky130_fd_sc_hd__mux2_1 _11201_ (.A0(net474),
    .A1(_02807_),
    .S(net26),
    .X(_00163_));
 sky130_fd_sc_hd__a22o_1 _11202_ (.A1(net939),
    .A2(net51),
    .B1(net48),
    .B2(net874),
    .X(_02808_));
 sky130_fd_sc_hd__a21o_1 _11203_ (.A1(net853),
    .A2(net22),
    .B1(_02808_),
    .X(_02809_));
 sky130_fd_sc_hd__mux2_1 _11204_ (.A0(net470),
    .A1(_02809_),
    .S(net26),
    .X(_00164_));
 sky130_fd_sc_hd__a22o_1 _11205_ (.A1(net765),
    .A2(net51),
    .B1(net48),
    .B2(\in_data[90] ),
    .X(_02810_));
 sky130_fd_sc_hd__a21o_1 _11206_ (.A1(net824),
    .A2(net22),
    .B1(_02810_),
    .X(_02811_));
 sky130_fd_sc_hd__mux2_1 _11207_ (.A0(net466),
    .A1(_02811_),
    .S(net26),
    .X(_00165_));
 sky130_fd_sc_hd__a22o_1 _11208_ (.A1(net866),
    .A2(net51),
    .B1(net48),
    .B2(\in_data[91] ),
    .X(_02812_));
 sky130_fd_sc_hd__a21o_1 _11209_ (.A1(net807),
    .A2(net22),
    .B1(_02812_),
    .X(_02813_));
 sky130_fd_sc_hd__mux2_1 _11210_ (.A0(net463),
    .A1(_02813_),
    .S(net26),
    .X(_00166_));
 sky130_fd_sc_hd__a22o_1 _11211_ (.A1(net860),
    .A2(_02753_),
    .B1(net48),
    .B2(\in_data[92] ),
    .X(_02814_));
 sky130_fd_sc_hd__a21o_1 _11212_ (.A1(net827),
    .A2(net22),
    .B1(_02814_),
    .X(_02815_));
 sky130_fd_sc_hd__mux2_1 _11213_ (.A0(net460),
    .A1(_02815_),
    .S(net26),
    .X(_00167_));
 sky130_fd_sc_hd__a22o_1 _11214_ (.A1(net821),
    .A2(net51),
    .B1(net48),
    .B2(\in_data[93] ),
    .X(_02816_));
 sky130_fd_sc_hd__a21o_1 _11215_ (.A1(net826),
    .A2(_02757_),
    .B1(_02816_),
    .X(_02817_));
 sky130_fd_sc_hd__mux2_1 _11216_ (.A0(net459),
    .A1(_02817_),
    .S(net26),
    .X(_00168_));
 sky130_fd_sc_hd__a22o_1 _11217_ (.A1(net766),
    .A2(net51),
    .B1(net48),
    .B2(\in_data[94] ),
    .X(_02818_));
 sky130_fd_sc_hd__a21o_1 _11218_ (.A1(net847),
    .A2(net22),
    .B1(_02818_),
    .X(_02819_));
 sky130_fd_sc_hd__mux2_1 _11219_ (.A0(net457),
    .A1(_02819_),
    .S(net26),
    .X(_00169_));
 sky130_fd_sc_hd__a22o_1 _11220_ (.A1(net794),
    .A2(net51),
    .B1(net48),
    .B2(\in_data[95] ),
    .X(_02820_));
 sky130_fd_sc_hd__a21o_1 _11221_ (.A1(net848),
    .A2(net22),
    .B1(_02820_),
    .X(_02821_));
 sky130_fd_sc_hd__mux2_1 _11222_ (.A0(net959),
    .A1(_02821_),
    .S(net26),
    .X(_00170_));
 sky130_fd_sc_hd__or2_4 _11223_ (.A(net604),
    .B(net610),
    .X(_02822_));
 sky130_fd_sc_hd__nor2_4 _11224_ (.A(net591),
    .B(_02822_),
    .Y(_02823_));
 sky130_fd_sc_hd__a22o_1 _11225_ (.A1(net598),
    .A2(t2y[0]),
    .B1(t0y[0]),
    .B2(net607),
    .X(_02824_));
 sky130_fd_sc_hd__a221o_2 _11226_ (.A1(net587),
    .A2(t1x[0]),
    .B1(v2z[0]),
    .B2(net601),
    .C1(_02824_),
    .X(_02825_));
 sky130_fd_sc_hd__a31o_1 _11227_ (.A1(net59),
    .A2(v0z[0]),
    .A3(net19),
    .B1(_02825_),
    .X(_02826_));
 sky130_fd_sc_hd__mux2_1 _11228_ (.A0(net450),
    .A1(_02826_),
    .S(net25),
    .X(_00171_));
 sky130_fd_sc_hd__a22o_1 _11229_ (.A1(net598),
    .A2(t2y[1]),
    .B1(t0y[1]),
    .B2(net607),
    .X(_02827_));
 sky130_fd_sc_hd__a221o_2 _11230_ (.A1(net587),
    .A2(t1x[1]),
    .B1(v2z[1]),
    .B2(net601),
    .C1(_02827_),
    .X(_02828_));
 sky130_fd_sc_hd__a31o_1 _11231_ (.A1(net59),
    .A2(v0z[1]),
    .A3(net19),
    .B1(_02828_),
    .X(_02829_));
 sky130_fd_sc_hd__mux2_1 _11232_ (.A0(net445),
    .A1(_02829_),
    .S(net25),
    .X(_00172_));
 sky130_fd_sc_hd__a22o_1 _11233_ (.A1(net598),
    .A2(t2y[2]),
    .B1(t0y[2]),
    .B2(net607),
    .X(_02830_));
 sky130_fd_sc_hd__a221o_2 _11234_ (.A1(net587),
    .A2(t1x[2]),
    .B1(v2z[2]),
    .B2(net601),
    .C1(_02830_),
    .X(_02831_));
 sky130_fd_sc_hd__a31o_1 _11235_ (.A1(net59),
    .A2(v0z[2]),
    .A3(net19),
    .B1(_02831_),
    .X(_02832_));
 sky130_fd_sc_hd__mux2_1 _11236_ (.A0(net440),
    .A1(_02832_),
    .S(net25),
    .X(_00173_));
 sky130_fd_sc_hd__a22o_1 _11237_ (.A1(net598),
    .A2(t2y[3]),
    .B1(t0y[3]),
    .B2(net607),
    .X(_02833_));
 sky130_fd_sc_hd__a221o_2 _11238_ (.A1(net587),
    .A2(t1x[3]),
    .B1(v2z[3]),
    .B2(net606),
    .C1(_02833_),
    .X(_02834_));
 sky130_fd_sc_hd__a31o_1 _11239_ (.A1(net59),
    .A2(v0z[3]),
    .A3(net19),
    .B1(_02834_),
    .X(_02835_));
 sky130_fd_sc_hd__mux2_1 _11240_ (.A0(net436),
    .A1(_02835_),
    .S(net25),
    .X(_00174_));
 sky130_fd_sc_hd__a22o_1 _11241_ (.A1(net598),
    .A2(t2y[4]),
    .B1(t0y[4]),
    .B2(net607),
    .X(_02836_));
 sky130_fd_sc_hd__a221o_2 _11242_ (.A1(net587),
    .A2(t1x[4]),
    .B1(v2z[4]),
    .B2(net601),
    .C1(_02836_),
    .X(_02837_));
 sky130_fd_sc_hd__a31o_1 _11243_ (.A1(net59),
    .A2(v0z[4]),
    .A3(net19),
    .B1(_02837_),
    .X(_02838_));
 sky130_fd_sc_hd__mux2_1 _11244_ (.A0(net431),
    .A1(_02838_),
    .S(net25),
    .X(_00175_));
 sky130_fd_sc_hd__a22o_1 _11245_ (.A1(net598),
    .A2(t2y[5]),
    .B1(t0y[5]),
    .B2(net607),
    .X(_02839_));
 sky130_fd_sc_hd__a221o_2 _11246_ (.A1(net592),
    .A2(t1x[5]),
    .B1(v2z[5]),
    .B2(net601),
    .C1(_02839_),
    .X(_02840_));
 sky130_fd_sc_hd__a31o_1 _11247_ (.A1(net59),
    .A2(v0z[5]),
    .A3(net19),
    .B1(_02840_),
    .X(_02841_));
 sky130_fd_sc_hd__mux2_1 _11248_ (.A0(net426),
    .A1(_02841_),
    .S(net25),
    .X(_00176_));
 sky130_fd_sc_hd__a22o_1 _11249_ (.A1(net598),
    .A2(t2y[6]),
    .B1(t0y[6]),
    .B2(net607),
    .X(_02842_));
 sky130_fd_sc_hd__a221o_2 _11250_ (.A1(net588),
    .A2(t1x[6]),
    .B1(v2z[6]),
    .B2(net601),
    .C1(_02842_),
    .X(_02843_));
 sky130_fd_sc_hd__a31o_1 _11251_ (.A1(net59),
    .A2(v0z[6]),
    .A3(net19),
    .B1(_02843_),
    .X(_02844_));
 sky130_fd_sc_hd__mux2_1 _11252_ (.A0(net421),
    .A1(_02844_),
    .S(net25),
    .X(_00177_));
 sky130_fd_sc_hd__a22o_1 _11253_ (.A1(net598),
    .A2(t2y[7]),
    .B1(t0y[7]),
    .B2(net607),
    .X(_02845_));
 sky130_fd_sc_hd__a221o_2 _11254_ (.A1(net588),
    .A2(t1x[7]),
    .B1(v2z[7]),
    .B2(net606),
    .C1(_02845_),
    .X(_02846_));
 sky130_fd_sc_hd__a31o_1 _11255_ (.A1(net59),
    .A2(v0z[7]),
    .A3(net19),
    .B1(_02846_),
    .X(_02847_));
 sky130_fd_sc_hd__mux2_1 _11256_ (.A0(net417),
    .A1(_02847_),
    .S(net26),
    .X(_00178_));
 sky130_fd_sc_hd__a22o_1 _11257_ (.A1(net593),
    .A2(t2y[8]),
    .B1(t0y[8]),
    .B2(net608),
    .X(_02848_));
 sky130_fd_sc_hd__a221o_2 _11258_ (.A1(net588),
    .A2(t1x[8]),
    .B1(v2z[8]),
    .B2(net602),
    .C1(_02848_),
    .X(_02849_));
 sky130_fd_sc_hd__a31o_1 _11259_ (.A1(net59),
    .A2(v0z[8]),
    .A3(net19),
    .B1(_02849_),
    .X(_02850_));
 sky130_fd_sc_hd__mux2_1 _11260_ (.A0(net413),
    .A1(_02850_),
    .S(net25),
    .X(_00179_));
 sky130_fd_sc_hd__a22o_1 _11261_ (.A1(net593),
    .A2(t2y[9]),
    .B1(t0y[9]),
    .B2(net608),
    .X(_02851_));
 sky130_fd_sc_hd__a221o_2 _11262_ (.A1(net588),
    .A2(t1x[9]),
    .B1(v2z[9]),
    .B2(net602),
    .C1(_02851_),
    .X(_02852_));
 sky130_fd_sc_hd__a31o_1 _11263_ (.A1(net59),
    .A2(v0z[9]),
    .A3(net19),
    .B1(_02852_),
    .X(_02853_));
 sky130_fd_sc_hd__mux2_1 _11264_ (.A0(net408),
    .A1(_02853_),
    .S(net26),
    .X(_00180_));
 sky130_fd_sc_hd__a22o_1 _11265_ (.A1(net593),
    .A2(t2y[10]),
    .B1(t0y[10]),
    .B2(net608),
    .X(_02854_));
 sky130_fd_sc_hd__a221o_2 _11266_ (.A1(net588),
    .A2(t1x[10]),
    .B1(v2z[10]),
    .B2(net602),
    .C1(_02854_),
    .X(_02855_));
 sky130_fd_sc_hd__a31o_1 _11267_ (.A1(net58),
    .A2(v0z[10]),
    .A3(net17),
    .B1(_02855_),
    .X(_02856_));
 sky130_fd_sc_hd__mux2_1 _11268_ (.A0(net404),
    .A1(_02856_),
    .S(net26),
    .X(_00181_));
 sky130_fd_sc_hd__a22o_1 _11269_ (.A1(net593),
    .A2(t2y[11]),
    .B1(t0y[11]),
    .B2(net608),
    .X(_02857_));
 sky130_fd_sc_hd__a221o_2 _11270_ (.A1(net588),
    .A2(t1x[11]),
    .B1(v2z[11]),
    .B2(net602),
    .C1(_02857_),
    .X(_02858_));
 sky130_fd_sc_hd__a31o_1 _11271_ (.A1(net58),
    .A2(v0z[11]),
    .A3(net17),
    .B1(_02858_),
    .X(_02859_));
 sky130_fd_sc_hd__mux2_1 _11272_ (.A0(net400),
    .A1(_02859_),
    .S(net27),
    .X(_00182_));
 sky130_fd_sc_hd__a22o_1 _11273_ (.A1(net593),
    .A2(t2y[12]),
    .B1(t0y[12]),
    .B2(net608),
    .X(_02860_));
 sky130_fd_sc_hd__a221o_2 _11274_ (.A1(net589),
    .A2(t1x[12]),
    .B1(v2z[12]),
    .B2(net602),
    .C1(_02860_),
    .X(_02861_));
 sky130_fd_sc_hd__a31o_1 _11275_ (.A1(net58),
    .A2(v0z[12]),
    .A3(net17),
    .B1(_02861_),
    .X(_02862_));
 sky130_fd_sc_hd__mux2_1 _11276_ (.A0(net396),
    .A1(_02862_),
    .S(net27),
    .X(_00183_));
 sky130_fd_sc_hd__a22o_1 _11277_ (.A1(net593),
    .A2(t2y[13]),
    .B1(t0y[13]),
    .B2(net608),
    .X(_02863_));
 sky130_fd_sc_hd__a221o_2 _11278_ (.A1(net589),
    .A2(t1x[13]),
    .B1(v2z[13]),
    .B2(net602),
    .C1(_02863_),
    .X(_02864_));
 sky130_fd_sc_hd__a31o_1 _11279_ (.A1(net58),
    .A2(v0z[13]),
    .A3(net17),
    .B1(_02864_),
    .X(_02865_));
 sky130_fd_sc_hd__mux2_1 _11280_ (.A0(net390),
    .A1(_02865_),
    .S(net27),
    .X(_00184_));
 sky130_fd_sc_hd__a22o_1 _11281_ (.A1(net593),
    .A2(t2y[14]),
    .B1(t0y[14]),
    .B2(net609),
    .X(_02866_));
 sky130_fd_sc_hd__a221o_2 _11282_ (.A1(net588),
    .A2(t1x[14]),
    .B1(v2z[14]),
    .B2(net602),
    .C1(_02866_),
    .X(_02867_));
 sky130_fd_sc_hd__a31o_1 _11283_ (.A1(net58),
    .A2(v0z[14]),
    .A3(net17),
    .B1(_02867_),
    .X(_02868_));
 sky130_fd_sc_hd__mux2_1 _11284_ (.A0(net386),
    .A1(_02868_),
    .S(net26),
    .X(_00185_));
 sky130_fd_sc_hd__a22o_1 _11285_ (.A1(net593),
    .A2(t2y[15]),
    .B1(t0y[15]),
    .B2(net608),
    .X(_02869_));
 sky130_fd_sc_hd__a221o_2 _11286_ (.A1(net589),
    .A2(t1x[15]),
    .B1(v2z[15]),
    .B2(net603),
    .C1(_02869_),
    .X(_02870_));
 sky130_fd_sc_hd__a31o_1 _11287_ (.A1(net58),
    .A2(v0z[15]),
    .A3(net17),
    .B1(_02870_),
    .X(_02871_));
 sky130_fd_sc_hd__mux2_1 _11288_ (.A0(net381),
    .A1(_02871_),
    .S(net27),
    .X(_00186_));
 sky130_fd_sc_hd__a22o_1 _11289_ (.A1(net593),
    .A2(t2y[16]),
    .B1(t0y[16]),
    .B2(net609),
    .X(_02872_));
 sky130_fd_sc_hd__a221o_2 _11290_ (.A1(net589),
    .A2(t1x[16]),
    .B1(v2z[16]),
    .B2(net603),
    .C1(_02872_),
    .X(_02873_));
 sky130_fd_sc_hd__a31o_1 _11291_ (.A1(net58),
    .A2(v0z[16]),
    .A3(net17),
    .B1(_02873_),
    .X(_02874_));
 sky130_fd_sc_hd__mux2_1 _11292_ (.A0(net375),
    .A1(_02874_),
    .S(net27),
    .X(_00187_));
 sky130_fd_sc_hd__a22o_1 _11293_ (.A1(net593),
    .A2(t2y[17]),
    .B1(t0y[17]),
    .B2(net608),
    .X(_02875_));
 sky130_fd_sc_hd__a221o_2 _11294_ (.A1(net589),
    .A2(t1x[17]),
    .B1(v2z[17]),
    .B2(net603),
    .C1(_02875_),
    .X(_02876_));
 sky130_fd_sc_hd__a31o_1 _11295_ (.A1(net58),
    .A2(v0z[17]),
    .A3(net18),
    .B1(_02876_),
    .X(_02877_));
 sky130_fd_sc_hd__mux2_1 _11296_ (.A0(net371),
    .A1(_02877_),
    .S(net27),
    .X(_00188_));
 sky130_fd_sc_hd__a22o_1 _11297_ (.A1(net593),
    .A2(t2y[18]),
    .B1(t0y[18]),
    .B2(net609),
    .X(_02878_));
 sky130_fd_sc_hd__a221o_2 _11298_ (.A1(net591),
    .A2(t1x[18]),
    .B1(v2z[18]),
    .B2(net603),
    .C1(_02878_),
    .X(_02879_));
 sky130_fd_sc_hd__a31o_1 _11299_ (.A1(net58),
    .A2(v0z[18]),
    .A3(net18),
    .B1(_02879_),
    .X(_02880_));
 sky130_fd_sc_hd__mux2_1 _11300_ (.A0(net631),
    .A1(_02880_),
    .S(net27),
    .X(_00189_));
 sky130_fd_sc_hd__a22o_1 _11301_ (.A1(net593),
    .A2(t2y[19]),
    .B1(t0y[19]),
    .B2(net609),
    .X(_02881_));
 sky130_fd_sc_hd__a221o_2 _11302_ (.A1(net591),
    .A2(t1x[19]),
    .B1(v2z[19]),
    .B2(net603),
    .C1(_02881_),
    .X(_02882_));
 sky130_fd_sc_hd__a31o_1 _11303_ (.A1(net58),
    .A2(v0z[19]),
    .A3(net18),
    .B1(_02882_),
    .X(_02883_));
 sky130_fd_sc_hd__mux2_1 _11304_ (.A0(net365),
    .A1(_02883_),
    .S(net27),
    .X(_00190_));
 sky130_fd_sc_hd__a22o_1 _11305_ (.A1(net593),
    .A2(t2y[20]),
    .B1(t0y[20]),
    .B2(net610),
    .X(_02884_));
 sky130_fd_sc_hd__a221o_2 _11306_ (.A1(net591),
    .A2(t1x[20]),
    .B1(v2z[20]),
    .B2(net604),
    .C1(_02884_),
    .X(_02885_));
 sky130_fd_sc_hd__a31o_1 _11307_ (.A1(net58),
    .A2(v0z[20]),
    .A3(net17),
    .B1(_02885_),
    .X(_02886_));
 sky130_fd_sc_hd__mux2_1 _11308_ (.A0(net364),
    .A1(_02886_),
    .S(net27),
    .X(_00191_));
 sky130_fd_sc_hd__a22o_1 _11309_ (.A1(net594),
    .A2(t2y[21]),
    .B1(t0y[21]),
    .B2(net610),
    .X(_02887_));
 sky130_fd_sc_hd__a221o_2 _11310_ (.A1(net591),
    .A2(t1x[21]),
    .B1(v2z[21]),
    .B2(net604),
    .C1(_02887_),
    .X(_02888_));
 sky130_fd_sc_hd__a31o_1 _11311_ (.A1(net58),
    .A2(v0z[21]),
    .A3(net17),
    .B1(_02888_),
    .X(_02889_));
 sky130_fd_sc_hd__mux2_1 _11312_ (.A0(net360),
    .A1(_02889_),
    .S(net27),
    .X(_00192_));
 sky130_fd_sc_hd__a22o_1 _11313_ (.A1(net594),
    .A2(t2y[22]),
    .B1(t0y[22]),
    .B2(net610),
    .X(_02890_));
 sky130_fd_sc_hd__a221o_2 _11314_ (.A1(net591),
    .A2(t1x[22]),
    .B1(v2z[22]),
    .B2(net604),
    .C1(_02890_),
    .X(_02891_));
 sky130_fd_sc_hd__a31o_1 _11315_ (.A1(net58),
    .A2(v0z[22]),
    .A3(net17),
    .B1(_02891_),
    .X(_02892_));
 sky130_fd_sc_hd__mux2_1 _11316_ (.A0(net355),
    .A1(_02892_),
    .S(net27),
    .X(_00193_));
 sky130_fd_sc_hd__a22o_1 _11317_ (.A1(net593),
    .A2(t2y[23]),
    .B1(t0y[23]),
    .B2(net610),
    .X(_02893_));
 sky130_fd_sc_hd__a221o_2 _11318_ (.A1(net591),
    .A2(t1x[23]),
    .B1(v2z[23]),
    .B2(net604),
    .C1(_02893_),
    .X(_02894_));
 sky130_fd_sc_hd__a31o_2 _11319_ (.A1(net59),
    .A2(v0z[23]),
    .A3(net18),
    .B1(_02894_),
    .X(_02895_));
 sky130_fd_sc_hd__mux2_1 _11320_ (.A0(net887),
    .A1(_02895_),
    .S(net27),
    .X(_00194_));
 sky130_fd_sc_hd__a22o_1 _11321_ (.A1(net593),
    .A2(t2y[24]),
    .B1(t0y[24]),
    .B2(net610),
    .X(_02896_));
 sky130_fd_sc_hd__a221o_2 _11322_ (.A1(net590),
    .A2(t1x[24]),
    .B1(v2z[24]),
    .B2(net604),
    .C1(_02896_),
    .X(_02897_));
 sky130_fd_sc_hd__a31o_2 _11323_ (.A1(net59),
    .A2(v0z[24]),
    .A3(net18),
    .B1(_02897_),
    .X(_02898_));
 sky130_fd_sc_hd__mux2_1 _11324_ (.A0(net345),
    .A1(_02898_),
    .S(net27),
    .X(_00195_));
 sky130_fd_sc_hd__a22o_1 _11325_ (.A1(net593),
    .A2(t2y[25]),
    .B1(t0y[25]),
    .B2(net611),
    .X(_02899_));
 sky130_fd_sc_hd__a221o_2 _11326_ (.A1(net590),
    .A2(t1x[25]),
    .B1(v2z[25]),
    .B2(net605),
    .C1(_02899_),
    .X(_02900_));
 sky130_fd_sc_hd__a31o_2 _11327_ (.A1(net58),
    .A2(v0z[25]),
    .A3(net18),
    .B1(_02900_),
    .X(_02901_));
 sky130_fd_sc_hd__mux2_1 _11328_ (.A0(net341),
    .A1(_02901_),
    .S(net27),
    .X(_00196_));
 sky130_fd_sc_hd__a22o_1 _11329_ (.A1(net594),
    .A2(t2y[26]),
    .B1(t0y[26]),
    .B2(net611),
    .X(_02902_));
 sky130_fd_sc_hd__a221o_2 _11330_ (.A1(net590),
    .A2(t1x[26]),
    .B1(v2z[26]),
    .B2(net604),
    .C1(_02902_),
    .X(_02903_));
 sky130_fd_sc_hd__a31o_2 _11331_ (.A1(net58),
    .A2(v0z[26]),
    .A3(net18),
    .B1(_02903_),
    .X(_02904_));
 sky130_fd_sc_hd__mux2_1 _11332_ (.A0(net339),
    .A1(_02904_),
    .S(net27),
    .X(_00197_));
 sky130_fd_sc_hd__a22o_1 _11333_ (.A1(net594),
    .A2(t2y[27]),
    .B1(t0y[27]),
    .B2(net610),
    .X(_02905_));
 sky130_fd_sc_hd__a221o_2 _11334_ (.A1(net590),
    .A2(t1x[27]),
    .B1(v2z[27]),
    .B2(net605),
    .C1(_02905_),
    .X(_02906_));
 sky130_fd_sc_hd__a31o_2 _11335_ (.A1(net61),
    .A2(v0z[27]),
    .A3(net20),
    .B1(_02906_),
    .X(_02907_));
 sky130_fd_sc_hd__mux2_1 _11336_ (.A0(net334),
    .A1(_02907_),
    .S(_02756_),
    .X(_00198_));
 sky130_fd_sc_hd__a22o_1 _11337_ (.A1(net594),
    .A2(t2y[28]),
    .B1(t0y[28]),
    .B2(net610),
    .X(_02908_));
 sky130_fd_sc_hd__a221o_2 _11338_ (.A1(net590),
    .A2(t1x[28]),
    .B1(v2z[28]),
    .B2(net605),
    .C1(_02908_),
    .X(_02909_));
 sky130_fd_sc_hd__a31o_2 _11339_ (.A1(net61),
    .A2(v0z[28]),
    .A3(net20),
    .B1(_02909_),
    .X(_02910_));
 sky130_fd_sc_hd__mux2_1 _11340_ (.A0(net331),
    .A1(_02910_),
    .S(_02756_),
    .X(_00199_));
 sky130_fd_sc_hd__a22o_1 _11341_ (.A1(net594),
    .A2(t2y[29]),
    .B1(t0y[29]),
    .B2(net610),
    .X(_02911_));
 sky130_fd_sc_hd__a221o_2 _11342_ (.A1(net590),
    .A2(t1x[29]),
    .B1(v2z[29]),
    .B2(net605),
    .C1(_02911_),
    .X(_02912_));
 sky130_fd_sc_hd__a31o_2 _11343_ (.A1(net61),
    .A2(v0z[29]),
    .A3(net20),
    .B1(_02912_),
    .X(_02913_));
 sky130_fd_sc_hd__mux2_1 _11344_ (.A0(net329),
    .A1(_02913_),
    .S(_02756_),
    .X(_00200_));
 sky130_fd_sc_hd__a22o_1 _11345_ (.A1(net594),
    .A2(t2y[30]),
    .B1(t0y[30]),
    .B2(net611),
    .X(_02914_));
 sky130_fd_sc_hd__a221o_2 _11346_ (.A1(net590),
    .A2(t1x[30]),
    .B1(v2z[30]),
    .B2(net605),
    .C1(_02914_),
    .X(_02915_));
 sky130_fd_sc_hd__a31o_2 _11347_ (.A1(net61),
    .A2(v0z[30]),
    .A3(net20),
    .B1(_02915_),
    .X(_02916_));
 sky130_fd_sc_hd__mux2_1 _11348_ (.A0(net327),
    .A1(_02916_),
    .S(_02756_),
    .X(_00201_));
 sky130_fd_sc_hd__a22o_1 _11349_ (.A1(net594),
    .A2(t2y[31]),
    .B1(t0y[31]),
    .B2(net611),
    .X(_02917_));
 sky130_fd_sc_hd__a221o_4 _11350_ (.A1(net590),
    .A2(t1x[31]),
    .B1(v2z[31]),
    .B2(net605),
    .C1(_02917_),
    .X(_02918_));
 sky130_fd_sc_hd__a31o_1 _11351_ (.A1(net58),
    .A2(v0z[31]),
    .A3(net17),
    .B1(_02918_),
    .X(_02919_));
 sky130_fd_sc_hd__mux2_1 _11352_ (.A0(net965),
    .A1(_02919_),
    .S(net27),
    .X(_00202_));
 sky130_fd_sc_hd__o31ai_2 _11353_ (.A1(net587),
    .A2(net601),
    .A3(net46),
    .B1(net646),
    .Y(_02920_));
 sky130_fd_sc_hd__a22o_1 _11354_ (.A1(net585),
    .A2(\in_data[0] ),
    .B1(net46),
    .B2(net806),
    .X(_02921_));
 sky130_fd_sc_hd__a21o_1 _11355_ (.A1(net846),
    .A2(net29),
    .B1(_02921_),
    .X(_02922_));
 sky130_fd_sc_hd__mux2_1 _11356_ (.A0(_02922_),
    .A1(net322),
    .S(net11),
    .X(_00203_));
 sky130_fd_sc_hd__a22o_1 _11357_ (.A1(net585),
    .A2(net870),
    .B1(net46),
    .B2(net859),
    .X(_02923_));
 sky130_fd_sc_hd__a21o_1 _11358_ (.A1(net843),
    .A2(net29),
    .B1(_02923_),
    .X(_02924_));
 sky130_fd_sc_hd__mux2_1 _11359_ (.A0(_02924_),
    .A1(net318),
    .S(net11),
    .X(_00204_));
 sky130_fd_sc_hd__a22o_1 _11360_ (.A1(net587),
    .A2(net868),
    .B1(net46),
    .B2(net855),
    .X(_02925_));
 sky130_fd_sc_hd__a21o_1 _11361_ (.A1(net822),
    .A2(net29),
    .B1(_02925_),
    .X(_02926_));
 sky130_fd_sc_hd__mux2_1 _11362_ (.A0(_02926_),
    .A1(net313),
    .S(net11),
    .X(_00205_));
 sky130_fd_sc_hd__a22o_1 _11363_ (.A1(net585),
    .A2(net876),
    .B1(net46),
    .B2(net842),
    .X(_02927_));
 sky130_fd_sc_hd__a21o_1 _11364_ (.A1(net838),
    .A2(net29),
    .B1(_02927_),
    .X(_02928_));
 sky130_fd_sc_hd__mux2_1 _11365_ (.A0(_02928_),
    .A1(net309),
    .S(net11),
    .X(_00206_));
 sky130_fd_sc_hd__a22o_1 _11366_ (.A1(net585),
    .A2(\in_data[4] ),
    .B1(net45),
    .B2(net823),
    .X(_02929_));
 sky130_fd_sc_hd__a21o_1 _11367_ (.A1(net811),
    .A2(net29),
    .B1(_02929_),
    .X(_02930_));
 sky130_fd_sc_hd__mux2_1 _11368_ (.A0(_02930_),
    .A1(net304),
    .S(net11),
    .X(_00207_));
 sky130_fd_sc_hd__a22o_1 _11369_ (.A1(net585),
    .A2(net901),
    .B1(net45),
    .B2(net785),
    .X(_02931_));
 sky130_fd_sc_hd__a21o_1 _11370_ (.A1(net832),
    .A2(net29),
    .B1(_02931_),
    .X(_02932_));
 sky130_fd_sc_hd__mux2_1 _11371_ (.A0(_02932_),
    .A1(net299),
    .S(net11),
    .X(_00208_));
 sky130_fd_sc_hd__a22o_1 _11372_ (.A1(net585),
    .A2(net877),
    .B1(net45),
    .B2(net850),
    .X(_02933_));
 sky130_fd_sc_hd__a21o_1 _11373_ (.A1(net825),
    .A2(net29),
    .B1(_02933_),
    .X(_02934_));
 sky130_fd_sc_hd__mux2_1 _11374_ (.A0(_02934_),
    .A1(net294),
    .S(net11),
    .X(_00209_));
 sky130_fd_sc_hd__a22o_1 _11375_ (.A1(net586),
    .A2(net906),
    .B1(net46),
    .B2(net828),
    .X(_02935_));
 sky130_fd_sc_hd__a21o_1 _11376_ (.A1(net795),
    .A2(net29),
    .B1(_02935_),
    .X(_02936_));
 sky130_fd_sc_hd__mux2_1 _11377_ (.A0(_02936_),
    .A1(net289),
    .S(net11),
    .X(_00210_));
 sky130_fd_sc_hd__a22o_1 _11378_ (.A1(net585),
    .A2(net894),
    .B1(net45),
    .B2(net829),
    .X(_02937_));
 sky130_fd_sc_hd__a21o_1 _11379_ (.A1(net944),
    .A2(net29),
    .B1(_02937_),
    .X(_02938_));
 sky130_fd_sc_hd__mux2_1 _11380_ (.A0(_02938_),
    .A1(net284),
    .S(net11),
    .X(_00211_));
 sky130_fd_sc_hd__a22o_1 _11381_ (.A1(net585),
    .A2(net888),
    .B1(net45),
    .B2(net845),
    .X(_02939_));
 sky130_fd_sc_hd__a21o_1 _11382_ (.A1(net954),
    .A2(net29),
    .B1(_02939_),
    .X(_02940_));
 sky130_fd_sc_hd__mux2_1 _11383_ (.A0(_02940_),
    .A1(net278),
    .S(net11),
    .X(_00212_));
 sky130_fd_sc_hd__a22o_1 _11384_ (.A1(net585),
    .A2(net924),
    .B1(net45),
    .B2(net856),
    .X(_02941_));
 sky130_fd_sc_hd__a21o_1 _11385_ (.A1(net962),
    .A2(net29),
    .B1(_02941_),
    .X(_02942_));
 sky130_fd_sc_hd__mux2_1 _11386_ (.A0(_02942_),
    .A1(net273),
    .S(net11),
    .X(_00213_));
 sky130_fd_sc_hd__a22o_1 _11387_ (.A1(net585),
    .A2(net890),
    .B1(net45),
    .B2(net857),
    .X(_02943_));
 sky130_fd_sc_hd__a21o_1 _11388_ (.A1(net907),
    .A2(net29),
    .B1(_02943_),
    .X(_02944_));
 sky130_fd_sc_hd__mux2_1 _11389_ (.A0(_02944_),
    .A1(net268),
    .S(net11),
    .X(_00214_));
 sky130_fd_sc_hd__a22o_1 _11390_ (.A1(net585),
    .A2(net896),
    .B1(net45),
    .B2(net769),
    .X(_02945_));
 sky130_fd_sc_hd__a21o_1 _11391_ (.A1(net949),
    .A2(net29),
    .B1(_02945_),
    .X(_02946_));
 sky130_fd_sc_hd__mux2_1 _11392_ (.A0(_02946_),
    .A1(net263),
    .S(net11),
    .X(_00215_));
 sky130_fd_sc_hd__a22o_1 _11393_ (.A1(net585),
    .A2(net900),
    .B1(net46),
    .B2(net816),
    .X(_02947_));
 sky130_fd_sc_hd__a21o_1 _11394_ (.A1(net938),
    .A2(net28),
    .B1(_02947_),
    .X(_02948_));
 sky130_fd_sc_hd__mux2_1 _11395_ (.A0(_02948_),
    .A1(net258),
    .S(net11),
    .X(_00216_));
 sky130_fd_sc_hd__a22o_1 _11396_ (.A1(net587),
    .A2(net912),
    .B1(net49),
    .B2(net844),
    .X(_02949_));
 sky130_fd_sc_hd__a21o_1 _11397_ (.A1(net950),
    .A2(net28),
    .B1(_02949_),
    .X(_02950_));
 sky130_fd_sc_hd__mux2_1 _11398_ (.A0(_02950_),
    .A1(net257),
    .S(net11),
    .X(_00217_));
 sky130_fd_sc_hd__a22o_1 _11399_ (.A1(net585),
    .A2(net911),
    .B1(net47),
    .B2(net799),
    .X(_02951_));
 sky130_fd_sc_hd__a21o_1 _11400_ (.A1(net915),
    .A2(net28),
    .B1(_02951_),
    .X(_02952_));
 sky130_fd_sc_hd__mux2_1 _11401_ (.A0(_02952_),
    .A1(net252),
    .S(net11),
    .X(_00218_));
 sky130_fd_sc_hd__a22o_1 _11402_ (.A1(net585),
    .A2(\in_data[16] ),
    .B1(net47),
    .B2(\in_data[48] ),
    .X(_02953_));
 sky130_fd_sc_hd__a21o_1 _11403_ (.A1(\in_data[80] ),
    .A2(net28),
    .B1(_02953_),
    .X(_02954_));
 sky130_fd_sc_hd__mux2_1 _11404_ (.A0(_02954_),
    .A1(net630),
    .S(net13),
    .X(_00219_));
 sky130_fd_sc_hd__a22o_1 _11405_ (.A1(net586),
    .A2(\in_data[17] ),
    .B1(net49),
    .B2(\in_data[49] ),
    .X(_02955_));
 sky130_fd_sc_hd__a21o_1 _11406_ (.A1(\in_data[81] ),
    .A2(net28),
    .B1(_02955_),
    .X(_02956_));
 sky130_fd_sc_hd__mux2_1 _11407_ (.A0(_02956_),
    .A1(net247),
    .S(net13),
    .X(_00220_));
 sky130_fd_sc_hd__a22o_1 _11408_ (.A1(net586),
    .A2(\in_data[18] ),
    .B1(net47),
    .B2(\in_data[50] ),
    .X(_02957_));
 sky130_fd_sc_hd__a21o_1 _11409_ (.A1(\in_data[82] ),
    .A2(net28),
    .B1(_02957_),
    .X(_02958_));
 sky130_fd_sc_hd__mux2_1 _11410_ (.A0(_02958_),
    .A1(net242),
    .S(net13),
    .X(_00221_));
 sky130_fd_sc_hd__a22o_1 _11411_ (.A1(net586),
    .A2(\in_data[19] ),
    .B1(net47),
    .B2(\in_data[51] ),
    .X(_02959_));
 sky130_fd_sc_hd__a21o_2 _11412_ (.A1(\in_data[83] ),
    .A2(net28),
    .B1(_02959_),
    .X(_02960_));
 sky130_fd_sc_hd__mux2_1 _11413_ (.A0(_02960_),
    .A1(net237),
    .S(net13),
    .X(_00222_));
 sky130_fd_sc_hd__a22o_1 _11414_ (.A1(net586),
    .A2(\in_data[20] ),
    .B1(net47),
    .B2(\in_data[52] ),
    .X(_02961_));
 sky130_fd_sc_hd__a21o_1 _11415_ (.A1(\in_data[84] ),
    .A2(net28),
    .B1(_02961_),
    .X(_02962_));
 sky130_fd_sc_hd__mux2_1 _11416_ (.A0(_02962_),
    .A1(net232),
    .S(net13),
    .X(_00223_));
 sky130_fd_sc_hd__a22o_1 _11417_ (.A1(net586),
    .A2(\in_data[21] ),
    .B1(net47),
    .B2(\in_data[53] ),
    .X(_02963_));
 sky130_fd_sc_hd__a21o_1 _11418_ (.A1(\in_data[85] ),
    .A2(net28),
    .B1(_02963_),
    .X(_02964_));
 sky130_fd_sc_hd__mux2_1 _11419_ (.A0(_02964_),
    .A1(net227),
    .S(net12),
    .X(_00224_));
 sky130_fd_sc_hd__a22o_1 _11420_ (.A1(net586),
    .A2(\in_data[22] ),
    .B1(net49),
    .B2(\in_data[54] ),
    .X(_02965_));
 sky130_fd_sc_hd__a21o_1 _11421_ (.A1(\in_data[86] ),
    .A2(net28),
    .B1(_02965_),
    .X(_02966_));
 sky130_fd_sc_hd__mux2_1 _11422_ (.A0(_02966_),
    .A1(net223),
    .S(net13),
    .X(_00225_));
 sky130_fd_sc_hd__a22o_1 _11423_ (.A1(net587),
    .A2(\in_data[23] ),
    .B1(net47),
    .B2(\in_data[55] ),
    .X(_02967_));
 sky130_fd_sc_hd__a21o_2 _11424_ (.A1(\in_data[87] ),
    .A2(net29),
    .B1(_02967_),
    .X(_02968_));
 sky130_fd_sc_hd__mux2_1 _11425_ (.A0(_02968_),
    .A1(net218),
    .S(net12),
    .X(_00226_));
 sky130_fd_sc_hd__a22o_1 _11426_ (.A1(net586),
    .A2(\in_data[24] ),
    .B1(net48),
    .B2(\in_data[56] ),
    .X(_02969_));
 sky130_fd_sc_hd__a21o_1 _11427_ (.A1(\in_data[88] ),
    .A2(net28),
    .B1(_02969_),
    .X(_02970_));
 sky130_fd_sc_hd__mux2_1 _11428_ (.A0(_02970_),
    .A1(net214),
    .S(net12),
    .X(_00227_));
 sky130_fd_sc_hd__a22o_1 _11429_ (.A1(net586),
    .A2(\in_data[25] ),
    .B1(net48),
    .B2(\in_data[57] ),
    .X(_02971_));
 sky130_fd_sc_hd__a21o_2 _11430_ (.A1(\in_data[89] ),
    .A2(net28),
    .B1(_02971_),
    .X(_02972_));
 sky130_fd_sc_hd__mux2_1 _11431_ (.A0(_02972_),
    .A1(net210),
    .S(net12),
    .X(_00228_));
 sky130_fd_sc_hd__a22o_1 _11432_ (.A1(net586),
    .A2(\in_data[26] ),
    .B1(net48),
    .B2(\in_data[58] ),
    .X(_02973_));
 sky130_fd_sc_hd__a21o_1 _11433_ (.A1(\in_data[90] ),
    .A2(net28),
    .B1(_02973_),
    .X(_02974_));
 sky130_fd_sc_hd__mux2_1 _11434_ (.A0(_02974_),
    .A1(net207),
    .S(net12),
    .X(_00229_));
 sky130_fd_sc_hd__a22o_1 _11435_ (.A1(net586),
    .A2(\in_data[27] ),
    .B1(net48),
    .B2(\in_data[59] ),
    .X(_02975_));
 sky130_fd_sc_hd__a21o_2 _11436_ (.A1(\in_data[91] ),
    .A2(net28),
    .B1(_02975_),
    .X(_02976_));
 sky130_fd_sc_hd__mux2_1 _11437_ (.A0(_02976_),
    .A1(net204),
    .S(net12),
    .X(_00230_));
 sky130_fd_sc_hd__a22o_1 _11438_ (.A1(net586),
    .A2(\in_data[28] ),
    .B1(net48),
    .B2(\in_data[60] ),
    .X(_02977_));
 sky130_fd_sc_hd__a21o_1 _11439_ (.A1(\in_data[92] ),
    .A2(net28),
    .B1(_02977_),
    .X(_02978_));
 sky130_fd_sc_hd__mux2_1 _11440_ (.A0(_02978_),
    .A1(net201),
    .S(net12),
    .X(_00231_));
 sky130_fd_sc_hd__a22o_1 _11441_ (.A1(net586),
    .A2(\in_data[29] ),
    .B1(net49),
    .B2(\in_data[61] ),
    .X(_02979_));
 sky130_fd_sc_hd__a21o_1 _11442_ (.A1(\in_data[93] ),
    .A2(net28),
    .B1(_02979_),
    .X(_02980_));
 sky130_fd_sc_hd__mux2_1 _11443_ (.A0(_02980_),
    .A1(net910),
    .S(net12),
    .X(_00232_));
 sky130_fd_sc_hd__a22o_1 _11444_ (.A1(net586),
    .A2(\in_data[30] ),
    .B1(net48),
    .B2(\in_data[62] ),
    .X(_02981_));
 sky130_fd_sc_hd__a21o_2 _11445_ (.A1(\in_data[94] ),
    .A2(net29),
    .B1(_02981_),
    .X(_02982_));
 sky130_fd_sc_hd__mux2_1 _11446_ (.A0(_02982_),
    .A1(net940),
    .S(net13),
    .X(_00233_));
 sky130_fd_sc_hd__a22o_1 _11447_ (.A1(net586),
    .A2(\in_data[31] ),
    .B1(net48),
    .B2(\in_data[63] ),
    .X(_02983_));
 sky130_fd_sc_hd__a21o_2 _11448_ (.A1(\in_data[95] ),
    .A2(_02755_),
    .B1(_02983_),
    .X(_02984_));
 sky130_fd_sc_hd__mux2_1 _11449_ (.A0(_02984_),
    .A1(net194),
    .S(net12),
    .X(_00234_));
 sky130_fd_sc_hd__a22o_1 _11450_ (.A1(net607),
    .A2(t1y[0]),
    .B1(t0x[0]),
    .B2(net601),
    .X(_02985_));
 sky130_fd_sc_hd__a221o_1 _11451_ (.A1(net592),
    .A2(t2x[0]),
    .B1(v1z[0]),
    .B2(net17),
    .C1(_02985_),
    .X(_02986_));
 sky130_fd_sc_hd__mux2_1 _11452_ (.A0(_02986_),
    .A1(net625),
    .S(net12),
    .X(_00235_));
 sky130_fd_sc_hd__a22o_1 _11453_ (.A1(\state[2] ),
    .A2(t1y[1]),
    .B1(t0x[1]),
    .B2(net601),
    .X(_02987_));
 sky130_fd_sc_hd__a221o_1 _11454_ (.A1(net587),
    .A2(t2x[1]),
    .B1(v1z[1]),
    .B2(net17),
    .C1(_02987_),
    .X(_02988_));
 sky130_fd_sc_hd__mux2_1 _11455_ (.A0(_02988_),
    .A1(net192),
    .S(net12),
    .X(_00236_));
 sky130_fd_sc_hd__a22o_1 _11456_ (.A1(net607),
    .A2(t1y[2]),
    .B1(t0x[2]),
    .B2(net601),
    .X(_02989_));
 sky130_fd_sc_hd__a221o_1 _11457_ (.A1(net587),
    .A2(t2x[2]),
    .B1(v1z[2]),
    .B2(net18),
    .C1(_02989_),
    .X(_02990_));
 sky130_fd_sc_hd__mux2_1 _11458_ (.A0(_02990_),
    .A1(net187),
    .S(net12),
    .X(_00237_));
 sky130_fd_sc_hd__a22o_1 _11459_ (.A1(net607),
    .A2(t1y[3]),
    .B1(t0x[3]),
    .B2(net606),
    .X(_02991_));
 sky130_fd_sc_hd__a221o_1 _11460_ (.A1(net587),
    .A2(t2x[3]),
    .B1(v1z[3]),
    .B2(net17),
    .C1(_02991_),
    .X(_02992_));
 sky130_fd_sc_hd__mux2_1 _11461_ (.A0(_02992_),
    .A1(net185),
    .S(net12),
    .X(_00238_));
 sky130_fd_sc_hd__a22o_1 _11462_ (.A1(net607),
    .A2(t1y[4]),
    .B1(t0x[4]),
    .B2(net601),
    .X(_02993_));
 sky130_fd_sc_hd__a221o_1 _11463_ (.A1(net587),
    .A2(t2x[4]),
    .B1(v1z[4]),
    .B2(net17),
    .C1(_02993_),
    .X(_02994_));
 sky130_fd_sc_hd__mux2_1 _11464_ (.A0(_02994_),
    .A1(net180),
    .S(net12),
    .X(_00239_));
 sky130_fd_sc_hd__a22o_1 _11465_ (.A1(net607),
    .A2(t1y[5]),
    .B1(t0x[5]),
    .B2(net601),
    .X(_02995_));
 sky130_fd_sc_hd__a221o_1 _11466_ (.A1(net587),
    .A2(t2x[5]),
    .B1(v1z[5]),
    .B2(net17),
    .C1(_02995_),
    .X(_02996_));
 sky130_fd_sc_hd__mux2_1 _11467_ (.A0(_02996_),
    .A1(net175),
    .S(net12),
    .X(_00240_));
 sky130_fd_sc_hd__a22o_1 _11468_ (.A1(net607),
    .A2(t1y[6]),
    .B1(t0x[6]),
    .B2(net601),
    .X(_02997_));
 sky130_fd_sc_hd__a221o_1 _11469_ (.A1(net588),
    .A2(t2x[6]),
    .B1(v1z[6]),
    .B2(net18),
    .C1(_02997_),
    .X(_02998_));
 sky130_fd_sc_hd__mux2_1 _11470_ (.A0(_02998_),
    .A1(net167),
    .S(net12),
    .X(_00241_));
 sky130_fd_sc_hd__a22o_1 _11471_ (.A1(net607),
    .A2(t1y[7]),
    .B1(t0x[7]),
    .B2(net601),
    .X(_02999_));
 sky130_fd_sc_hd__a221o_1 _11472_ (.A1(net588),
    .A2(t2x[7]),
    .B1(v1z[7]),
    .B2(net18),
    .C1(_02999_),
    .X(_03000_));
 sky130_fd_sc_hd__mux2_1 _11473_ (.A0(_03000_),
    .A1(net162),
    .S(net14),
    .X(_00242_));
 sky130_fd_sc_hd__a22o_1 _11474_ (.A1(net608),
    .A2(t1y[8]),
    .B1(t0x[8]),
    .B2(net602),
    .X(_03001_));
 sky130_fd_sc_hd__a221o_1 _11475_ (.A1(net588),
    .A2(t2x[8]),
    .B1(v1z[8]),
    .B2(net20),
    .C1(_03001_),
    .X(_03002_));
 sky130_fd_sc_hd__mux2_1 _11476_ (.A0(_03002_),
    .A1(net157),
    .S(net14),
    .X(_00243_));
 sky130_fd_sc_hd__a22o_1 _11477_ (.A1(net608),
    .A2(t1y[9]),
    .B1(t0x[9]),
    .B2(net602),
    .X(_03003_));
 sky130_fd_sc_hd__a221o_1 _11478_ (.A1(net588),
    .A2(t2x[9]),
    .B1(v1z[9]),
    .B2(net20),
    .C1(_03003_),
    .X(_03004_));
 sky130_fd_sc_hd__mux2_1 _11479_ (.A0(_03004_),
    .A1(net152),
    .S(net14),
    .X(_00244_));
 sky130_fd_sc_hd__a22o_1 _11480_ (.A1(net608),
    .A2(t1y[10]),
    .B1(t0x[10]),
    .B2(net602),
    .X(_03005_));
 sky130_fd_sc_hd__a221o_1 _11481_ (.A1(net588),
    .A2(t2x[10]),
    .B1(v1z[10]),
    .B2(net20),
    .C1(_03005_),
    .X(_03006_));
 sky130_fd_sc_hd__mux2_1 _11482_ (.A0(_03006_),
    .A1(net147),
    .S(net14),
    .X(_00245_));
 sky130_fd_sc_hd__a22o_1 _11483_ (.A1(net608),
    .A2(t1y[11]),
    .B1(t0x[11]),
    .B2(net602),
    .X(_03007_));
 sky130_fd_sc_hd__a221o_1 _11484_ (.A1(net588),
    .A2(t2x[11]),
    .B1(v1z[11]),
    .B2(net20),
    .C1(_03007_),
    .X(_03008_));
 sky130_fd_sc_hd__mux2_1 _11485_ (.A0(_03008_),
    .A1(net144),
    .S(net14),
    .X(_00246_));
 sky130_fd_sc_hd__a22o_1 _11486_ (.A1(net608),
    .A2(t1y[12]),
    .B1(t0x[12]),
    .B2(net602),
    .X(_03009_));
 sky130_fd_sc_hd__a221o_1 _11487_ (.A1(net589),
    .A2(t2x[12]),
    .B1(v1z[12]),
    .B2(net20),
    .C1(_03009_),
    .X(_03010_));
 sky130_fd_sc_hd__mux2_1 _11488_ (.A0(_03010_),
    .A1(net138),
    .S(net14),
    .X(_00247_));
 sky130_fd_sc_hd__a22o_1 _11489_ (.A1(net608),
    .A2(t1y[13]),
    .B1(t0x[13]),
    .B2(net602),
    .X(_03011_));
 sky130_fd_sc_hd__a221o_1 _11490_ (.A1(net589),
    .A2(t2x[13]),
    .B1(v1z[13]),
    .B2(net20),
    .C1(_03011_),
    .X(_03012_));
 sky130_fd_sc_hd__mux2_1 _11491_ (.A0(_03012_),
    .A1(net133),
    .S(net14),
    .X(_00248_));
 sky130_fd_sc_hd__a22o_1 _11492_ (.A1(net609),
    .A2(t1y[14]),
    .B1(t0x[14]),
    .B2(net602),
    .X(_03013_));
 sky130_fd_sc_hd__a221o_1 _11493_ (.A1(net589),
    .A2(t2x[14]),
    .B1(v1z[14]),
    .B2(net20),
    .C1(_03013_),
    .X(_03014_));
 sky130_fd_sc_hd__mux2_1 _11494_ (.A0(_03014_),
    .A1(net129),
    .S(net14),
    .X(_00249_));
 sky130_fd_sc_hd__a22o_1 _11495_ (.A1(net608),
    .A2(t1y[15]),
    .B1(t0x[15]),
    .B2(net602),
    .X(_03015_));
 sky130_fd_sc_hd__a221o_1 _11496_ (.A1(net588),
    .A2(t2x[15]),
    .B1(v1z[15]),
    .B2(net20),
    .C1(_03015_),
    .X(_03016_));
 sky130_fd_sc_hd__mux2_1 _11497_ (.A0(_03016_),
    .A1(net124),
    .S(net14),
    .X(_00250_));
 sky130_fd_sc_hd__a22o_1 _11498_ (.A1(net608),
    .A2(t1y[16]),
    .B1(t0x[16]),
    .B2(net603),
    .X(_03017_));
 sky130_fd_sc_hd__a221o_1 _11499_ (.A1(net588),
    .A2(t2x[16]),
    .B1(v1z[16]),
    .B2(net20),
    .C1(_03017_),
    .X(_03018_));
 sky130_fd_sc_hd__mux2_1 _11500_ (.A0(_03018_),
    .A1(net119),
    .S(net14),
    .X(_00251_));
 sky130_fd_sc_hd__a22o_1 _11501_ (.A1(net609),
    .A2(t1y[17]),
    .B1(t0x[17]),
    .B2(net602),
    .X(_03019_));
 sky130_fd_sc_hd__a221o_1 _11502_ (.A1(net588),
    .A2(t2x[17]),
    .B1(v1z[17]),
    .B2(net20),
    .C1(_03019_),
    .X(_03020_));
 sky130_fd_sc_hd__mux2_1 _11503_ (.A0(_03020_),
    .A1(net115),
    .S(net14),
    .X(_00252_));
 sky130_fd_sc_hd__a22o_1 _11504_ (.A1(net609),
    .A2(t1y[18]),
    .B1(t0x[18]),
    .B2(net603),
    .X(_03021_));
 sky130_fd_sc_hd__a221o_1 _11505_ (.A1(net591),
    .A2(t2x[18]),
    .B1(v1z[18]),
    .B2(net21),
    .C1(_03021_),
    .X(_03022_));
 sky130_fd_sc_hd__mux2_1 _11506_ (.A0(_03022_),
    .A1(net108),
    .S(net15),
    .X(_00253_));
 sky130_fd_sc_hd__a22o_1 _11507_ (.A1(net609),
    .A2(t1y[19]),
    .B1(t0x[19]),
    .B2(net603),
    .X(_03023_));
 sky130_fd_sc_hd__a221o_1 _11508_ (.A1(net591),
    .A2(t2x[19]),
    .B1(v1z[19]),
    .B2(net21),
    .C1(_03023_),
    .X(_03024_));
 sky130_fd_sc_hd__mux2_1 _11509_ (.A0(_03024_),
    .A1(net103),
    .S(net14),
    .X(_00254_));
 sky130_fd_sc_hd__a22o_1 _11510_ (.A1(net610),
    .A2(t1y[20]),
    .B1(t0x[20]),
    .B2(net604),
    .X(_03025_));
 sky130_fd_sc_hd__a221o_1 _11511_ (.A1(net591),
    .A2(t2x[20]),
    .B1(v1z[20]),
    .B2(net21),
    .C1(_03025_),
    .X(_03026_));
 sky130_fd_sc_hd__mux2_1 _11512_ (.A0(_03026_),
    .A1(net99),
    .S(net14),
    .X(_00255_));
 sky130_fd_sc_hd__a22o_1 _11513_ (.A1(net610),
    .A2(t1y[21]),
    .B1(t0x[21]),
    .B2(net604),
    .X(_03027_));
 sky130_fd_sc_hd__a221o_1 _11514_ (.A1(net591),
    .A2(t2x[21]),
    .B1(v1z[21]),
    .B2(net21),
    .C1(_03027_),
    .X(_03028_));
 sky130_fd_sc_hd__mux2_1 _11515_ (.A0(_03028_),
    .A1(net93),
    .S(net14),
    .X(_00256_));
 sky130_fd_sc_hd__a22o_1 _11516_ (.A1(net610),
    .A2(t1y[22]),
    .B1(t0x[22]),
    .B2(net604),
    .X(_03029_));
 sky130_fd_sc_hd__a221o_1 _11517_ (.A1(net591),
    .A2(t2x[22]),
    .B1(v1z[22]),
    .B2(net21),
    .C1(_03029_),
    .X(_03030_));
 sky130_fd_sc_hd__mux2_1 _11518_ (.A0(_03030_),
    .A1(net89),
    .S(net14),
    .X(_00257_));
 sky130_fd_sc_hd__a22o_1 _11519_ (.A1(net610),
    .A2(t1y[23]),
    .B1(t0x[23]),
    .B2(net604),
    .X(_03031_));
 sky130_fd_sc_hd__a221o_1 _11520_ (.A1(net591),
    .A2(t2x[23]),
    .B1(v1z[23]),
    .B2(net21),
    .C1(_03031_),
    .X(_03032_));
 sky130_fd_sc_hd__mux2_1 _11521_ (.A0(_03032_),
    .A1(net85),
    .S(net14),
    .X(_00258_));
 sky130_fd_sc_hd__a22o_1 _11522_ (.A1(net610),
    .A2(t1y[24]),
    .B1(t0x[24]),
    .B2(net604),
    .X(_03033_));
 sky130_fd_sc_hd__a221o_1 _11523_ (.A1(net590),
    .A2(t2x[24]),
    .B1(v1z[24]),
    .B2(net21),
    .C1(_03033_),
    .X(_03034_));
 sky130_fd_sc_hd__mux2_1 _11524_ (.A0(_03034_),
    .A1(net81),
    .S(net15),
    .X(_00259_));
 sky130_fd_sc_hd__a22o_1 _11525_ (.A1(net611),
    .A2(t1y[25]),
    .B1(t0x[25]),
    .B2(net604),
    .X(_03035_));
 sky130_fd_sc_hd__a221o_1 _11526_ (.A1(net590),
    .A2(t2x[25]),
    .B1(v1z[25]),
    .B2(net21),
    .C1(_03035_),
    .X(_03036_));
 sky130_fd_sc_hd__mux2_1 _11527_ (.A0(_03036_),
    .A1(net78),
    .S(net15),
    .X(_00260_));
 sky130_fd_sc_hd__a22o_1 _11528_ (.A1(net610),
    .A2(t1y[26]),
    .B1(t0x[26]),
    .B2(net604),
    .X(_03037_));
 sky130_fd_sc_hd__a221o_1 _11529_ (.A1(net590),
    .A2(t2x[26]),
    .B1(v1z[26]),
    .B2(net21),
    .C1(_03037_),
    .X(_03038_));
 sky130_fd_sc_hd__mux2_1 _11530_ (.A0(_03038_),
    .A1(net75),
    .S(net15),
    .X(_00261_));
 sky130_fd_sc_hd__a22o_1 _11531_ (.A1(net611),
    .A2(t1y[27]),
    .B1(t0x[27]),
    .B2(net604),
    .X(_03039_));
 sky130_fd_sc_hd__a221o_1 _11532_ (.A1(net590),
    .A2(t2x[27]),
    .B1(v1z[27]),
    .B2(net21),
    .C1(_03039_),
    .X(_03040_));
 sky130_fd_sc_hd__mux2_1 _11533_ (.A0(_03040_),
    .A1(net74),
    .S(net15),
    .X(_00262_));
 sky130_fd_sc_hd__a22o_1 _11534_ (.A1(net611),
    .A2(t1y[28]),
    .B1(t0x[28]),
    .B2(net604),
    .X(_03041_));
 sky130_fd_sc_hd__a221o_1 _11535_ (.A1(net590),
    .A2(t2x[28]),
    .B1(v1z[28]),
    .B2(net20),
    .C1(_03041_),
    .X(_03042_));
 sky130_fd_sc_hd__mux2_1 _11536_ (.A0(_03042_),
    .A1(net71),
    .S(net15),
    .X(_00263_));
 sky130_fd_sc_hd__a22o_1 _11537_ (.A1(net611),
    .A2(t1y[29]),
    .B1(t0x[29]),
    .B2(net605),
    .X(_03043_));
 sky130_fd_sc_hd__a221o_1 _11538_ (.A1(net590),
    .A2(t2x[29]),
    .B1(v1z[29]),
    .B2(net20),
    .C1(_03043_),
    .X(_03044_));
 sky130_fd_sc_hd__mux2_1 _11539_ (.A0(_03044_),
    .A1(net68),
    .S(net15),
    .X(_00264_));
 sky130_fd_sc_hd__a22o_1 _11540_ (.A1(net611),
    .A2(t1y[30]),
    .B1(t0x[30]),
    .B2(net605),
    .X(_03045_));
 sky130_fd_sc_hd__a221o_1 _11541_ (.A1(net590),
    .A2(t2x[30]),
    .B1(v1z[30]),
    .B2(net21),
    .C1(_03045_),
    .X(_03046_));
 sky130_fd_sc_hd__mux2_1 _11542_ (.A0(_03046_),
    .A1(net65),
    .S(net15),
    .X(_00265_));
 sky130_fd_sc_hd__a22o_1 _11543_ (.A1(net611),
    .A2(t1y[31]),
    .B1(t0x[31]),
    .B2(net605),
    .X(_03047_));
 sky130_fd_sc_hd__a221o_1 _11544_ (.A1(net590),
    .A2(t2x[31]),
    .B1(v1z[31]),
    .B2(net21),
    .C1(_03047_),
    .X(_03048_));
 sky130_fd_sc_hd__mux2_1 _11545_ (.A0(_03048_),
    .A1(net62),
    .S(net15),
    .X(_00266_));
 sky130_fd_sc_hd__nor2_8 _11546_ (.A(net599),
    .B(_02822_),
    .Y(_03049_));
 sky130_fd_sc_hd__or2_2 _11547_ (.A(net599),
    .B(_02822_),
    .X(_03050_));
 sky130_fd_sc_hd__nor2_1 _11548_ (.A(net592),
    .B(\state[9] ),
    .Y(_03051_));
 sky130_fd_sc_hd__or2_4 _11549_ (.A(net592),
    .B(\state[9] ),
    .X(_03052_));
 sky130_fd_sc_hd__nor2_1 _11550_ (.A(net10),
    .B(_03052_),
    .Y(_03053_));
 sky130_fd_sc_hd__nand2_2 _11551_ (.A(_03049_),
    .B(net43),
    .Y(_03054_));
 sky130_fd_sc_hd__o21a_4 _11552_ (.A1(net595),
    .A2(_03054_),
    .B1(net645),
    .X(_03055_));
 sky130_fd_sc_hd__o21ai_4 _11553_ (.A1(net595),
    .A2(_03054_),
    .B1(net645),
    .Y(_03056_));
 sky130_fd_sc_hd__nor2_4 _11554_ (.A(\state[9] ),
    .B(_02822_),
    .Y(_03057_));
 sky130_fd_sc_hd__or2_4 _11555_ (.A(\state[9] ),
    .B(_02822_),
    .X(_03058_));
 sky130_fd_sc_hd__and3_1 _11556_ (.A(net435),
    .B(net431),
    .C(net540),
    .X(_03059_));
 sky130_fd_sc_hd__and4_1 _11557_ (.A(net435),
    .B(net430),
    .C(net535),
    .D(net540),
    .X(_03060_));
 sky130_fd_sc_hd__nand2_1 _11558_ (.A(net426),
    .B(net544),
    .Y(_03061_));
 sky130_fd_sc_hd__a22o_1 _11559_ (.A1(net435),
    .A2(net535),
    .B1(net540),
    .B2(net430),
    .X(_03062_));
 sky130_fd_sc_hd__and2b_1 _11560_ (.A_N(_03060_),
    .B(_03062_),
    .X(_03063_));
 sky130_fd_sc_hd__a31o_1 _11561_ (.A1(net426),
    .A2(net544),
    .A3(_03062_),
    .B1(_03060_),
    .X(_03064_));
 sky130_fd_sc_hd__nand2_1 _11562_ (.A(net413),
    .B(net552),
    .Y(_03065_));
 sky130_fd_sc_hd__a22o_1 _11563_ (.A1(net421),
    .A2(net545),
    .B1(net548),
    .B2(net417),
    .X(_03066_));
 sky130_fd_sc_hd__and3_1 _11564_ (.A(net421),
    .B(net417),
    .C(net548),
    .X(_03067_));
 sky130_fd_sc_hd__a21bo_1 _11565_ (.A1(net545),
    .A2(_03067_),
    .B1_N(_03066_),
    .X(_03068_));
 sky130_fd_sc_hd__xor2_2 _11566_ (.A(_03065_),
    .B(_03068_),
    .X(_03069_));
 sky130_fd_sc_hd__nand2_1 _11567_ (.A(_03064_),
    .B(_03069_),
    .Y(_03070_));
 sky130_fd_sc_hd__and4_1 _11568_ (.A(net421),
    .B(net417),
    .C(net548),
    .D(net552),
    .X(_03071_));
 sky130_fd_sc_hd__nand2_1 _11569_ (.A(net413),
    .B(net558),
    .Y(_03072_));
 sky130_fd_sc_hd__a22o_1 _11570_ (.A1(net421),
    .A2(net548),
    .B1(net552),
    .B2(net417),
    .X(_03073_));
 sky130_fd_sc_hd__and2b_1 _11571_ (.A_N(_03071_),
    .B(_03073_),
    .X(_03074_));
 sky130_fd_sc_hd__a31o_1 _11572_ (.A1(net413),
    .A2(net558),
    .A3(_03073_),
    .B1(_03071_),
    .X(_03075_));
 sky130_fd_sc_hd__xor2_2 _11573_ (.A(_03064_),
    .B(_03069_),
    .X(_03076_));
 sky130_fd_sc_hd__nand2_1 _11574_ (.A(_03075_),
    .B(_03076_),
    .Y(_03077_));
 sky130_fd_sc_hd__nand2_1 _11575_ (.A(net400),
    .B(net564),
    .Y(_03078_));
 sky130_fd_sc_hd__a22o_1 _11576_ (.A1(net412),
    .A2(net552),
    .B1(net560),
    .B2(net405),
    .X(_03079_));
 sky130_fd_sc_hd__and3_1 _11577_ (.A(net408),
    .B(net404),
    .C(net560),
    .X(_03080_));
 sky130_fd_sc_hd__a21bo_1 _11578_ (.A1(net552),
    .A2(_03080_),
    .B1_N(_03079_),
    .X(_03081_));
 sky130_fd_sc_hd__xor2_2 _11579_ (.A(_03078_),
    .B(_03081_),
    .X(_03082_));
 sky130_fd_sc_hd__and4_1 _11580_ (.A(net408),
    .B(net404),
    .C(net560),
    .D(net564),
    .X(_03083_));
 sky130_fd_sc_hd__nand2_1 _11581_ (.A(net400),
    .B(net567),
    .Y(_03084_));
 sky130_fd_sc_hd__a22o_1 _11582_ (.A1(net408),
    .A2(net560),
    .B1(net564),
    .B2(net404),
    .X(_03085_));
 sky130_fd_sc_hd__and2b_1 _11583_ (.A_N(_03083_),
    .B(_03085_),
    .X(_03086_));
 sky130_fd_sc_hd__a31o_1 _11584_ (.A1(net400),
    .A2(net567),
    .A3(_03085_),
    .B1(_03083_),
    .X(_03087_));
 sky130_fd_sc_hd__xor2_1 _11585_ (.A(_03082_),
    .B(_03087_),
    .X(_03088_));
 sky130_fd_sc_hd__a22o_1 _11586_ (.A1(net396),
    .A2(net567),
    .B1(net572),
    .B2(net390),
    .X(_03089_));
 sky130_fd_sc_hd__and4_1 _11587_ (.A(net396),
    .B(net390),
    .C(net567),
    .D(net575),
    .X(_03090_));
 sky130_fd_sc_hd__inv_2 _11588_ (.A(_03090_),
    .Y(_03091_));
 sky130_fd_sc_hd__and4_1 _11589_ (.A(net386),
    .B(net577),
    .C(_03089_),
    .D(_03091_),
    .X(_03092_));
 sky130_fd_sc_hd__a22oi_1 _11590_ (.A1(net386),
    .A2(net577),
    .B1(_03089_),
    .B2(_03091_),
    .Y(_03093_));
 sky130_fd_sc_hd__nor2_1 _11591_ (.A(_03092_),
    .B(_03093_),
    .Y(_03094_));
 sky130_fd_sc_hd__and2_1 _11592_ (.A(_03088_),
    .B(_03094_),
    .X(_03095_));
 sky130_fd_sc_hd__xnor2_1 _11593_ (.A(_03088_),
    .B(_03094_),
    .Y(_03096_));
 sky130_fd_sc_hd__a21o_1 _11594_ (.A1(_03070_),
    .A2(_03077_),
    .B1(_03096_),
    .X(_03097_));
 sky130_fd_sc_hd__xnor2_1 _11595_ (.A(_03084_),
    .B(_03086_),
    .Y(_03098_));
 sky130_fd_sc_hd__and4_1 _11596_ (.A(net408),
    .B(net404),
    .C(net564),
    .D(net567),
    .X(_03099_));
 sky130_fd_sc_hd__nand2_1 _11597_ (.A(net400),
    .B(net572),
    .Y(_03100_));
 sky130_fd_sc_hd__a22o_1 _11598_ (.A1(net408),
    .A2(net564),
    .B1(net567),
    .B2(net404),
    .X(_03101_));
 sky130_fd_sc_hd__and2b_1 _11599_ (.A_N(_03099_),
    .B(_03101_),
    .X(_03102_));
 sky130_fd_sc_hd__a31o_1 _11600_ (.A1(net400),
    .A2(net572),
    .A3(_03101_),
    .B1(_03099_),
    .X(_03103_));
 sky130_fd_sc_hd__and2_1 _11601_ (.A(_03098_),
    .B(_03103_),
    .X(_03104_));
 sky130_fd_sc_hd__xor2_1 _11602_ (.A(_03098_),
    .B(_03103_),
    .X(_03105_));
 sky130_fd_sc_hd__a22o_1 _11603_ (.A1(net396),
    .A2(net572),
    .B1(net577),
    .B2(net390),
    .X(_03106_));
 sky130_fd_sc_hd__and4_1 _11604_ (.A(net396),
    .B(net390),
    .C(net575),
    .D(net577),
    .X(_03107_));
 sky130_fd_sc_hd__inv_2 _11605_ (.A(_03107_),
    .Y(_03108_));
 sky130_fd_sc_hd__and4_1 _11606_ (.A(net386),
    .B(net581),
    .C(_03106_),
    .D(_03108_),
    .X(_03109_));
 sky130_fd_sc_hd__a22oi_1 _11607_ (.A1(net386),
    .A2(net581),
    .B1(_03106_),
    .B2(_03108_),
    .Y(_03110_));
 sky130_fd_sc_hd__nor2_1 _11608_ (.A(_03109_),
    .B(_03110_),
    .Y(_03111_));
 sky130_fd_sc_hd__and2_1 _11609_ (.A(_03105_),
    .B(_03111_),
    .X(_03112_));
 sky130_fd_sc_hd__nand3_2 _11610_ (.A(_03070_),
    .B(_03077_),
    .C(_03096_),
    .Y(_03113_));
 sky130_fd_sc_hd__o211ai_4 _11611_ (.A1(_03104_),
    .A2(_03112_),
    .B1(_03113_),
    .C1(_03097_),
    .Y(_03114_));
 sky130_fd_sc_hd__nor2_1 _11612_ (.A(_03107_),
    .B(_03109_),
    .Y(_03115_));
 sky130_fd_sc_hd__nand2_1 _11613_ (.A(net381),
    .B(net581),
    .Y(_03116_));
 sky130_fd_sc_hd__or2_1 _11614_ (.A(_03115_),
    .B(_03116_),
    .X(_03117_));
 sky130_fd_sc_hd__a22o_1 _11615_ (.A1(net577),
    .A2(net381),
    .B1(net375),
    .B2(net584),
    .X(_03118_));
 sky130_fd_sc_hd__and4_1 _11616_ (.A(net577),
    .B(net381),
    .C(net375),
    .D(net581),
    .X(_03119_));
 sky130_fd_sc_hd__nand4_2 _11617_ (.A(net577),
    .B(net381),
    .C(net375),
    .D(net582),
    .Y(_03120_));
 sky130_fd_sc_hd__o211a_1 _11618_ (.A1(_03090_),
    .A2(_03092_),
    .B1(_03118_),
    .C1(_03120_),
    .X(_03121_));
 sky130_fd_sc_hd__o211ai_1 _11619_ (.A1(_03090_),
    .A2(_03092_),
    .B1(_03118_),
    .C1(_03120_),
    .Y(_03122_));
 sky130_fd_sc_hd__a211o_1 _11620_ (.A1(_03118_),
    .A2(_03120_),
    .B1(_03090_),
    .C1(_03092_),
    .X(_03123_));
 sky130_fd_sc_hd__nand2_1 _11621_ (.A(_03122_),
    .B(_03123_),
    .Y(_03124_));
 sky130_fd_sc_hd__or2_1 _11622_ (.A(_03117_),
    .B(_03124_),
    .X(_03125_));
 sky130_fd_sc_hd__xnor2_1 _11623_ (.A(_03117_),
    .B(_03124_),
    .Y(_03126_));
 sky130_fd_sc_hd__a21oi_1 _11624_ (.A1(_03097_),
    .A2(_03114_),
    .B1(_03126_),
    .Y(_03127_));
 sky130_fd_sc_hd__and4_1 _11625_ (.A(net435),
    .B(net430),
    .C(net530),
    .D(net535),
    .X(_03128_));
 sky130_fd_sc_hd__a22oi_1 _11626_ (.A1(net435),
    .A2(net530),
    .B1(net536),
    .B2(net430),
    .Y(_03129_));
 sky130_fd_sc_hd__and4bb_1 _11627_ (.A_N(_03128_),
    .B_N(_03129_),
    .C(net426),
    .D(net540),
    .X(_03130_));
 sky130_fd_sc_hd__a22o_1 _11628_ (.A1(net421),
    .A2(net540),
    .B1(net544),
    .B2(net417),
    .X(_03131_));
 sky130_fd_sc_hd__nand4_2 _11629_ (.A(net421),
    .B(net417),
    .C(net540),
    .D(net544),
    .Y(_03132_));
 sky130_fd_sc_hd__nand4_2 _11630_ (.A(net413),
    .B(net548),
    .C(_03131_),
    .D(_03132_),
    .Y(_03133_));
 sky130_fd_sc_hd__a22o_1 _11631_ (.A1(net413),
    .A2(net548),
    .B1(_03131_),
    .B2(_03132_),
    .X(_03134_));
 sky130_fd_sc_hd__o211a_1 _11632_ (.A1(_03128_),
    .A2(_03130_),
    .B1(_03133_),
    .C1(_03134_),
    .X(_03135_));
 sky130_fd_sc_hd__a32o_1 _11633_ (.A1(net413),
    .A2(net552),
    .A3(_03066_),
    .B1(_03067_),
    .B2(net545),
    .X(_03136_));
 sky130_fd_sc_hd__a211o_1 _11634_ (.A1(_03133_),
    .A2(_03134_),
    .B1(_03128_),
    .C1(_03130_),
    .X(_03137_));
 sky130_fd_sc_hd__nand2b_1 _11635_ (.A_N(_03135_),
    .B(_03137_),
    .Y(_03138_));
 sky130_fd_sc_hd__a21o_1 _11636_ (.A1(_03136_),
    .A2(_03137_),
    .B1(_03135_),
    .X(_03139_));
 sky130_fd_sc_hd__and2_1 _11637_ (.A(net400),
    .B(net557),
    .X(_03140_));
 sky130_fd_sc_hd__a22o_1 _11638_ (.A1(net548),
    .A2(net408),
    .B1(net405),
    .B2(net552),
    .X(_03141_));
 sky130_fd_sc_hd__nand4_1 _11639_ (.A(net548),
    .B(net408),
    .C(net405),
    .D(net552),
    .Y(_03142_));
 sky130_fd_sc_hd__nand3_1 _11640_ (.A(_03140_),
    .B(_03141_),
    .C(_03142_),
    .Y(_03143_));
 sky130_fd_sc_hd__a21o_1 _11641_ (.A1(_03141_),
    .A2(_03142_),
    .B1(_03140_),
    .X(_03144_));
 sky130_fd_sc_hd__a32o_1 _11642_ (.A1(net400),
    .A2(net564),
    .A3(_03079_),
    .B1(_03080_),
    .B2(net552),
    .X(_03145_));
 sky130_fd_sc_hd__nand3_2 _11643_ (.A(_03143_),
    .B(_03144_),
    .C(_03145_),
    .Y(_03146_));
 sky130_fd_sc_hd__a21o_1 _11644_ (.A1(_03143_),
    .A2(_03144_),
    .B1(_03145_),
    .X(_03147_));
 sky130_fd_sc_hd__nand2_1 _11645_ (.A(net386),
    .B(net572),
    .Y(_03148_));
 sky130_fd_sc_hd__a22oi_1 _11646_ (.A1(net396),
    .A2(net564),
    .B1(net567),
    .B2(net390),
    .Y(_03149_));
 sky130_fd_sc_hd__and4_1 _11647_ (.A(net396),
    .B(net390),
    .C(net564),
    .D(net567),
    .X(_03150_));
 sky130_fd_sc_hd__nor2_1 _11648_ (.A(_03149_),
    .B(_03150_),
    .Y(_03151_));
 sky130_fd_sc_hd__xnor2_1 _11649_ (.A(_03148_),
    .B(_03151_),
    .Y(_03152_));
 sky130_fd_sc_hd__nand3_2 _11650_ (.A(_03146_),
    .B(_03147_),
    .C(_03152_),
    .Y(_03153_));
 sky130_fd_sc_hd__a21o_1 _11651_ (.A1(_03146_),
    .A2(_03147_),
    .B1(_03152_),
    .X(_03154_));
 sky130_fd_sc_hd__nand3_1 _11652_ (.A(_03139_),
    .B(_03153_),
    .C(_03154_),
    .Y(_03155_));
 sky130_fd_sc_hd__a21oi_2 _11653_ (.A1(_03082_),
    .A2(_03087_),
    .B1(_03095_),
    .Y(_03156_));
 sky130_fd_sc_hd__a21o_1 _11654_ (.A1(_03153_),
    .A2(_03154_),
    .B1(_03139_),
    .X(_03157_));
 sky130_fd_sc_hd__nand2_1 _11655_ (.A(_03155_),
    .B(_03157_),
    .Y(_03158_));
 sky130_fd_sc_hd__o21ai_2 _11656_ (.A1(_03156_),
    .A2(_03158_),
    .B1(_03155_),
    .Y(_03159_));
 sky130_fd_sc_hd__a31o_1 _11657_ (.A1(net386),
    .A2(net575),
    .A3(_03151_),
    .B1(_03150_),
    .X(_03160_));
 sky130_fd_sc_hd__nand2_1 _11658_ (.A(net371),
    .B(net581),
    .Y(_03161_));
 sky130_fd_sc_hd__and4_1 _11659_ (.A(net572),
    .B(net580),
    .C(net381),
    .D(net375),
    .X(_03162_));
 sky130_fd_sc_hd__a22o_1 _11660_ (.A1(net572),
    .A2(net381),
    .B1(net375),
    .B2(net580),
    .X(_03163_));
 sky130_fd_sc_hd__and2b_1 _11661_ (.A_N(_03162_),
    .B(_03163_),
    .X(_03164_));
 sky130_fd_sc_hd__xnor2_1 _11662_ (.A(_03161_),
    .B(_03164_),
    .Y(_03165_));
 sky130_fd_sc_hd__or2_1 _11663_ (.A(_03160_),
    .B(_03165_),
    .X(_03166_));
 sky130_fd_sc_hd__and2_1 _11664_ (.A(_03160_),
    .B(_03165_),
    .X(_03167_));
 sky130_fd_sc_hd__inv_2 _11665_ (.A(_03167_),
    .Y(_03168_));
 sky130_fd_sc_hd__nand2_1 _11666_ (.A(_03166_),
    .B(_03168_),
    .Y(_03169_));
 sky130_fd_sc_hd__nor2_1 _11667_ (.A(_03119_),
    .B(_03121_),
    .Y(_03170_));
 sky130_fd_sc_hd__xnor2_1 _11668_ (.A(_03169_),
    .B(_03170_),
    .Y(_03171_));
 sky130_fd_sc_hd__and2b_1 _11669_ (.A_N(_03171_),
    .B(_03159_),
    .X(_03172_));
 sky130_fd_sc_hd__xor2_1 _11670_ (.A(_03159_),
    .B(_03171_),
    .X(_03173_));
 sky130_fd_sc_hd__nor2_1 _11671_ (.A(_03125_),
    .B(_03173_),
    .Y(_03174_));
 sky130_fd_sc_hd__xor2_1 _11672_ (.A(_03125_),
    .B(_03173_),
    .X(_03175_));
 sky130_fd_sc_hd__and4_1 _11673_ (.A(net435),
    .B(net430),
    .C(net525),
    .D(net530),
    .X(_03176_));
 sky130_fd_sc_hd__nand2_1 _11674_ (.A(net426),
    .B(net535),
    .Y(_03177_));
 sky130_fd_sc_hd__a22o_1 _11675_ (.A1(net435),
    .A2(net525),
    .B1(net530),
    .B2(net430),
    .X(_03178_));
 sky130_fd_sc_hd__and2b_1 _11676_ (.A_N(_03176_),
    .B(_03178_),
    .X(_03179_));
 sky130_fd_sc_hd__a31o_1 _11677_ (.A1(net426),
    .A2(net535),
    .A3(_03178_),
    .B1(_03176_),
    .X(_03180_));
 sky130_fd_sc_hd__a22o_1 _11678_ (.A1(net421),
    .A2(net536),
    .B1(net541),
    .B2(net417),
    .X(_03181_));
 sky130_fd_sc_hd__nand4_2 _11679_ (.A(net421),
    .B(net417),
    .C(net536),
    .D(net540),
    .Y(_03182_));
 sky130_fd_sc_hd__nand4_2 _11680_ (.A(net413),
    .B(net545),
    .C(_03181_),
    .D(_03182_),
    .Y(_03183_));
 sky130_fd_sc_hd__a22o_1 _11681_ (.A1(net413),
    .A2(net545),
    .B1(_03181_),
    .B2(_03182_),
    .X(_03184_));
 sky130_fd_sc_hd__nand3_1 _11682_ (.A(_03180_),
    .B(_03183_),
    .C(_03184_),
    .Y(_03185_));
 sky130_fd_sc_hd__nand2_1 _11683_ (.A(_03132_),
    .B(_03133_),
    .Y(_03186_));
 sky130_fd_sc_hd__a21o_1 _11684_ (.A1(_03183_),
    .A2(_03184_),
    .B1(_03180_),
    .X(_03187_));
 sky130_fd_sc_hd__and3_1 _11685_ (.A(_03185_),
    .B(_03186_),
    .C(_03187_),
    .X(_03188_));
 sky130_fd_sc_hd__a21bo_1 _11686_ (.A1(_03186_),
    .A2(_03187_),
    .B1_N(_03185_),
    .X(_03189_));
 sky130_fd_sc_hd__nand2_1 _11687_ (.A(net386),
    .B(net567),
    .Y(_03190_));
 sky130_fd_sc_hd__and4_1 _11688_ (.A(net560),
    .B(net396),
    .C(net390),
    .D(net564),
    .X(_03191_));
 sky130_fd_sc_hd__a22o_1 _11689_ (.A1(net560),
    .A2(net396),
    .B1(net390),
    .B2(net564),
    .X(_03192_));
 sky130_fd_sc_hd__and2b_1 _11690_ (.A_N(_03191_),
    .B(_03192_),
    .X(_03193_));
 sky130_fd_sc_hd__xnor2_1 _11691_ (.A(_03190_),
    .B(_03193_),
    .Y(_03194_));
 sky130_fd_sc_hd__nand4_1 _11692_ (.A(net545),
    .B(net548),
    .C(net408),
    .D(net404),
    .Y(_03195_));
 sky130_fd_sc_hd__a22o_1 _11693_ (.A1(net545),
    .A2(net408),
    .B1(net404),
    .B2(net548),
    .X(_03196_));
 sky130_fd_sc_hd__nand4_1 _11694_ (.A(net400),
    .B(net552),
    .C(_03195_),
    .D(_03196_),
    .Y(_03197_));
 sky130_fd_sc_hd__a22o_1 _11695_ (.A1(net400),
    .A2(net552),
    .B1(_03195_),
    .B2(_03196_),
    .X(_03198_));
 sky130_fd_sc_hd__a21bo_1 _11696_ (.A1(_03140_),
    .A2(_03141_),
    .B1_N(_03142_),
    .X(_03199_));
 sky130_fd_sc_hd__nand3_1 _11697_ (.A(_03197_),
    .B(_03198_),
    .C(_03199_),
    .Y(_03200_));
 sky130_fd_sc_hd__a21o_1 _11698_ (.A1(_03197_),
    .A2(_03198_),
    .B1(_03199_),
    .X(_03201_));
 sky130_fd_sc_hd__nand3_1 _11699_ (.A(_03194_),
    .B(_03200_),
    .C(_03201_),
    .Y(_03202_));
 sky130_fd_sc_hd__a21o_1 _11700_ (.A1(_03200_),
    .A2(_03201_),
    .B1(_03194_),
    .X(_03203_));
 sky130_fd_sc_hd__and3_1 _11701_ (.A(_03189_),
    .B(_03202_),
    .C(_03203_),
    .X(_03204_));
 sky130_fd_sc_hd__a21oi_2 _11702_ (.A1(_03202_),
    .A2(_03203_),
    .B1(_03189_),
    .Y(_03205_));
 sky130_fd_sc_hd__a211oi_4 _11703_ (.A1(_03146_),
    .A2(_03153_),
    .B1(_03204_),
    .C1(_03205_),
    .Y(_03206_));
 sky130_fd_sc_hd__o211a_1 _11704_ (.A1(_03204_),
    .A2(_03205_),
    .B1(_03146_),
    .C1(_03153_),
    .X(_03207_));
 sky130_fd_sc_hd__nand2_1 _11705_ (.A(_03182_),
    .B(_03183_),
    .Y(_03208_));
 sky130_fd_sc_hd__and4_1 _11706_ (.A(net436),
    .B(net430),
    .C(net520),
    .D(net525),
    .X(_03209_));
 sky130_fd_sc_hd__a22oi_1 _11707_ (.A1(net436),
    .A2(net520),
    .B1(net525),
    .B2(net430),
    .Y(_03210_));
 sky130_fd_sc_hd__and4bb_1 _11708_ (.A_N(_03209_),
    .B_N(_03210_),
    .C(net426),
    .D(net530),
    .X(_03211_));
 sky130_fd_sc_hd__nor2_1 _11709_ (.A(_03209_),
    .B(_03211_),
    .Y(_03212_));
 sky130_fd_sc_hd__nand2_1 _11710_ (.A(net414),
    .B(net541),
    .Y(_03213_));
 sky130_fd_sc_hd__and4_1 _11711_ (.A(net530),
    .B(net422),
    .C(net418),
    .D(net536),
    .X(_03214_));
 sky130_fd_sc_hd__a22o_1 _11712_ (.A1(net530),
    .A2(net422),
    .B1(net418),
    .B2(net536),
    .X(_03215_));
 sky130_fd_sc_hd__and2b_1 _11713_ (.A_N(_03214_),
    .B(_03215_),
    .X(_03216_));
 sky130_fd_sc_hd__xnor2_2 _11714_ (.A(_03213_),
    .B(_03216_),
    .Y(_03217_));
 sky130_fd_sc_hd__nand2b_1 _11715_ (.A_N(_03212_),
    .B(_03217_),
    .Y(_03218_));
 sky130_fd_sc_hd__xnor2_2 _11716_ (.A(_03212_),
    .B(_03217_),
    .Y(_03219_));
 sky130_fd_sc_hd__nand2_1 _11717_ (.A(_03208_),
    .B(_03219_),
    .Y(_03220_));
 sky130_fd_sc_hd__xor2_2 _11718_ (.A(_03208_),
    .B(_03219_),
    .X(_03221_));
 sky130_fd_sc_hd__nand2_1 _11719_ (.A(net427),
    .B(net525),
    .Y(_03222_));
 sky130_fd_sc_hd__a22oi_2 _11720_ (.A1(net516),
    .A2(net437),
    .B1(net432),
    .B2(net520),
    .Y(_03223_));
 sky130_fd_sc_hd__and4_1 _11721_ (.A(net515),
    .B(net435),
    .C(net432),
    .D(net520),
    .X(_03224_));
 sky130_fd_sc_hd__nor2_1 _11722_ (.A(_03223_),
    .B(_03224_),
    .Y(_03225_));
 sky130_fd_sc_hd__xnor2_2 _11723_ (.A(_03222_),
    .B(_03225_),
    .Y(_03226_));
 sky130_fd_sc_hd__and2_1 _11724_ (.A(net441),
    .B(net511),
    .X(_03227_));
 sky130_fd_sc_hd__nand4_2 _11725_ (.A(net449),
    .B(net503),
    .C(net444),
    .D(net507),
    .Y(_03228_));
 sky130_fd_sc_hd__a22o_1 _11726_ (.A1(net449),
    .A2(net503),
    .B1(net444),
    .B2(net507),
    .X(_03229_));
 sky130_fd_sc_hd__nand3_1 _11727_ (.A(_03227_),
    .B(_03228_),
    .C(_03229_),
    .Y(_03230_));
 sky130_fd_sc_hd__a21o_1 _11728_ (.A1(_03228_),
    .A2(_03229_),
    .B1(_03227_),
    .X(_03231_));
 sky130_fd_sc_hd__nand4_2 _11729_ (.A(net449),
    .B(net444),
    .C(net507),
    .D(net511),
    .Y(_03232_));
 sky130_fd_sc_hd__and2_1 _11730_ (.A(net441),
    .B(net515),
    .X(_03233_));
 sky130_fd_sc_hd__a22o_1 _11731_ (.A1(net449),
    .A2(net507),
    .B1(net511),
    .B2(net444),
    .X(_03234_));
 sky130_fd_sc_hd__nand3_1 _11732_ (.A(_03232_),
    .B(_03233_),
    .C(_03234_),
    .Y(_03235_));
 sky130_fd_sc_hd__a21bo_1 _11733_ (.A1(_03233_),
    .A2(_03234_),
    .B1_N(_03232_),
    .X(_03236_));
 sky130_fd_sc_hd__nand3_2 _11734_ (.A(_03230_),
    .B(_03231_),
    .C(_03236_),
    .Y(_03237_));
 sky130_fd_sc_hd__a21o_1 _11735_ (.A1(_03230_),
    .A2(_03231_),
    .B1(_03236_),
    .X(_03238_));
 sky130_fd_sc_hd__nand3_2 _11736_ (.A(_03226_),
    .B(_03237_),
    .C(_03238_),
    .Y(_03239_));
 sky130_fd_sc_hd__a21o_1 _11737_ (.A1(_03237_),
    .A2(_03238_),
    .B1(_03226_),
    .X(_03240_));
 sky130_fd_sc_hd__nand4_1 _11738_ (.A(net448),
    .B(net444),
    .C(net511),
    .D(net515),
    .Y(_03241_));
 sky130_fd_sc_hd__and2_1 _11739_ (.A(net441),
    .B(net520),
    .X(_03242_));
 sky130_fd_sc_hd__a22o_1 _11740_ (.A1(net448),
    .A2(net511),
    .B1(net515),
    .B2(net443),
    .X(_03243_));
 sky130_fd_sc_hd__nand3_1 _11741_ (.A(_03241_),
    .B(_03242_),
    .C(_03243_),
    .Y(_03244_));
 sky130_fd_sc_hd__a21bo_1 _11742_ (.A1(_03242_),
    .A2(_03243_),
    .B1_N(_03241_),
    .X(_03245_));
 sky130_fd_sc_hd__a21o_1 _11743_ (.A1(_03232_),
    .A2(_03234_),
    .B1(_03233_),
    .X(_03246_));
 sky130_fd_sc_hd__nand3_2 _11744_ (.A(_03235_),
    .B(_03245_),
    .C(_03246_),
    .Y(_03247_));
 sky130_fd_sc_hd__a21o_1 _11745_ (.A1(_03235_),
    .A2(_03246_),
    .B1(_03245_),
    .X(_03248_));
 sky130_fd_sc_hd__o2bb2a_1 _11746_ (.A1_N(net427),
    .A2_N(net530),
    .B1(_03209_),
    .B2(_03210_),
    .X(_03249_));
 sky130_fd_sc_hd__nor2_1 _11747_ (.A(_03211_),
    .B(_03249_),
    .Y(_03250_));
 sky130_fd_sc_hd__nand3_2 _11748_ (.A(_03247_),
    .B(_03248_),
    .C(_03250_),
    .Y(_03251_));
 sky130_fd_sc_hd__a21bo_1 _11749_ (.A1(_03248_),
    .A2(_03250_),
    .B1_N(_03247_),
    .X(_03252_));
 sky130_fd_sc_hd__nand3_4 _11750_ (.A(_03239_),
    .B(_03240_),
    .C(_03252_),
    .Y(_03253_));
 sky130_fd_sc_hd__a21o_1 _11751_ (.A1(_03239_),
    .A2(_03240_),
    .B1(_03252_),
    .X(_03254_));
 sky130_fd_sc_hd__and3_1 _11752_ (.A(_03221_),
    .B(_03253_),
    .C(_03254_),
    .X(_03255_));
 sky130_fd_sc_hd__nand3_2 _11753_ (.A(_03221_),
    .B(_03253_),
    .C(_03254_),
    .Y(_03256_));
 sky130_fd_sc_hd__a21oi_2 _11754_ (.A1(_03253_),
    .A2(_03254_),
    .B1(_03221_),
    .Y(_03257_));
 sky130_fd_sc_hd__nand4_1 _11755_ (.A(net448),
    .B(net443),
    .C(net515),
    .D(net520),
    .Y(_03258_));
 sky130_fd_sc_hd__and2_1 _11756_ (.A(net440),
    .B(net525),
    .X(_03259_));
 sky130_fd_sc_hd__a22o_1 _11757_ (.A1(net448),
    .A2(net515),
    .B1(net520),
    .B2(net443),
    .X(_03260_));
 sky130_fd_sc_hd__nand3_1 _11758_ (.A(_03258_),
    .B(_03259_),
    .C(_03260_),
    .Y(_03261_));
 sky130_fd_sc_hd__a21bo_1 _11759_ (.A1(_03259_),
    .A2(_03260_),
    .B1_N(_03258_),
    .X(_03262_));
 sky130_fd_sc_hd__a21o_1 _11760_ (.A1(_03241_),
    .A2(_03243_),
    .B1(_03242_),
    .X(_03263_));
 sky130_fd_sc_hd__nand3_1 _11761_ (.A(_03244_),
    .B(_03262_),
    .C(_03263_),
    .Y(_03264_));
 sky130_fd_sc_hd__a21o_1 _11762_ (.A1(_03244_),
    .A2(_03263_),
    .B1(_03262_),
    .X(_03265_));
 sky130_fd_sc_hd__xnor2_2 _11763_ (.A(_03177_),
    .B(_03179_),
    .Y(_03266_));
 sky130_fd_sc_hd__nand3_2 _11764_ (.A(_03264_),
    .B(_03265_),
    .C(_03266_),
    .Y(_03267_));
 sky130_fd_sc_hd__a21bo_1 _11765_ (.A1(_03265_),
    .A2(_03266_),
    .B1_N(_03264_),
    .X(_03268_));
 sky130_fd_sc_hd__a21o_1 _11766_ (.A1(_03247_),
    .A2(_03248_),
    .B1(_03250_),
    .X(_03269_));
 sky130_fd_sc_hd__nand3_4 _11767_ (.A(_03251_),
    .B(_03268_),
    .C(_03269_),
    .Y(_03270_));
 sky130_fd_sc_hd__a21o_1 _11768_ (.A1(_03251_),
    .A2(_03269_),
    .B1(_03268_),
    .X(_03271_));
 sky130_fd_sc_hd__a21oi_1 _11769_ (.A1(_03185_),
    .A2(_03187_),
    .B1(_03186_),
    .Y(_03272_));
 sky130_fd_sc_hd__nor2_1 _11770_ (.A(_03188_),
    .B(_03272_),
    .Y(_03273_));
 sky130_fd_sc_hd__and3_1 _11771_ (.A(_03270_),
    .B(_03271_),
    .C(_03273_),
    .X(_03274_));
 sky130_fd_sc_hd__nand3_2 _11772_ (.A(_03270_),
    .B(_03271_),
    .C(_03273_),
    .Y(_03275_));
 sky130_fd_sc_hd__a211oi_4 _11773_ (.A1(_03270_),
    .A2(_03275_),
    .B1(_03255_),
    .C1(_03257_),
    .Y(_03276_));
 sky130_fd_sc_hd__o211a_2 _11774_ (.A1(_03255_),
    .A2(_03257_),
    .B1(_03270_),
    .C1(_03275_),
    .X(_03277_));
 sky130_fd_sc_hd__nor4_2 _11775_ (.A(_03206_),
    .B(_03207_),
    .C(_03276_),
    .D(_03277_),
    .Y(_03278_));
 sky130_fd_sc_hd__or4_2 _11776_ (.A(_03206_),
    .B(_03207_),
    .C(_03276_),
    .D(_03277_),
    .X(_03279_));
 sky130_fd_sc_hd__o22ai_4 _11777_ (.A1(_03206_),
    .A2(_03207_),
    .B1(_03276_),
    .B2(_03277_),
    .Y(_03280_));
 sky130_fd_sc_hd__nand4_1 _11778_ (.A(net448),
    .B(net444),
    .C(net520),
    .D(net525),
    .Y(_03281_));
 sky130_fd_sc_hd__and2_1 _11779_ (.A(net440),
    .B(net530),
    .X(_03282_));
 sky130_fd_sc_hd__a22o_1 _11780_ (.A1(net448),
    .A2(net520),
    .B1(net525),
    .B2(net443),
    .X(_03283_));
 sky130_fd_sc_hd__nand3_1 _11781_ (.A(_03281_),
    .B(_03282_),
    .C(_03283_),
    .Y(_03284_));
 sky130_fd_sc_hd__a21bo_1 _11782_ (.A1(_03282_),
    .A2(_03283_),
    .B1_N(_03281_),
    .X(_03285_));
 sky130_fd_sc_hd__a21o_1 _11783_ (.A1(_03258_),
    .A2(_03260_),
    .B1(_03259_),
    .X(_03286_));
 sky130_fd_sc_hd__nand3_1 _11784_ (.A(_03261_),
    .B(_03285_),
    .C(_03286_),
    .Y(_03287_));
 sky130_fd_sc_hd__a21o_1 _11785_ (.A1(_03261_),
    .A2(_03286_),
    .B1(_03285_),
    .X(_03288_));
 sky130_fd_sc_hd__o2bb2a_1 _11786_ (.A1_N(net426),
    .A2_N(net540),
    .B1(_03128_),
    .B2(_03129_),
    .X(_03289_));
 sky130_fd_sc_hd__nor2_1 _11787_ (.A(_03130_),
    .B(_03289_),
    .Y(_03290_));
 sky130_fd_sc_hd__nand3_2 _11788_ (.A(_03287_),
    .B(_03288_),
    .C(_03290_),
    .Y(_03291_));
 sky130_fd_sc_hd__a21bo_1 _11789_ (.A1(_03288_),
    .A2(_03290_),
    .B1_N(_03287_),
    .X(_03292_));
 sky130_fd_sc_hd__a21o_1 _11790_ (.A1(_03264_),
    .A2(_03265_),
    .B1(_03266_),
    .X(_03293_));
 sky130_fd_sc_hd__nand3_4 _11791_ (.A(_03267_),
    .B(_03292_),
    .C(_03293_),
    .Y(_03294_));
 sky130_fd_sc_hd__a21o_1 _11792_ (.A1(_03267_),
    .A2(_03293_),
    .B1(_03292_),
    .X(_03295_));
 sky130_fd_sc_hd__xnor2_2 _11793_ (.A(_03136_),
    .B(_03138_),
    .Y(_03296_));
 sky130_fd_sc_hd__and3_1 _11794_ (.A(_03294_),
    .B(_03295_),
    .C(_03296_),
    .X(_03297_));
 sky130_fd_sc_hd__nand3_2 _11795_ (.A(_03294_),
    .B(_03295_),
    .C(_03296_),
    .Y(_03298_));
 sky130_fd_sc_hd__a21oi_2 _11796_ (.A1(_03270_),
    .A2(_03271_),
    .B1(_03273_),
    .Y(_03299_));
 sky130_fd_sc_hd__a211oi_4 _11797_ (.A1(_03294_),
    .A2(_03298_),
    .B1(_03299_),
    .C1(_03274_),
    .Y(_03300_));
 sky130_fd_sc_hd__o211a_1 _11798_ (.A1(_03274_),
    .A2(_03299_),
    .B1(_03298_),
    .C1(_03294_),
    .X(_03301_));
 sky130_fd_sc_hd__xnor2_2 _11799_ (.A(_03156_),
    .B(_03158_),
    .Y(_03302_));
 sky130_fd_sc_hd__nor3_2 _11800_ (.A(_03300_),
    .B(_03301_),
    .C(_03302_),
    .Y(_03303_));
 sky130_fd_sc_hd__or3_2 _11801_ (.A(_03300_),
    .B(_03301_),
    .C(_03302_),
    .X(_03304_));
 sky130_fd_sc_hd__o211a_1 _11802_ (.A1(_03300_),
    .A2(_03303_),
    .B1(_03279_),
    .C1(_03280_),
    .X(_03305_));
 sky130_fd_sc_hd__o211ai_2 _11803_ (.A1(_03300_),
    .A2(_03303_),
    .B1(_03279_),
    .C1(_03280_),
    .Y(_03306_));
 sky130_fd_sc_hd__a211o_1 _11804_ (.A1(_03279_),
    .A2(_03280_),
    .B1(_03300_),
    .C1(_03303_),
    .X(_03307_));
 sky130_fd_sc_hd__and3_2 _11805_ (.A(_03175_),
    .B(_03306_),
    .C(_03307_),
    .X(_03308_));
 sky130_fd_sc_hd__a21oi_2 _11806_ (.A1(_03306_),
    .A2(_03307_),
    .B1(_03175_),
    .Y(_03309_));
 sky130_fd_sc_hd__nand4_1 _11807_ (.A(net449),
    .B(net444),
    .C(net525),
    .D(net530),
    .Y(_03310_));
 sky130_fd_sc_hd__and2_1 _11808_ (.A(net440),
    .B(net535),
    .X(_03311_));
 sky130_fd_sc_hd__a22o_1 _11809_ (.A1(net449),
    .A2(net525),
    .B1(net530),
    .B2(net444),
    .X(_03312_));
 sky130_fd_sc_hd__nand3_1 _11810_ (.A(_03310_),
    .B(_03311_),
    .C(_03312_),
    .Y(_03313_));
 sky130_fd_sc_hd__a21bo_1 _11811_ (.A1(_03311_),
    .A2(_03312_),
    .B1_N(_03310_),
    .X(_03314_));
 sky130_fd_sc_hd__a21o_1 _11812_ (.A1(_03281_),
    .A2(_03283_),
    .B1(_03282_),
    .X(_03315_));
 sky130_fd_sc_hd__nand3_1 _11813_ (.A(_03284_),
    .B(_03314_),
    .C(_03315_),
    .Y(_03316_));
 sky130_fd_sc_hd__a21o_1 _11814_ (.A1(_03284_),
    .A2(_03315_),
    .B1(_03314_),
    .X(_03317_));
 sky130_fd_sc_hd__xnor2_2 _11815_ (.A(_03061_),
    .B(_03063_),
    .Y(_03318_));
 sky130_fd_sc_hd__nand3_2 _11816_ (.A(_03316_),
    .B(_03317_),
    .C(_03318_),
    .Y(_03319_));
 sky130_fd_sc_hd__a21bo_1 _11817_ (.A1(_03317_),
    .A2(_03318_),
    .B1_N(_03316_),
    .X(_03320_));
 sky130_fd_sc_hd__a21o_1 _11818_ (.A1(_03287_),
    .A2(_03288_),
    .B1(_03290_),
    .X(_03321_));
 sky130_fd_sc_hd__nand3_4 _11819_ (.A(_03291_),
    .B(_03320_),
    .C(_03321_),
    .Y(_03322_));
 sky130_fd_sc_hd__a21o_1 _11820_ (.A1(_03291_),
    .A2(_03321_),
    .B1(_03320_),
    .X(_03323_));
 sky130_fd_sc_hd__xor2_2 _11821_ (.A(_03075_),
    .B(_03076_),
    .X(_03324_));
 sky130_fd_sc_hd__and3_1 _11822_ (.A(_03322_),
    .B(_03323_),
    .C(_03324_),
    .X(_03325_));
 sky130_fd_sc_hd__nand3_2 _11823_ (.A(_03322_),
    .B(_03323_),
    .C(_03324_),
    .Y(_03326_));
 sky130_fd_sc_hd__a21oi_2 _11824_ (.A1(_03294_),
    .A2(_03295_),
    .B1(_03296_),
    .Y(_03327_));
 sky130_fd_sc_hd__a211o_2 _11825_ (.A1(_03322_),
    .A2(_03326_),
    .B1(_03327_),
    .C1(_03297_),
    .X(_03328_));
 sky130_fd_sc_hd__inv_2 _11826_ (.A(_03328_),
    .Y(_03329_));
 sky130_fd_sc_hd__o211ai_4 _11827_ (.A1(_03297_),
    .A2(_03327_),
    .B1(_03326_),
    .C1(_03322_),
    .Y(_03330_));
 sky130_fd_sc_hd__a211o_1 _11828_ (.A1(_03097_),
    .A2(_03113_),
    .B1(_03112_),
    .C1(_03104_),
    .X(_03331_));
 sky130_fd_sc_hd__and4_1 _11829_ (.A(_03114_),
    .B(_03328_),
    .C(_03330_),
    .D(_03331_),
    .X(_03332_));
 sky130_fd_sc_hd__nand4_2 _11830_ (.A(_03114_),
    .B(_03328_),
    .C(_03330_),
    .D(_03331_),
    .Y(_03333_));
 sky130_fd_sc_hd__o21ai_2 _11831_ (.A1(_03300_),
    .A2(_03301_),
    .B1(_03302_),
    .Y(_03334_));
 sky130_fd_sc_hd__o211ai_4 _11832_ (.A1(_03329_),
    .A2(_03332_),
    .B1(_03334_),
    .C1(_03304_),
    .Y(_03335_));
 sky130_fd_sc_hd__and3_1 _11833_ (.A(_03097_),
    .B(_03114_),
    .C(_03126_),
    .X(_03336_));
 sky130_fd_sc_hd__nor2_1 _11834_ (.A(_03127_),
    .B(_03336_),
    .Y(_03337_));
 sky130_fd_sc_hd__a211o_1 _11835_ (.A1(_03304_),
    .A2(_03334_),
    .B1(_03332_),
    .C1(_03329_),
    .X(_03338_));
 sky130_fd_sc_hd__nand3_4 _11836_ (.A(_03335_),
    .B(_03337_),
    .C(_03338_),
    .Y(_03339_));
 sky130_fd_sc_hd__a211oi_4 _11837_ (.A1(_03335_),
    .A2(_03339_),
    .B1(_03308_),
    .C1(_03309_),
    .Y(_03340_));
 sky130_fd_sc_hd__o211a_1 _11838_ (.A1(_03308_),
    .A2(_03309_),
    .B1(_03335_),
    .C1(_03339_),
    .X(_03341_));
 sky130_fd_sc_hd__nor3b_2 _11839_ (.A(_03340_),
    .B(_03341_),
    .C_N(_03127_),
    .Y(_03342_));
 sky130_fd_sc_hd__or3b_1 _11840_ (.A(_03340_),
    .B(_03341_),
    .C_N(_03127_),
    .X(_03343_));
 sky130_fd_sc_hd__o21bai_1 _11841_ (.A1(_03340_),
    .A2(_03341_),
    .B1_N(_03127_),
    .Y(_03344_));
 sky130_fd_sc_hd__nand4_1 _11842_ (.A(net449),
    .B(net444),
    .C(net530),
    .D(net535),
    .Y(_03345_));
 sky130_fd_sc_hd__and2_1 _11843_ (.A(net440),
    .B(net540),
    .X(_03346_));
 sky130_fd_sc_hd__a22o_1 _11844_ (.A1(net449),
    .A2(net530),
    .B1(net535),
    .B2(net444),
    .X(_03347_));
 sky130_fd_sc_hd__nand3_1 _11845_ (.A(_03345_),
    .B(_03346_),
    .C(_03347_),
    .Y(_03348_));
 sky130_fd_sc_hd__a21bo_1 _11846_ (.A1(_03346_),
    .A2(_03347_),
    .B1_N(_03345_),
    .X(_03349_));
 sky130_fd_sc_hd__a21o_1 _11847_ (.A1(_03310_),
    .A2(_03312_),
    .B1(_03311_),
    .X(_03350_));
 sky130_fd_sc_hd__nand3_2 _11848_ (.A(_03313_),
    .B(_03349_),
    .C(_03350_),
    .Y(_03351_));
 sky130_fd_sc_hd__a21o_1 _11849_ (.A1(_03313_),
    .A2(_03350_),
    .B1(_03349_),
    .X(_03352_));
 sky130_fd_sc_hd__nand2_1 _11850_ (.A(net426),
    .B(net548),
    .Y(_03353_));
 sky130_fd_sc_hd__a22o_1 _11851_ (.A1(net436),
    .A2(net540),
    .B1(net544),
    .B2(net431),
    .X(_03354_));
 sky130_fd_sc_hd__a21bo_1 _11852_ (.A1(net544),
    .A2(_03059_),
    .B1_N(_03354_),
    .X(_03355_));
 sky130_fd_sc_hd__xor2_1 _11853_ (.A(_03353_),
    .B(_03355_),
    .X(_03356_));
 sky130_fd_sc_hd__nand3_1 _11854_ (.A(_03351_),
    .B(_03352_),
    .C(_03356_),
    .Y(_03357_));
 sky130_fd_sc_hd__a21bo_1 _11855_ (.A1(_03352_),
    .A2(_03356_),
    .B1_N(_03351_),
    .X(_03358_));
 sky130_fd_sc_hd__a21o_1 _11856_ (.A1(_03316_),
    .A2(_03317_),
    .B1(_03318_),
    .X(_03359_));
 sky130_fd_sc_hd__nand3_4 _11857_ (.A(_03319_),
    .B(_03358_),
    .C(_03359_),
    .Y(_03360_));
 sky130_fd_sc_hd__a21o_1 _11858_ (.A1(_03319_),
    .A2(_03359_),
    .B1(_03358_),
    .X(_03361_));
 sky130_fd_sc_hd__and4_1 _11859_ (.A(net422),
    .B(net418),
    .C(net552),
    .D(net558),
    .X(_03362_));
 sky130_fd_sc_hd__nand2_1 _11860_ (.A(net413),
    .B(net565),
    .Y(_03363_));
 sky130_fd_sc_hd__a22o_1 _11861_ (.A1(net422),
    .A2(net552),
    .B1(net558),
    .B2(net418),
    .X(_03364_));
 sky130_fd_sc_hd__and2b_1 _11862_ (.A_N(_03362_),
    .B(_03364_),
    .X(_03365_));
 sky130_fd_sc_hd__a31o_1 _11863_ (.A1(net413),
    .A2(net565),
    .A3(_03364_),
    .B1(_03362_),
    .X(_03366_));
 sky130_fd_sc_hd__a32o_1 _11864_ (.A1(net427),
    .A2(net548),
    .A3(_03354_),
    .B1(_03059_),
    .B2(net544),
    .X(_03367_));
 sky130_fd_sc_hd__xnor2_2 _11865_ (.A(_03072_),
    .B(_03074_),
    .Y(_03368_));
 sky130_fd_sc_hd__nand2_1 _11866_ (.A(_03367_),
    .B(_03368_),
    .Y(_03369_));
 sky130_fd_sc_hd__xor2_2 _11867_ (.A(_03367_),
    .B(_03368_),
    .X(_03370_));
 sky130_fd_sc_hd__nand2_1 _11868_ (.A(_03366_),
    .B(_03370_),
    .Y(_03371_));
 sky130_fd_sc_hd__xor2_2 _11869_ (.A(_03366_),
    .B(_03370_),
    .X(_03372_));
 sky130_fd_sc_hd__nand3_4 _11870_ (.A(_03360_),
    .B(_03361_),
    .C(_03372_),
    .Y(_03373_));
 sky130_fd_sc_hd__a21oi_2 _11871_ (.A1(_03322_),
    .A2(_03323_),
    .B1(_03324_),
    .Y(_03374_));
 sky130_fd_sc_hd__a211oi_4 _11872_ (.A1(_03360_),
    .A2(_03373_),
    .B1(_03374_),
    .C1(_03325_),
    .Y(_03375_));
 sky130_fd_sc_hd__o211a_1 _11873_ (.A1(_03325_),
    .A2(_03374_),
    .B1(_03373_),
    .C1(_03360_),
    .X(_03376_));
 sky130_fd_sc_hd__xnor2_1 _11874_ (.A(_03100_),
    .B(_03102_),
    .Y(_03377_));
 sky130_fd_sc_hd__and4_1 _11875_ (.A(net408),
    .B(net404),
    .C(net567),
    .D(net572),
    .X(_03378_));
 sky130_fd_sc_hd__inv_2 _11876_ (.A(_03378_),
    .Y(_03379_));
 sky130_fd_sc_hd__a22o_1 _11877_ (.A1(net408),
    .A2(net567),
    .B1(net572),
    .B2(net404),
    .X(_03380_));
 sky130_fd_sc_hd__and4b_1 _11878_ (.A_N(_03378_),
    .B(_03380_),
    .C(net400),
    .D(net577),
    .X(_03381_));
 sky130_fd_sc_hd__or2_1 _11879_ (.A(_03378_),
    .B(_03381_),
    .X(_03382_));
 sky130_fd_sc_hd__and2_1 _11880_ (.A(_03377_),
    .B(_03382_),
    .X(_03383_));
 sky130_fd_sc_hd__xor2_1 _11881_ (.A(_03377_),
    .B(_03382_),
    .X(_03384_));
 sky130_fd_sc_hd__a22o_1 _11882_ (.A1(net396),
    .A2(net577),
    .B1(net581),
    .B2(net390),
    .X(_03385_));
 sky130_fd_sc_hd__inv_2 _11883_ (.A(_03385_),
    .Y(_03386_));
 sky130_fd_sc_hd__and4_1 _11884_ (.A(net396),
    .B(net390),
    .C(net577),
    .D(net581),
    .X(_03387_));
 sky130_fd_sc_hd__nor2_1 _11885_ (.A(_03386_),
    .B(_03387_),
    .Y(_03388_));
 sky130_fd_sc_hd__and2_1 _11886_ (.A(_03384_),
    .B(_03388_),
    .X(_03389_));
 sky130_fd_sc_hd__xnor2_1 _11887_ (.A(_03105_),
    .B(_03111_),
    .Y(_03390_));
 sky130_fd_sc_hd__a21o_1 _11888_ (.A1(_03369_),
    .A2(_03371_),
    .B1(_03390_),
    .X(_03391_));
 sky130_fd_sc_hd__nand3_1 _11889_ (.A(_03369_),
    .B(_03371_),
    .C(_03390_),
    .Y(_03392_));
 sky130_fd_sc_hd__o211ai_2 _11890_ (.A1(_03383_),
    .A2(_03389_),
    .B1(_03391_),
    .C1(_03392_),
    .Y(_03393_));
 sky130_fd_sc_hd__a211o_1 _11891_ (.A1(_03391_),
    .A2(_03392_),
    .B1(_03383_),
    .C1(_03389_),
    .X(_03394_));
 sky130_fd_sc_hd__and4bb_2 _11892_ (.A_N(_03375_),
    .B_N(_03376_),
    .C(_03393_),
    .D(_03394_),
    .X(_03395_));
 sky130_fd_sc_hd__a22o_1 _11893_ (.A1(_03328_),
    .A2(_03330_),
    .B1(_03331_),
    .B2(_03114_),
    .X(_03396_));
 sky130_fd_sc_hd__o211a_1 _11894_ (.A1(_03375_),
    .A2(_03395_),
    .B1(_03396_),
    .C1(_03333_),
    .X(_03397_));
 sky130_fd_sc_hd__o211ai_1 _11895_ (.A1(_03375_),
    .A2(_03395_),
    .B1(_03396_),
    .C1(_03333_),
    .Y(_03398_));
 sky130_fd_sc_hd__a211o_1 _11896_ (.A1(_03333_),
    .A2(_03396_),
    .B1(_03395_),
    .C1(_03375_),
    .X(_03399_));
 sky130_fd_sc_hd__xnor2_1 _11897_ (.A(_03115_),
    .B(_03116_),
    .Y(_03400_));
 sky130_fd_sc_hd__a21oi_1 _11898_ (.A1(_03391_),
    .A2(_03393_),
    .B1(_03400_),
    .Y(_03401_));
 sky130_fd_sc_hd__and3_1 _11899_ (.A(_03391_),
    .B(_03393_),
    .C(_03400_),
    .X(_03402_));
 sky130_fd_sc_hd__nor2_1 _11900_ (.A(_03401_),
    .B(_03402_),
    .Y(_03403_));
 sky130_fd_sc_hd__and3_2 _11901_ (.A(_03398_),
    .B(_03399_),
    .C(_03403_),
    .X(_03404_));
 sky130_fd_sc_hd__a21o_1 _11902_ (.A1(_03335_),
    .A2(_03338_),
    .B1(_03337_),
    .X(_03405_));
 sky130_fd_sc_hd__o211a_1 _11903_ (.A1(_03397_),
    .A2(_03404_),
    .B1(_03405_),
    .C1(_03339_),
    .X(_03406_));
 sky130_fd_sc_hd__a211oi_2 _11904_ (.A1(_03339_),
    .A2(_03405_),
    .B1(_03404_),
    .C1(_03397_),
    .Y(_03407_));
 sky130_fd_sc_hd__nor3b_2 _11905_ (.A(_03406_),
    .B(_03407_),
    .C_N(_03401_),
    .Y(_03408_));
 sky130_fd_sc_hd__o211a_1 _11906_ (.A1(_03406_),
    .A2(_03408_),
    .B1(_03343_),
    .C1(_03344_),
    .X(_03409_));
 sky130_fd_sc_hd__inv_2 _11907_ (.A(_03409_),
    .Y(_03410_));
 sky130_fd_sc_hd__a211o_1 _11908_ (.A1(_03343_),
    .A2(_03344_),
    .B1(_03406_),
    .C1(_03408_),
    .X(_03411_));
 sky130_fd_sc_hd__nand2b_2 _11909_ (.A_N(_03409_),
    .B(_03411_),
    .Y(_03412_));
 sky130_fd_sc_hd__o21ba_1 _11910_ (.A1(_03406_),
    .A2(_03407_),
    .B1_N(_03401_),
    .X(_03413_));
 sky130_fd_sc_hd__nand4_1 _11911_ (.A(net449),
    .B(net444),
    .C(net535),
    .D(net540),
    .Y(_03414_));
 sky130_fd_sc_hd__and2_1 _11912_ (.A(net440),
    .B(net544),
    .X(_03415_));
 sky130_fd_sc_hd__a22o_1 _11913_ (.A1(net448),
    .A2(net535),
    .B1(net540),
    .B2(net443),
    .X(_03416_));
 sky130_fd_sc_hd__nand3_1 _11914_ (.A(_03414_),
    .B(_03415_),
    .C(_03416_),
    .Y(_03417_));
 sky130_fd_sc_hd__a21bo_1 _11915_ (.A1(_03415_),
    .A2(_03416_),
    .B1_N(_03414_),
    .X(_03418_));
 sky130_fd_sc_hd__a21o_1 _11916_ (.A1(_03345_),
    .A2(_03347_),
    .B1(_03346_),
    .X(_03419_));
 sky130_fd_sc_hd__nand3_1 _11917_ (.A(_03348_),
    .B(_03418_),
    .C(_03419_),
    .Y(_03420_));
 sky130_fd_sc_hd__a21o_1 _11918_ (.A1(_03348_),
    .A2(_03419_),
    .B1(_03418_),
    .X(_03421_));
 sky130_fd_sc_hd__nand2_1 _11919_ (.A(net427),
    .B(net552),
    .Y(_03422_));
 sky130_fd_sc_hd__a22oi_2 _11920_ (.A1(net435),
    .A2(net544),
    .B1(net549),
    .B2(net430),
    .Y(_03423_));
 sky130_fd_sc_hd__and4_1 _11921_ (.A(net435),
    .B(net430),
    .C(net544),
    .D(net549),
    .X(_03424_));
 sky130_fd_sc_hd__nor2_1 _11922_ (.A(_03423_),
    .B(_03424_),
    .Y(_03425_));
 sky130_fd_sc_hd__xnor2_1 _11923_ (.A(_03422_),
    .B(_03425_),
    .Y(_03426_));
 sky130_fd_sc_hd__nand3_1 _11924_ (.A(_03420_),
    .B(_03421_),
    .C(_03426_),
    .Y(_03427_));
 sky130_fd_sc_hd__a21bo_1 _11925_ (.A1(_03421_),
    .A2(_03426_),
    .B1_N(_03420_),
    .X(_03428_));
 sky130_fd_sc_hd__a21o_1 _11926_ (.A1(_03351_),
    .A2(_03352_),
    .B1(_03356_),
    .X(_03429_));
 sky130_fd_sc_hd__and3_1 _11927_ (.A(_03357_),
    .B(_03428_),
    .C(_03429_),
    .X(_03430_));
 sky130_fd_sc_hd__nand3_1 _11928_ (.A(_03357_),
    .B(_03428_),
    .C(_03429_),
    .Y(_03431_));
 sky130_fd_sc_hd__a21o_1 _11929_ (.A1(_03357_),
    .A2(_03429_),
    .B1(_03428_),
    .X(_03432_));
 sky130_fd_sc_hd__and4_1 _11930_ (.A(net422),
    .B(net418),
    .C(net558),
    .D(net565),
    .X(_03433_));
 sky130_fd_sc_hd__nand2_1 _11931_ (.A(net413),
    .B(net570),
    .Y(_03434_));
 sky130_fd_sc_hd__a22o_1 _11932_ (.A1(net422),
    .A2(net558),
    .B1(net561),
    .B2(net418),
    .X(_03435_));
 sky130_fd_sc_hd__and2b_1 _11933_ (.A_N(_03433_),
    .B(_03435_),
    .X(_03436_));
 sky130_fd_sc_hd__a31o_1 _11934_ (.A1(net414),
    .A2(net566),
    .A3(_03435_),
    .B1(_03433_),
    .X(_03437_));
 sky130_fd_sc_hd__o21ba_1 _11935_ (.A1(_03422_),
    .A2(_03423_),
    .B1_N(_03424_),
    .X(_03438_));
 sky130_fd_sc_hd__xnor2_1 _11936_ (.A(_03363_),
    .B(_03365_),
    .Y(_03439_));
 sky130_fd_sc_hd__nand2b_1 _11937_ (.A_N(_03438_),
    .B(_03439_),
    .Y(_03440_));
 sky130_fd_sc_hd__xnor2_1 _11938_ (.A(_03438_),
    .B(_03439_),
    .Y(_03441_));
 sky130_fd_sc_hd__nand2_1 _11939_ (.A(_03437_),
    .B(_03441_),
    .Y(_03442_));
 sky130_fd_sc_hd__xor2_1 _11940_ (.A(_03437_),
    .B(_03441_),
    .X(_03443_));
 sky130_fd_sc_hd__and3_2 _11941_ (.A(_03431_),
    .B(_03432_),
    .C(_03443_),
    .X(_03444_));
 sky130_fd_sc_hd__a21o_1 _11942_ (.A1(_03360_),
    .A2(_03361_),
    .B1(_03372_),
    .X(_03445_));
 sky130_fd_sc_hd__o211a_1 _11943_ (.A1(_03430_),
    .A2(_03444_),
    .B1(_03445_),
    .C1(_03373_),
    .X(_03446_));
 sky130_fd_sc_hd__o211ai_2 _11944_ (.A1(_03430_),
    .A2(_03444_),
    .B1(_03445_),
    .C1(_03373_),
    .Y(_03447_));
 sky130_fd_sc_hd__a211oi_1 _11945_ (.A1(_03373_),
    .A2(_03445_),
    .B1(_03444_),
    .C1(_03430_),
    .Y(_03448_));
 sky130_fd_sc_hd__nor2_1 _11946_ (.A(_03446_),
    .B(_03448_),
    .Y(_03449_));
 sky130_fd_sc_hd__a22oi_1 _11947_ (.A1(net400),
    .A2(net577),
    .B1(_03379_),
    .B2(_03380_),
    .Y(_03450_));
 sky130_fd_sc_hd__nor2_1 _11948_ (.A(_03381_),
    .B(_03450_),
    .Y(_03451_));
 sky130_fd_sc_hd__and4_1 _11949_ (.A(net408),
    .B(net404),
    .C(net572),
    .D(net577),
    .X(_03452_));
 sky130_fd_sc_hd__inv_2 _11950_ (.A(_03452_),
    .Y(_03453_));
 sky130_fd_sc_hd__a22o_1 _11951_ (.A1(net408),
    .A2(net572),
    .B1(net577),
    .B2(net404),
    .X(_03454_));
 sky130_fd_sc_hd__and4_1 _11952_ (.A(net400),
    .B(net581),
    .C(_03453_),
    .D(_03454_),
    .X(_03455_));
 sky130_fd_sc_hd__or2_1 _11953_ (.A(_03452_),
    .B(_03455_),
    .X(_03456_));
 sky130_fd_sc_hd__nand2_1 _11954_ (.A(_03451_),
    .B(_03456_),
    .Y(_03457_));
 sky130_fd_sc_hd__nand2_1 _11955_ (.A(net396),
    .B(net581),
    .Y(_03458_));
 sky130_fd_sc_hd__xor2_1 _11956_ (.A(_03451_),
    .B(_03456_),
    .X(_03459_));
 sky130_fd_sc_hd__nand2b_1 _11957_ (.A_N(_03458_),
    .B(_03459_),
    .Y(_03460_));
 sky130_fd_sc_hd__xnor2_1 _11958_ (.A(_03384_),
    .B(_03388_),
    .Y(_03461_));
 sky130_fd_sc_hd__a21oi_2 _11959_ (.A1(_03440_),
    .A2(_03442_),
    .B1(_03461_),
    .Y(_03462_));
 sky130_fd_sc_hd__and3_1 _11960_ (.A(_03440_),
    .B(_03442_),
    .C(_03461_),
    .X(_03463_));
 sky130_fd_sc_hd__a211oi_2 _11961_ (.A1(_03457_),
    .A2(_03460_),
    .B1(_03462_),
    .C1(_03463_),
    .Y(_03464_));
 sky130_fd_sc_hd__o211a_1 _11962_ (.A1(_03462_),
    .A2(_03463_),
    .B1(_03457_),
    .C1(_03460_),
    .X(_03465_));
 sky130_fd_sc_hd__nor2_1 _11963_ (.A(_03464_),
    .B(_03465_),
    .Y(_03466_));
 sky130_fd_sc_hd__or4_2 _11964_ (.A(_03446_),
    .B(_03448_),
    .C(_03464_),
    .D(_03465_),
    .X(_03467_));
 sky130_fd_sc_hd__a2bb2oi_1 _11965_ (.A1_N(_03375_),
    .A2_N(_03376_),
    .B1(_03393_),
    .B2(_03394_),
    .Y(_03468_));
 sky130_fd_sc_hd__a211o_2 _11966_ (.A1(_03447_),
    .A2(_03467_),
    .B1(_03468_),
    .C1(_03395_),
    .X(_03469_));
 sky130_fd_sc_hd__o211ai_2 _11967_ (.A1(_03395_),
    .A2(_03468_),
    .B1(_03467_),
    .C1(_03447_),
    .Y(_03470_));
 sky130_fd_sc_hd__o21ai_2 _11968_ (.A1(_03462_),
    .A2(_03464_),
    .B1(_03387_),
    .Y(_03471_));
 sky130_fd_sc_hd__or3_1 _11969_ (.A(_03387_),
    .B(_03462_),
    .C(_03464_),
    .X(_03472_));
 sky130_fd_sc_hd__and2_1 _11970_ (.A(_03471_),
    .B(_03472_),
    .X(_03473_));
 sky130_fd_sc_hd__nand3_2 _11971_ (.A(_03469_),
    .B(_03470_),
    .C(_03473_),
    .Y(_03474_));
 sky130_fd_sc_hd__a21oi_1 _11972_ (.A1(_03398_),
    .A2(_03399_),
    .B1(_03403_),
    .Y(_03475_));
 sky130_fd_sc_hd__a211o_1 _11973_ (.A1(_03469_),
    .A2(_03474_),
    .B1(_03475_),
    .C1(_03404_),
    .X(_03476_));
 sky130_fd_sc_hd__o211a_1 _11974_ (.A1(_03404_),
    .A2(_03475_),
    .B1(_03474_),
    .C1(_03469_),
    .X(_03477_));
 sky130_fd_sc_hd__o211ai_1 _11975_ (.A1(_03404_),
    .A2(_03475_),
    .B1(_03474_),
    .C1(_03469_),
    .Y(_03478_));
 sky130_fd_sc_hd__and2_1 _11976_ (.A(_03476_),
    .B(_03478_),
    .X(_03479_));
 sky130_fd_sc_hd__or3b_1 _11977_ (.A(_03477_),
    .B(_03471_),
    .C_N(_03476_),
    .X(_03480_));
 sky130_fd_sc_hd__a211oi_2 _11978_ (.A1(_03476_),
    .A2(_03480_),
    .B1(_03408_),
    .C1(_03413_),
    .Y(_03481_));
 sky130_fd_sc_hd__xnor2_1 _11979_ (.A(_03471_),
    .B(_03479_),
    .Y(_03482_));
 sky130_fd_sc_hd__and2b_1 _11980_ (.A_N(_03481_),
    .B(_03482_),
    .X(_03483_));
 sky130_fd_sc_hd__a21o_1 _11981_ (.A1(_03469_),
    .A2(_03470_),
    .B1(_03473_),
    .X(_03484_));
 sky130_fd_sc_hd__and2_1 _11982_ (.A(_03474_),
    .B(_03484_),
    .X(_03485_));
 sky130_fd_sc_hd__nand4_1 _11983_ (.A(net448),
    .B(net443),
    .C(net540),
    .D(net544),
    .Y(_03486_));
 sky130_fd_sc_hd__and2_1 _11984_ (.A(net440),
    .B(net549),
    .X(_03487_));
 sky130_fd_sc_hd__a22o_1 _11985_ (.A1(net449),
    .A2(net540),
    .B1(net544),
    .B2(net443),
    .X(_03488_));
 sky130_fd_sc_hd__nand3_1 _11986_ (.A(_03486_),
    .B(_03487_),
    .C(_03488_),
    .Y(_03489_));
 sky130_fd_sc_hd__a21bo_1 _11987_ (.A1(_03487_),
    .A2(_03488_),
    .B1_N(_03486_),
    .X(_03490_));
 sky130_fd_sc_hd__a21o_1 _11988_ (.A1(_03414_),
    .A2(_03416_),
    .B1(_03415_),
    .X(_03491_));
 sky130_fd_sc_hd__nand3_1 _11989_ (.A(_03417_),
    .B(_03490_),
    .C(_03491_),
    .Y(_03492_));
 sky130_fd_sc_hd__a22oi_2 _11990_ (.A1(net435),
    .A2(net549),
    .B1(net553),
    .B2(net430),
    .Y(_03493_));
 sky130_fd_sc_hd__and4_1 _11991_ (.A(net435),
    .B(net430),
    .C(net549),
    .D(net553),
    .X(_03494_));
 sky130_fd_sc_hd__nor2_1 _11992_ (.A(_03493_),
    .B(_03494_),
    .Y(_03495_));
 sky130_fd_sc_hd__nand2_1 _11993_ (.A(net427),
    .B(net557),
    .Y(_03496_));
 sky130_fd_sc_hd__xnor2_1 _11994_ (.A(_03495_),
    .B(_03496_),
    .Y(_03497_));
 sky130_fd_sc_hd__a21o_1 _11995_ (.A1(_03417_),
    .A2(_03491_),
    .B1(_03490_),
    .X(_03498_));
 sky130_fd_sc_hd__nand3_1 _11996_ (.A(_03492_),
    .B(_03497_),
    .C(_03498_),
    .Y(_03499_));
 sky130_fd_sc_hd__a21bo_1 _11997_ (.A1(_03497_),
    .A2(_03498_),
    .B1_N(_03492_),
    .X(_03500_));
 sky130_fd_sc_hd__a21o_1 _11998_ (.A1(_03420_),
    .A2(_03421_),
    .B1(_03426_),
    .X(_03501_));
 sky130_fd_sc_hd__nand3_2 _11999_ (.A(_03427_),
    .B(_03500_),
    .C(_03501_),
    .Y(_03502_));
 sky130_fd_sc_hd__o21ba_1 _12000_ (.A1(_03493_),
    .A2(_03496_),
    .B1_N(_03494_),
    .X(_03503_));
 sky130_fd_sc_hd__xnor2_1 _12001_ (.A(_03434_),
    .B(_03436_),
    .Y(_03504_));
 sky130_fd_sc_hd__and2b_1 _12002_ (.A_N(_03503_),
    .B(_03504_),
    .X(_03505_));
 sky130_fd_sc_hd__xnor2_1 _12003_ (.A(_03503_),
    .B(_03504_),
    .Y(_03506_));
 sky130_fd_sc_hd__and4_1 _12004_ (.A(net422),
    .B(net417),
    .C(net561),
    .D(net570),
    .X(_03507_));
 sky130_fd_sc_hd__nand2_1 _12005_ (.A(net414),
    .B(net571),
    .Y(_03508_));
 sky130_fd_sc_hd__a22o_1 _12006_ (.A1(net422),
    .A2(net561),
    .B1(net570),
    .B2(net418),
    .X(_03509_));
 sky130_fd_sc_hd__and2b_1 _12007_ (.A_N(_03507_),
    .B(_03509_),
    .X(_03510_));
 sky130_fd_sc_hd__a31o_1 _12008_ (.A1(net414),
    .A2(net575),
    .A3(_03509_),
    .B1(_03507_),
    .X(_03511_));
 sky130_fd_sc_hd__xor2_1 _12009_ (.A(_03506_),
    .B(_03511_),
    .X(_03512_));
 sky130_fd_sc_hd__a21o_1 _12010_ (.A1(_03427_),
    .A2(_03501_),
    .B1(_03500_),
    .X(_03513_));
 sky130_fd_sc_hd__nand3_2 _12011_ (.A(_03502_),
    .B(_03512_),
    .C(_03513_),
    .Y(_03514_));
 sky130_fd_sc_hd__a21oi_1 _12012_ (.A1(_03431_),
    .A2(_03432_),
    .B1(_03443_),
    .Y(_03515_));
 sky130_fd_sc_hd__a211o_1 _12013_ (.A1(_03502_),
    .A2(_03514_),
    .B1(_03515_),
    .C1(_03444_),
    .X(_03516_));
 sky130_fd_sc_hd__a21oi_1 _12014_ (.A1(_03506_),
    .A2(_03511_),
    .B1(_03505_),
    .Y(_03517_));
 sky130_fd_sc_hd__xnor2_1 _12015_ (.A(_03458_),
    .B(_03459_),
    .Y(_03518_));
 sky130_fd_sc_hd__nand2b_1 _12016_ (.A_N(_03517_),
    .B(_03518_),
    .Y(_03519_));
 sky130_fd_sc_hd__xnor2_1 _12017_ (.A(_03517_),
    .B(_03518_),
    .Y(_03520_));
 sky130_fd_sc_hd__a22oi_1 _12018_ (.A1(net400),
    .A2(net581),
    .B1(_03453_),
    .B2(_03454_),
    .Y(_03521_));
 sky130_fd_sc_hd__nor2_1 _12019_ (.A(_03455_),
    .B(_03521_),
    .Y(_03522_));
 sky130_fd_sc_hd__and4_1 _12020_ (.A(net408),
    .B(net404),
    .C(net577),
    .D(net581),
    .X(_03523_));
 sky130_fd_sc_hd__and2_1 _12021_ (.A(_03522_),
    .B(_03523_),
    .X(_03524_));
 sky130_fd_sc_hd__nand2_1 _12022_ (.A(_03520_),
    .B(_03524_),
    .Y(_03525_));
 sky130_fd_sc_hd__xnor2_1 _12023_ (.A(_03520_),
    .B(_03524_),
    .Y(_03526_));
 sky130_fd_sc_hd__o211ai_1 _12024_ (.A1(_03444_),
    .A2(_03515_),
    .B1(_03514_),
    .C1(_03502_),
    .Y(_03527_));
 sky130_fd_sc_hd__nand2_1 _12025_ (.A(_03516_),
    .B(_03527_),
    .Y(_03528_));
 sky130_fd_sc_hd__or2_1 _12026_ (.A(_03526_),
    .B(_03528_),
    .X(_03529_));
 sky130_fd_sc_hd__xnor2_1 _12027_ (.A(_03449_),
    .B(_03466_),
    .Y(_03530_));
 sky130_fd_sc_hd__a21oi_2 _12028_ (.A1(_03516_),
    .A2(_03529_),
    .B1(_03530_),
    .Y(_03531_));
 sky130_fd_sc_hd__and3_1 _12029_ (.A(_03516_),
    .B(_03529_),
    .C(_03530_),
    .X(_03532_));
 sky130_fd_sc_hd__or2_1 _12030_ (.A(_03531_),
    .B(_03532_),
    .X(_03533_));
 sky130_fd_sc_hd__a21oi_2 _12031_ (.A1(_03519_),
    .A2(_03525_),
    .B1(_03533_),
    .Y(_03534_));
 sky130_fd_sc_hd__o21a_1 _12032_ (.A1(_03531_),
    .A2(_03534_),
    .B1(_03485_),
    .X(_03535_));
 sky130_fd_sc_hd__o211ai_2 _12033_ (.A1(_03408_),
    .A2(_03413_),
    .B1(_03476_),
    .C1(_03480_),
    .Y(_03536_));
 sky130_fd_sc_hd__a31o_1 _12034_ (.A1(_03482_),
    .A2(_03535_),
    .A3(_03536_),
    .B1(_03481_),
    .X(_03537_));
 sky130_fd_sc_hd__xnor2_4 _12035_ (.A(_03412_),
    .B(_03537_),
    .Y(_03538_));
 sky130_fd_sc_hd__and3_1 _12036_ (.A(_03519_),
    .B(_03525_),
    .C(_03533_),
    .X(_03539_));
 sky130_fd_sc_hd__nand4_1 _12037_ (.A(net448),
    .B(net443),
    .C(net544),
    .D(net549),
    .Y(_03540_));
 sky130_fd_sc_hd__and2_1 _12038_ (.A(net440),
    .B(net553),
    .X(_03541_));
 sky130_fd_sc_hd__a22o_1 _12039_ (.A1(net449),
    .A2(net544),
    .B1(net549),
    .B2(net444),
    .X(_03542_));
 sky130_fd_sc_hd__nand3_1 _12040_ (.A(_03540_),
    .B(_03541_),
    .C(_03542_),
    .Y(_03543_));
 sky130_fd_sc_hd__a21bo_1 _12041_ (.A1(_03541_),
    .A2(_03542_),
    .B1_N(_03540_),
    .X(_03544_));
 sky130_fd_sc_hd__a21o_1 _12042_ (.A1(_03486_),
    .A2(_03488_),
    .B1(_03487_),
    .X(_03545_));
 sky130_fd_sc_hd__nand3_1 _12043_ (.A(_03489_),
    .B(_03544_),
    .C(_03545_),
    .Y(_03546_));
 sky130_fd_sc_hd__and4_1 _12044_ (.A(net435),
    .B(net430),
    .C(net553),
    .D(net557),
    .X(_03547_));
 sky130_fd_sc_hd__a22o_1 _12045_ (.A1(net435),
    .A2(net553),
    .B1(net557),
    .B2(net430),
    .X(_03548_));
 sky130_fd_sc_hd__and2b_1 _12046_ (.A_N(_03547_),
    .B(_03548_),
    .X(_03549_));
 sky130_fd_sc_hd__nand2_1 _12047_ (.A(net427),
    .B(net561),
    .Y(_03550_));
 sky130_fd_sc_hd__xnor2_1 _12048_ (.A(_03549_),
    .B(_03550_),
    .Y(_03551_));
 sky130_fd_sc_hd__a21o_1 _12049_ (.A1(_03489_),
    .A2(_03545_),
    .B1(_03544_),
    .X(_03552_));
 sky130_fd_sc_hd__nand3_1 _12050_ (.A(_03546_),
    .B(_03551_),
    .C(_03552_),
    .Y(_03553_));
 sky130_fd_sc_hd__a21bo_1 _12051_ (.A1(_03551_),
    .A2(_03552_),
    .B1_N(_03546_),
    .X(_03554_));
 sky130_fd_sc_hd__a21o_1 _12052_ (.A1(_03492_),
    .A2(_03498_),
    .B1(_03497_),
    .X(_03555_));
 sky130_fd_sc_hd__and3_1 _12053_ (.A(_03499_),
    .B(_03554_),
    .C(_03555_),
    .X(_03556_));
 sky130_fd_sc_hd__a31o_1 _12054_ (.A1(net427),
    .A2(net561),
    .A3(_03548_),
    .B1(_03547_),
    .X(_03557_));
 sky130_fd_sc_hd__xnor2_1 _12055_ (.A(_03508_),
    .B(_03510_),
    .Y(_03558_));
 sky130_fd_sc_hd__and2_1 _12056_ (.A(_03557_),
    .B(_03558_),
    .X(_03559_));
 sky130_fd_sc_hd__xor2_1 _12057_ (.A(_03557_),
    .B(_03558_),
    .X(_03560_));
 sky130_fd_sc_hd__and4_1 _12058_ (.A(net421),
    .B(net417),
    .C(net566),
    .D(net571),
    .X(_03561_));
 sky130_fd_sc_hd__nand2_1 _12059_ (.A(net413),
    .B(net576),
    .Y(_03562_));
 sky130_fd_sc_hd__a22o_1 _12060_ (.A1(net421),
    .A2(net566),
    .B1(net571),
    .B2(net417),
    .X(_03563_));
 sky130_fd_sc_hd__and2b_1 _12061_ (.A_N(_03561_),
    .B(_03563_),
    .X(_03564_));
 sky130_fd_sc_hd__a31o_1 _12062_ (.A1(net413),
    .A2(net576),
    .A3(_03563_),
    .B1(_03561_),
    .X(_03565_));
 sky130_fd_sc_hd__xnor2_1 _12063_ (.A(_03560_),
    .B(_03565_),
    .Y(_03566_));
 sky130_fd_sc_hd__a21oi_1 _12064_ (.A1(_03499_),
    .A2(_03555_),
    .B1(_03554_),
    .Y(_03567_));
 sky130_fd_sc_hd__nor3_1 _12065_ (.A(_03556_),
    .B(_03566_),
    .C(_03567_),
    .Y(_03568_));
 sky130_fd_sc_hd__or3_1 _12066_ (.A(_03556_),
    .B(_03566_),
    .C(_03567_),
    .X(_03569_));
 sky130_fd_sc_hd__a21o_1 _12067_ (.A1(_03502_),
    .A2(_03513_),
    .B1(_03512_),
    .X(_03570_));
 sky130_fd_sc_hd__o211ai_2 _12068_ (.A1(_03556_),
    .A2(_03568_),
    .B1(_03570_),
    .C1(_03514_),
    .Y(_03571_));
 sky130_fd_sc_hd__a21o_1 _12069_ (.A1(_03560_),
    .A2(_03565_),
    .B1(_03559_),
    .X(_03572_));
 sky130_fd_sc_hd__nor2_1 _12070_ (.A(_03522_),
    .B(_03523_),
    .Y(_03573_));
 sky130_fd_sc_hd__or2_1 _12071_ (.A(_03524_),
    .B(_03573_),
    .X(_03574_));
 sky130_fd_sc_hd__and2b_1 _12072_ (.A_N(_03574_),
    .B(_03572_),
    .X(_03575_));
 sky130_fd_sc_hd__xnor2_1 _12073_ (.A(_03572_),
    .B(_03574_),
    .Y(_03576_));
 sky130_fd_sc_hd__a211o_1 _12074_ (.A1(_03514_),
    .A2(_03570_),
    .B1(_03568_),
    .C1(_03556_),
    .X(_03577_));
 sky130_fd_sc_hd__nand3_1 _12075_ (.A(_03571_),
    .B(_03576_),
    .C(_03577_),
    .Y(_03578_));
 sky130_fd_sc_hd__nand2_1 _12076_ (.A(_03571_),
    .B(_03578_),
    .Y(_03579_));
 sky130_fd_sc_hd__xor2_1 _12077_ (.A(_03526_),
    .B(_03528_),
    .X(_03580_));
 sky130_fd_sc_hd__nand2_1 _12078_ (.A(_03579_),
    .B(_03580_),
    .Y(_03581_));
 sky130_fd_sc_hd__xnor2_1 _12079_ (.A(_03579_),
    .B(_03580_),
    .Y(_03582_));
 sky130_fd_sc_hd__or3b_1 _12080_ (.A(_03574_),
    .B(_03582_),
    .C_N(_03572_),
    .X(_03583_));
 sky130_fd_sc_hd__a211o_1 _12081_ (.A1(_03581_),
    .A2(_03583_),
    .B1(_03534_),
    .C1(_03539_),
    .X(_03584_));
 sky130_fd_sc_hd__o211a_1 _12082_ (.A1(_03534_),
    .A2(_03539_),
    .B1(_03581_),
    .C1(_03583_),
    .X(_03585_));
 sky130_fd_sc_hd__xor2_1 _12083_ (.A(_03575_),
    .B(_03582_),
    .X(_03586_));
 sky130_fd_sc_hd__a21o_1 _12084_ (.A1(_03571_),
    .A2(_03577_),
    .B1(_03576_),
    .X(_03587_));
 sky130_fd_sc_hd__o21ai_1 _12085_ (.A1(_03556_),
    .A2(_03567_),
    .B1(_03566_),
    .Y(_03588_));
 sky130_fd_sc_hd__a21o_1 _12086_ (.A1(_03546_),
    .A2(_03552_),
    .B1(_03551_),
    .X(_03589_));
 sky130_fd_sc_hd__a21o_1 _12087_ (.A1(_03540_),
    .A2(_03542_),
    .B1(_03541_),
    .X(_03590_));
 sky130_fd_sc_hd__nand4_2 _12088_ (.A(net448),
    .B(net443),
    .C(net549),
    .D(net553),
    .Y(_03591_));
 sky130_fd_sc_hd__and2_1 _12089_ (.A(net440),
    .B(net557),
    .X(_03592_));
 sky130_fd_sc_hd__a22o_1 _12090_ (.A1(net448),
    .A2(net549),
    .B1(net553),
    .B2(net443),
    .X(_03593_));
 sky130_fd_sc_hd__nand3_1 _12091_ (.A(_03591_),
    .B(_03592_),
    .C(_03593_),
    .Y(_03594_));
 sky130_fd_sc_hd__a21bo_1 _12092_ (.A1(_03592_),
    .A2(_03593_),
    .B1_N(_03591_),
    .X(_03595_));
 sky130_fd_sc_hd__nand3_1 _12093_ (.A(_03543_),
    .B(_03590_),
    .C(_03595_),
    .Y(_03596_));
 sky130_fd_sc_hd__and4_1 _12094_ (.A(net435),
    .B(net430),
    .C(net557),
    .D(net561),
    .X(_03597_));
 sky130_fd_sc_hd__a22o_1 _12095_ (.A1(net435),
    .A2(net557),
    .B1(net561),
    .B2(net430),
    .X(_03598_));
 sky130_fd_sc_hd__and2b_1 _12096_ (.A_N(_03597_),
    .B(_03598_),
    .X(_03599_));
 sky130_fd_sc_hd__nand2_1 _12097_ (.A(net426),
    .B(net566),
    .Y(_03600_));
 sky130_fd_sc_hd__xnor2_1 _12098_ (.A(_03599_),
    .B(_03600_),
    .Y(_03601_));
 sky130_fd_sc_hd__a21o_1 _12099_ (.A1(_03543_),
    .A2(_03590_),
    .B1(_03595_),
    .X(_03602_));
 sky130_fd_sc_hd__nand3_1 _12100_ (.A(_03596_),
    .B(_03601_),
    .C(_03602_),
    .Y(_03603_));
 sky130_fd_sc_hd__a21bo_1 _12101_ (.A1(_03601_),
    .A2(_03602_),
    .B1_N(_03596_),
    .X(_03604_));
 sky130_fd_sc_hd__and3_2 _12102_ (.A(_03553_),
    .B(_03589_),
    .C(_03604_),
    .X(_03605_));
 sky130_fd_sc_hd__a31oi_2 _12103_ (.A1(net426),
    .A2(net566),
    .A3(_03598_),
    .B1(_03597_),
    .Y(_03606_));
 sky130_fd_sc_hd__xnor2_1 _12104_ (.A(_03562_),
    .B(_03564_),
    .Y(_03607_));
 sky130_fd_sc_hd__and2b_1 _12105_ (.A_N(_03606_),
    .B(_03607_),
    .X(_03608_));
 sky130_fd_sc_hd__xnor2_1 _12106_ (.A(_03606_),
    .B(_03607_),
    .Y(_03609_));
 sky130_fd_sc_hd__and4_1 _12107_ (.A(net421),
    .B(net417),
    .C(net571),
    .D(net576),
    .X(_03610_));
 sky130_fd_sc_hd__a22oi_1 _12108_ (.A1(net421),
    .A2(net571),
    .B1(net576),
    .B2(net417),
    .Y(_03611_));
 sky130_fd_sc_hd__and4bb_1 _12109_ (.A_N(_03610_),
    .B_N(_03611_),
    .C(net413),
    .D(net582),
    .X(_03612_));
 sky130_fd_sc_hd__nor2_1 _12110_ (.A(_03610_),
    .B(_03612_),
    .Y(_03613_));
 sky130_fd_sc_hd__and2b_1 _12111_ (.A_N(_03613_),
    .B(_03609_),
    .X(_03614_));
 sky130_fd_sc_hd__xor2_1 _12112_ (.A(_03609_),
    .B(_03613_),
    .X(_03615_));
 sky130_fd_sc_hd__a21oi_1 _12113_ (.A1(_03553_),
    .A2(_03589_),
    .B1(_03604_),
    .Y(_03616_));
 sky130_fd_sc_hd__nor3_1 _12114_ (.A(_03605_),
    .B(_03615_),
    .C(_03616_),
    .Y(_03617_));
 sky130_fd_sc_hd__or3_1 _12115_ (.A(_03605_),
    .B(_03615_),
    .C(_03616_),
    .X(_03618_));
 sky130_fd_sc_hd__o211a_1 _12116_ (.A1(_03605_),
    .A2(_03617_),
    .B1(_03569_),
    .C1(_03588_),
    .X(_03619_));
 sky130_fd_sc_hd__a22oi_1 _12117_ (.A1(net408),
    .A2(net577),
    .B1(net581),
    .B2(net404),
    .Y(_03620_));
 sky130_fd_sc_hd__nor2_1 _12118_ (.A(_03523_),
    .B(_03620_),
    .Y(_03621_));
 sky130_fd_sc_hd__o21ai_1 _12119_ (.A1(_03608_),
    .A2(_03614_),
    .B1(_03621_),
    .Y(_03622_));
 sky130_fd_sc_hd__or3_1 _12120_ (.A(_03608_),
    .B(_03614_),
    .C(_03621_),
    .X(_03623_));
 sky130_fd_sc_hd__nand2_1 _12121_ (.A(_03622_),
    .B(_03623_),
    .Y(_03624_));
 sky130_fd_sc_hd__a211oi_2 _12122_ (.A1(_03569_),
    .A2(_03588_),
    .B1(_03605_),
    .C1(_03617_),
    .Y(_03625_));
 sky130_fd_sc_hd__nor3_1 _12123_ (.A(_03619_),
    .B(_03624_),
    .C(_03625_),
    .Y(_03626_));
 sky130_fd_sc_hd__or3_1 _12124_ (.A(_03619_),
    .B(_03624_),
    .C(_03625_),
    .X(_03627_));
 sky130_fd_sc_hd__o211a_1 _12125_ (.A1(_03619_),
    .A2(_03626_),
    .B1(_03578_),
    .C1(_03587_),
    .X(_03628_));
 sky130_fd_sc_hd__a211oi_1 _12126_ (.A1(_03578_),
    .A2(_03587_),
    .B1(_03619_),
    .C1(_03626_),
    .Y(_03629_));
 sky130_fd_sc_hd__or3_1 _12127_ (.A(_03622_),
    .B(_03628_),
    .C(_03629_),
    .X(_03630_));
 sky130_fd_sc_hd__and2b_1 _12128_ (.A_N(_03628_),
    .B(_03630_),
    .X(_03631_));
 sky130_fd_sc_hd__nor2_1 _12129_ (.A(_03586_),
    .B(_03631_),
    .Y(_03632_));
 sky130_fd_sc_hd__nand2_1 _12130_ (.A(_03586_),
    .B(_03631_),
    .Y(_03633_));
 sky130_fd_sc_hd__o21ai_1 _12131_ (.A1(_03628_),
    .A2(_03629_),
    .B1(_03622_),
    .Y(_03634_));
 sky130_fd_sc_hd__o21ai_1 _12132_ (.A1(_03619_),
    .A2(_03625_),
    .B1(_03624_),
    .Y(_03635_));
 sky130_fd_sc_hd__o21ai_1 _12133_ (.A1(_03605_),
    .A2(_03616_),
    .B1(_03615_),
    .Y(_03636_));
 sky130_fd_sc_hd__a21o_1 _12134_ (.A1(_03596_),
    .A2(_03602_),
    .B1(_03601_),
    .X(_03637_));
 sky130_fd_sc_hd__a21o_1 _12135_ (.A1(_03591_),
    .A2(_03593_),
    .B1(_03592_),
    .X(_03638_));
 sky130_fd_sc_hd__nand4_1 _12136_ (.A(net450),
    .B(net445),
    .C(net553),
    .D(net557),
    .Y(_03639_));
 sky130_fd_sc_hd__and2_1 _12137_ (.A(net440),
    .B(net561),
    .X(_03640_));
 sky130_fd_sc_hd__a22o_1 _12138_ (.A1(net448),
    .A2(net553),
    .B1(net557),
    .B2(net443),
    .X(_03641_));
 sky130_fd_sc_hd__nand3_1 _12139_ (.A(_03639_),
    .B(_03640_),
    .C(_03641_),
    .Y(_03642_));
 sky130_fd_sc_hd__a21bo_1 _12140_ (.A1(_03640_),
    .A2(_03641_),
    .B1_N(_03639_),
    .X(_03643_));
 sky130_fd_sc_hd__nand3_1 _12141_ (.A(_03594_),
    .B(_03638_),
    .C(_03643_),
    .Y(_03644_));
 sky130_fd_sc_hd__a22oi_1 _12142_ (.A1(net436),
    .A2(net561),
    .B1(net566),
    .B2(net431),
    .Y(_03645_));
 sky130_fd_sc_hd__and4_1 _12143_ (.A(net436),
    .B(net431),
    .C(net561),
    .D(net566),
    .X(_03646_));
 sky130_fd_sc_hd__nor2_1 _12144_ (.A(_03645_),
    .B(_03646_),
    .Y(_03647_));
 sky130_fd_sc_hd__nand2_1 _12145_ (.A(net426),
    .B(net571),
    .Y(_03648_));
 sky130_fd_sc_hd__xnor2_1 _12146_ (.A(_03647_),
    .B(_03648_),
    .Y(_03649_));
 sky130_fd_sc_hd__a21o_1 _12147_ (.A1(_03594_),
    .A2(_03638_),
    .B1(_03643_),
    .X(_03650_));
 sky130_fd_sc_hd__nand3_1 _12148_ (.A(_03644_),
    .B(_03649_),
    .C(_03650_),
    .Y(_03651_));
 sky130_fd_sc_hd__a21bo_1 _12149_ (.A1(_03649_),
    .A2(_03650_),
    .B1_N(_03644_),
    .X(_03652_));
 sky130_fd_sc_hd__and3_1 _12150_ (.A(_03603_),
    .B(_03637_),
    .C(_03652_),
    .X(_03653_));
 sky130_fd_sc_hd__a31o_1 _12151_ (.A1(net426),
    .A2(net571),
    .A3(_03647_),
    .B1(_03646_),
    .X(_03654_));
 sky130_fd_sc_hd__o2bb2a_1 _12152_ (.A1_N(net413),
    .A2_N(net582),
    .B1(_03610_),
    .B2(_03611_),
    .X(_03655_));
 sky130_fd_sc_hd__nor2_1 _12153_ (.A(_03612_),
    .B(_03655_),
    .Y(_03656_));
 sky130_fd_sc_hd__xnor2_1 _12154_ (.A(_03654_),
    .B(_03656_),
    .Y(_03657_));
 sky130_fd_sc_hd__and4_1 _12155_ (.A(net421),
    .B(net417),
    .C(net576),
    .D(net582),
    .X(_03658_));
 sky130_fd_sc_hd__and2b_1 _12156_ (.A_N(_03657_),
    .B(_03658_),
    .X(_03659_));
 sky130_fd_sc_hd__xor2_1 _12157_ (.A(_03657_),
    .B(_03658_),
    .X(_03660_));
 sky130_fd_sc_hd__a21oi_1 _12158_ (.A1(_03603_),
    .A2(_03637_),
    .B1(_03652_),
    .Y(_03661_));
 sky130_fd_sc_hd__nor3_1 _12159_ (.A(_03653_),
    .B(_03660_),
    .C(_03661_),
    .Y(_03662_));
 sky130_fd_sc_hd__or3_1 _12160_ (.A(_03653_),
    .B(_03660_),
    .C(_03661_),
    .X(_03663_));
 sky130_fd_sc_hd__o211a_1 _12161_ (.A1(_03653_),
    .A2(_03662_),
    .B1(_03618_),
    .C1(_03636_),
    .X(_03664_));
 sky130_fd_sc_hd__nand2_1 _12162_ (.A(net412),
    .B(net582),
    .Y(_03665_));
 sky130_fd_sc_hd__a21oi_1 _12163_ (.A1(_03654_),
    .A2(_03656_),
    .B1(_03659_),
    .Y(_03666_));
 sky130_fd_sc_hd__nor2_1 _12164_ (.A(_03665_),
    .B(_03666_),
    .Y(_03667_));
 sky130_fd_sc_hd__xnor2_1 _12165_ (.A(_03665_),
    .B(_03666_),
    .Y(_03668_));
 sky130_fd_sc_hd__a211oi_1 _12166_ (.A1(_03618_),
    .A2(_03636_),
    .B1(_03653_),
    .C1(_03662_),
    .Y(_03669_));
 sky130_fd_sc_hd__nor3_1 _12167_ (.A(_03664_),
    .B(_03668_),
    .C(_03669_),
    .Y(_03670_));
 sky130_fd_sc_hd__or3_1 _12168_ (.A(_03664_),
    .B(_03668_),
    .C(_03669_),
    .X(_03671_));
 sky130_fd_sc_hd__o211a_1 _12169_ (.A1(_03664_),
    .A2(_03670_),
    .B1(_03627_),
    .C1(_03635_),
    .X(_03672_));
 sky130_fd_sc_hd__a211o_1 _12170_ (.A1(_03627_),
    .A2(_03635_),
    .B1(_03664_),
    .C1(_03670_),
    .X(_03673_));
 sky130_fd_sc_hd__nand2b_1 _12171_ (.A_N(_03672_),
    .B(_03673_),
    .Y(_03674_));
 sky130_fd_sc_hd__and3b_1 _12172_ (.A_N(_03672_),
    .B(_03673_),
    .C(_03667_),
    .X(_03675_));
 sky130_fd_sc_hd__o211a_1 _12173_ (.A1(_03672_),
    .A2(_03675_),
    .B1(_03630_),
    .C1(_03634_),
    .X(_03676_));
 sky130_fd_sc_hd__a211o_1 _12174_ (.A1(_03630_),
    .A2(_03634_),
    .B1(_03672_),
    .C1(_03675_),
    .X(_03677_));
 sky130_fd_sc_hd__xnor2_1 _12175_ (.A(_03667_),
    .B(_03674_),
    .Y(_03678_));
 sky130_fd_sc_hd__o21ai_1 _12176_ (.A1(_03664_),
    .A2(_03669_),
    .B1(_03668_),
    .Y(_03679_));
 sky130_fd_sc_hd__o21ai_1 _12177_ (.A1(_03653_),
    .A2(_03661_),
    .B1(_03660_),
    .Y(_03680_));
 sky130_fd_sc_hd__a21o_1 _12178_ (.A1(_03644_),
    .A2(_03650_),
    .B1(_03649_),
    .X(_03681_));
 sky130_fd_sc_hd__a21o_1 _12179_ (.A1(_03639_),
    .A2(_03641_),
    .B1(_03640_),
    .X(_03682_));
 sky130_fd_sc_hd__nand4_2 _12180_ (.A(net450),
    .B(net445),
    .C(net557),
    .D(net561),
    .Y(_03683_));
 sky130_fd_sc_hd__and2_1 _12181_ (.A(net440),
    .B(net566),
    .X(_03684_));
 sky130_fd_sc_hd__a22o_1 _12182_ (.A1(net450),
    .A2(net557),
    .B1(net561),
    .B2(net445),
    .X(_03685_));
 sky130_fd_sc_hd__nand3_1 _12183_ (.A(_03683_),
    .B(_03684_),
    .C(_03685_),
    .Y(_03686_));
 sky130_fd_sc_hd__a21bo_1 _12184_ (.A1(_03684_),
    .A2(_03685_),
    .B1_N(_03683_),
    .X(_03687_));
 sky130_fd_sc_hd__nand3_1 _12185_ (.A(_03642_),
    .B(_03682_),
    .C(_03687_),
    .Y(_03688_));
 sky130_fd_sc_hd__and4_1 _12186_ (.A(net436),
    .B(net431),
    .C(net566),
    .D(net571),
    .X(_03689_));
 sky130_fd_sc_hd__a22oi_1 _12187_ (.A1(net436),
    .A2(net566),
    .B1(net571),
    .B2(net431),
    .Y(_03690_));
 sky130_fd_sc_hd__nor2_1 _12188_ (.A(_03689_),
    .B(_03690_),
    .Y(_03691_));
 sky130_fd_sc_hd__nand2_1 _12189_ (.A(net426),
    .B(net576),
    .Y(_03692_));
 sky130_fd_sc_hd__and3_1 _12190_ (.A(net426),
    .B(net576),
    .C(_03691_),
    .X(_03693_));
 sky130_fd_sc_hd__xnor2_1 _12191_ (.A(_03691_),
    .B(_03692_),
    .Y(_03694_));
 sky130_fd_sc_hd__a21o_1 _12192_ (.A1(_03642_),
    .A2(_03682_),
    .B1(_03687_),
    .X(_03695_));
 sky130_fd_sc_hd__nand3_1 _12193_ (.A(_03688_),
    .B(_03694_),
    .C(_03695_),
    .Y(_03696_));
 sky130_fd_sc_hd__a21bo_1 _12194_ (.A1(_03694_),
    .A2(_03695_),
    .B1_N(_03688_),
    .X(_03697_));
 sky130_fd_sc_hd__and3_2 _12195_ (.A(_03651_),
    .B(_03681_),
    .C(_03697_),
    .X(_03698_));
 sky130_fd_sc_hd__a22oi_1 _12196_ (.A1(net421),
    .A2(net576),
    .B1(net582),
    .B2(net417),
    .Y(_03699_));
 sky130_fd_sc_hd__nor2_1 _12197_ (.A(_03658_),
    .B(_03699_),
    .Y(_03700_));
 sky130_fd_sc_hd__o21ai_2 _12198_ (.A1(_03689_),
    .A2(_03693_),
    .B1(_03700_),
    .Y(_03701_));
 sky130_fd_sc_hd__or3_1 _12199_ (.A(_03689_),
    .B(_03693_),
    .C(_03700_),
    .X(_03702_));
 sky130_fd_sc_hd__nand2_1 _12200_ (.A(_03701_),
    .B(_03702_),
    .Y(_03703_));
 sky130_fd_sc_hd__a21oi_2 _12201_ (.A1(_03651_),
    .A2(_03681_),
    .B1(_03697_),
    .Y(_03704_));
 sky130_fd_sc_hd__nor3_1 _12202_ (.A(_03698_),
    .B(_03703_),
    .C(_03704_),
    .Y(_03705_));
 sky130_fd_sc_hd__or3_1 _12203_ (.A(_03698_),
    .B(_03703_),
    .C(_03704_),
    .X(_03706_));
 sky130_fd_sc_hd__o211a_1 _12204_ (.A1(_03698_),
    .A2(_03705_),
    .B1(_03663_),
    .C1(_03680_),
    .X(_03707_));
 sky130_fd_sc_hd__a211oi_2 _12205_ (.A1(_03663_),
    .A2(_03680_),
    .B1(_03698_),
    .C1(_03705_),
    .Y(_03708_));
 sky130_fd_sc_hd__nor3_1 _12206_ (.A(_03701_),
    .B(_03707_),
    .C(_03708_),
    .Y(_03709_));
 sky130_fd_sc_hd__or3_1 _12207_ (.A(_03701_),
    .B(_03707_),
    .C(_03708_),
    .X(_03710_));
 sky130_fd_sc_hd__o211a_1 _12208_ (.A1(_03707_),
    .A2(_03709_),
    .B1(_03671_),
    .C1(_03679_),
    .X(_03711_));
 sky130_fd_sc_hd__a211o_1 _12209_ (.A1(_03671_),
    .A2(_03679_),
    .B1(_03707_),
    .C1(_03709_),
    .X(_03712_));
 sky130_fd_sc_hd__o21ai_1 _12210_ (.A1(_03707_),
    .A2(_03708_),
    .B1(_03701_),
    .Y(_03713_));
 sky130_fd_sc_hd__o21ai_2 _12211_ (.A1(_03698_),
    .A2(_03704_),
    .B1(_03703_),
    .Y(_03714_));
 sky130_fd_sc_hd__a21o_1 _12212_ (.A1(_03688_),
    .A2(_03695_),
    .B1(_03694_),
    .X(_03715_));
 sky130_fd_sc_hd__a21o_1 _12213_ (.A1(_03683_),
    .A2(_03685_),
    .B1(_03684_),
    .X(_03716_));
 sky130_fd_sc_hd__and4_1 _12214_ (.A(net450),
    .B(net445),
    .C(net561),
    .D(net566),
    .X(_03717_));
 sky130_fd_sc_hd__nand2_1 _12215_ (.A(net440),
    .B(net571),
    .Y(_03718_));
 sky130_fd_sc_hd__a22oi_2 _12216_ (.A1(net450),
    .A2(net561),
    .B1(net566),
    .B2(net445),
    .Y(_03719_));
 sky130_fd_sc_hd__or3_1 _12217_ (.A(_03717_),
    .B(_03718_),
    .C(_03719_),
    .X(_03720_));
 sky130_fd_sc_hd__o21bai_1 _12218_ (.A1(_03718_),
    .A2(_03719_),
    .B1_N(_03717_),
    .Y(_03721_));
 sky130_fd_sc_hd__nand3_1 _12219_ (.A(_03686_),
    .B(_03716_),
    .C(_03721_),
    .Y(_03722_));
 sky130_fd_sc_hd__a22oi_2 _12220_ (.A1(net436),
    .A2(net571),
    .B1(net576),
    .B2(net431),
    .Y(_03723_));
 sky130_fd_sc_hd__and4_1 _12221_ (.A(net436),
    .B(net431),
    .C(net571),
    .D(net576),
    .X(_03724_));
 sky130_fd_sc_hd__nor2_1 _12222_ (.A(_03723_),
    .B(_03724_),
    .Y(_03725_));
 sky130_fd_sc_hd__nand2_1 _12223_ (.A(net426),
    .B(net582),
    .Y(_03726_));
 sky130_fd_sc_hd__xnor2_1 _12224_ (.A(_03725_),
    .B(_03726_),
    .Y(_03727_));
 sky130_fd_sc_hd__a21o_1 _12225_ (.A1(_03686_),
    .A2(_03716_),
    .B1(_03721_),
    .X(_03728_));
 sky130_fd_sc_hd__and3_1 _12226_ (.A(_03722_),
    .B(_03727_),
    .C(_03728_),
    .X(_03729_));
 sky130_fd_sc_hd__a21bo_1 _12227_ (.A1(_03727_),
    .A2(_03728_),
    .B1_N(_03722_),
    .X(_03730_));
 sky130_fd_sc_hd__and3_1 _12228_ (.A(_03696_),
    .B(_03715_),
    .C(_03730_),
    .X(_03731_));
 sky130_fd_sc_hd__nand2_1 _12229_ (.A(net421),
    .B(net582),
    .Y(_03732_));
 sky130_fd_sc_hd__o21ba_1 _12230_ (.A1(_03723_),
    .A2(_03726_),
    .B1_N(_03724_),
    .X(_03733_));
 sky130_fd_sc_hd__nor2_1 _12231_ (.A(_03732_),
    .B(_03733_),
    .Y(_03734_));
 sky130_fd_sc_hd__xnor2_1 _12232_ (.A(_03732_),
    .B(_03733_),
    .Y(_03735_));
 sky130_fd_sc_hd__a21oi_1 _12233_ (.A1(_03696_),
    .A2(_03715_),
    .B1(_03730_),
    .Y(_03736_));
 sky130_fd_sc_hd__nor3_1 _12234_ (.A(_03731_),
    .B(_03735_),
    .C(_03736_),
    .Y(_03737_));
 sky130_fd_sc_hd__o211a_1 _12235_ (.A1(_03731_),
    .A2(_03737_),
    .B1(_03706_),
    .C1(_03714_),
    .X(_03738_));
 sky130_fd_sc_hd__o211ai_1 _12236_ (.A1(_03731_),
    .A2(_03737_),
    .B1(_03706_),
    .C1(_03714_),
    .Y(_03739_));
 sky130_fd_sc_hd__a211o_1 _12237_ (.A1(_03706_),
    .A2(_03714_),
    .B1(_03731_),
    .C1(_03737_),
    .X(_03740_));
 sky130_fd_sc_hd__and3_1 _12238_ (.A(_03734_),
    .B(_03739_),
    .C(_03740_),
    .X(_03741_));
 sky130_fd_sc_hd__o211a_1 _12239_ (.A1(_03738_),
    .A2(_03741_),
    .B1(_03710_),
    .C1(_03713_),
    .X(_03742_));
 sky130_fd_sc_hd__o21a_1 _12240_ (.A1(_03731_),
    .A2(_03736_),
    .B1(_03735_),
    .X(_03743_));
 sky130_fd_sc_hd__or2_1 _12241_ (.A(_03737_),
    .B(_03743_),
    .X(_03744_));
 sky130_fd_sc_hd__and4_1 _12242_ (.A(net436),
    .B(net431),
    .C(net576),
    .D(net582),
    .X(_03745_));
 sky130_fd_sc_hd__a21oi_1 _12243_ (.A1(_03722_),
    .A2(_03728_),
    .B1(_03727_),
    .Y(_03746_));
 sky130_fd_sc_hd__o21ai_1 _12244_ (.A1(_03717_),
    .A2(_03719_),
    .B1(_03718_),
    .Y(_03747_));
 sky130_fd_sc_hd__and4_1 _12245_ (.A(net450),
    .B(net445),
    .C(net566),
    .D(net571),
    .X(_03748_));
 sky130_fd_sc_hd__nand4_1 _12246_ (.A(net448),
    .B(net443),
    .C(net566),
    .D(net571),
    .Y(_03749_));
 sky130_fd_sc_hd__a22o_1 _12247_ (.A1(net448),
    .A2(net566),
    .B1(net571),
    .B2(net443),
    .X(_03750_));
 sky130_fd_sc_hd__and4_1 _12248_ (.A(net441),
    .B(\mul0.a[1] ),
    .C(_03749_),
    .D(_03750_),
    .X(_03751_));
 sky130_fd_sc_hd__nand4_1 _12249_ (.A(net440),
    .B(\mul0.a[1] ),
    .C(_03749_),
    .D(_03750_),
    .Y(_03752_));
 sky130_fd_sc_hd__o211a_1 _12250_ (.A1(_03748_),
    .A2(_03751_),
    .B1(_03720_),
    .C1(_03747_),
    .X(_03753_));
 sky130_fd_sc_hd__a22oi_1 _12251_ (.A1(net436),
    .A2(net576),
    .B1(net582),
    .B2(net431),
    .Y(_03754_));
 sky130_fd_sc_hd__nor2_1 _12252_ (.A(_03745_),
    .B(_03754_),
    .Y(_03755_));
 sky130_fd_sc_hd__a211o_1 _12253_ (.A1(_03720_),
    .A2(_03747_),
    .B1(_03748_),
    .C1(_03751_),
    .X(_03756_));
 sky130_fd_sc_hd__and2b_1 _12254_ (.A_N(_03753_),
    .B(_03756_),
    .X(_03757_));
 sky130_fd_sc_hd__a21oi_1 _12255_ (.A1(_03755_),
    .A2(_03756_),
    .B1(_03753_),
    .Y(_03758_));
 sky130_fd_sc_hd__or3_1 _12256_ (.A(_03729_),
    .B(_03746_),
    .C(_03758_),
    .X(_03759_));
 sky130_fd_sc_hd__o21ai_1 _12257_ (.A1(_03729_),
    .A2(_03746_),
    .B1(_03758_),
    .Y(_03760_));
 sky130_fd_sc_hd__and3_1 _12258_ (.A(_03745_),
    .B(_03759_),
    .C(_03760_),
    .X(_03761_));
 sky130_fd_sc_hd__xnor2_1 _12259_ (.A(_03755_),
    .B(_03757_),
    .Y(_03762_));
 sky130_fd_sc_hd__a22o_1 _12260_ (.A1(net440),
    .A2(net576),
    .B1(_03749_),
    .B2(_03750_),
    .X(_03763_));
 sky130_fd_sc_hd__and4_1 _12261_ (.A(net448),
    .B(net443),
    .C(net575),
    .D(net576),
    .X(_03764_));
 sky130_fd_sc_hd__a22o_1 _12262_ (.A1(net448),
    .A2(net575),
    .B1(\mul0.a[1] ),
    .B2(net443),
    .X(_03765_));
 sky130_fd_sc_hd__a31o_1 _12263_ (.A1(net440),
    .A2(net582),
    .A3(_03765_),
    .B1(_03764_),
    .X(_03766_));
 sky130_fd_sc_hd__nand3_2 _12264_ (.A(_03752_),
    .B(_03763_),
    .C(_03766_),
    .Y(_03767_));
 sky130_fd_sc_hd__a21o_1 _12265_ (.A1(_03752_),
    .A2(_03763_),
    .B1(_03766_),
    .X(_03768_));
 sky130_fd_sc_hd__a22oi_2 _12266_ (.A1(net436),
    .A2(net582),
    .B1(_03767_),
    .B2(_03768_),
    .Y(_03769_));
 sky130_fd_sc_hd__nand4_1 _12267_ (.A(net436),
    .B(net582),
    .C(_03767_),
    .D(_03768_),
    .Y(_03770_));
 sky130_fd_sc_hd__or2_1 _12268_ (.A(net440),
    .B(net575),
    .X(_03771_));
 sky130_fd_sc_hd__and4_1 _12269_ (.A(net450),
    .B(net443),
    .C(net576),
    .D(net582),
    .X(_03772_));
 sky130_fd_sc_hd__a21bo_1 _12270_ (.A1(_03718_),
    .A2(_03771_),
    .B1_N(_03772_),
    .X(_03773_));
 sky130_fd_sc_hd__nor2_1 _12271_ (.A(_03769_),
    .B(_03773_),
    .Y(_03774_));
 sky130_fd_sc_hd__a21boi_1 _12272_ (.A1(_03770_),
    .A2(_03774_),
    .B1_N(_03762_),
    .Y(_03775_));
 sky130_fd_sc_hd__o311a_1 _12273_ (.A1(_03762_),
    .A2(_03769_),
    .A3(_03773_),
    .B1(_03770_),
    .C1(_03767_),
    .X(_03776_));
 sky130_fd_sc_hd__a21oi_1 _12274_ (.A1(_03759_),
    .A2(_03760_),
    .B1(_03745_),
    .Y(_03777_));
 sky130_fd_sc_hd__or4_1 _12275_ (.A(_03761_),
    .B(_03775_),
    .C(_03776_),
    .D(_03777_),
    .X(_03778_));
 sky130_fd_sc_hd__a21boi_1 _12276_ (.A1(_03745_),
    .A2(_03760_),
    .B1_N(_03759_),
    .Y(_03779_));
 sky130_fd_sc_hd__o21a_1 _12277_ (.A1(_03744_),
    .A2(_03778_),
    .B1(_03779_),
    .X(_03780_));
 sky130_fd_sc_hd__a21oi_1 _12278_ (.A1(_03739_),
    .A2(_03740_),
    .B1(_03734_),
    .Y(_03781_));
 sky130_fd_sc_hd__a2111oi_1 _12279_ (.A1(_03744_),
    .A2(_03778_),
    .B1(_03780_),
    .C1(_03781_),
    .D1(_03741_),
    .Y(_03782_));
 sky130_fd_sc_hd__a21o_1 _12280_ (.A1(_03710_),
    .A2(_03713_),
    .B1(_03738_),
    .X(_03783_));
 sky130_fd_sc_hd__a21o_1 _12281_ (.A1(_03782_),
    .A2(_03783_),
    .B1(_03742_),
    .X(_03784_));
 sky130_fd_sc_hd__a21o_1 _12282_ (.A1(_03712_),
    .A2(_03784_),
    .B1(_03711_),
    .X(_03785_));
 sky130_fd_sc_hd__a31o_1 _12283_ (.A1(_03677_),
    .A2(_03678_),
    .A3(_03785_),
    .B1(_03676_),
    .X(_03786_));
 sky130_fd_sc_hd__a21oi_1 _12284_ (.A1(_03633_),
    .A2(_03786_),
    .B1(_03632_),
    .Y(_03787_));
 sky130_fd_sc_hd__o21ai_2 _12285_ (.A1(_03585_),
    .A2(_03787_),
    .B1(_03584_),
    .Y(_03788_));
 sky130_fd_sc_hd__or3_1 _12286_ (.A(_03485_),
    .B(_03531_),
    .C(_03534_),
    .X(_03789_));
 sky130_fd_sc_hd__and3b_1 _12287_ (.A_N(_03535_),
    .B(_03536_),
    .C(_03789_),
    .X(_03790_));
 sky130_fd_sc_hd__and3_2 _12288_ (.A(_03483_),
    .B(_03788_),
    .C(_03790_),
    .X(_03791_));
 sky130_fd_sc_hd__xnor2_4 _12289_ (.A(_03538_),
    .B(_03791_),
    .Y(_03792_));
 sky130_fd_sc_hd__nor2_1 _12290_ (.A(net9),
    .B(_03792_),
    .Y(_03793_));
 sky130_fd_sc_hd__nor2_2 _12291_ (.A(net600),
    .B(_03058_),
    .Y(_03794_));
 sky130_fd_sc_hd__a221o_1 _12292_ (.A1(net599),
    .A2(net802),
    .B1(_02738_),
    .B2(net6),
    .C1(_03793_),
    .X(_03795_));
 sky130_fd_sc_hd__mux2_1 _12293_ (.A0(net858),
    .A1(_03795_),
    .S(net3),
    .X(_00267_));
 sky130_fd_sc_hd__and4b_1 _12294_ (.A_N(_03412_),
    .B(_03483_),
    .C(_03535_),
    .D(_03536_),
    .X(_03796_));
 sky130_fd_sc_hd__a21oi_4 _12295_ (.A1(_03538_),
    .A2(_03791_),
    .B1(_03796_),
    .Y(_03797_));
 sky130_fd_sc_hd__a21o_1 _12296_ (.A1(_03538_),
    .A2(_03791_),
    .B1(_03796_),
    .X(_03798_));
 sky130_fd_sc_hd__nor2_1 _12297_ (.A(_03204_),
    .B(_03206_),
    .Y(_03799_));
 sky130_fd_sc_hd__a31o_1 _12298_ (.A1(net371),
    .A2(net581),
    .A3(_03163_),
    .B1(_03162_),
    .X(_03800_));
 sky130_fd_sc_hd__a31oi_2 _12299_ (.A1(net386),
    .A2(net567),
    .A3(_03192_),
    .B1(_03191_),
    .Y(_03801_));
 sky130_fd_sc_hd__nand4_1 _12300_ (.A(net567),
    .B(net572),
    .C(net381),
    .D(net375),
    .Y(_03802_));
 sky130_fd_sc_hd__a22o_1 _12301_ (.A1(net567),
    .A2(net381),
    .B1(net375),
    .B2(net572),
    .X(_03803_));
 sky130_fd_sc_hd__and4_1 _12302_ (.A(net577),
    .B(net371),
    .C(_03802_),
    .D(_03803_),
    .X(_03804_));
 sky130_fd_sc_hd__a22o_1 _12303_ (.A1(net580),
    .A2(net371),
    .B1(_03802_),
    .B2(_03803_),
    .X(_03805_));
 sky130_fd_sc_hd__and2b_1 _12304_ (.A_N(_03804_),
    .B(_03805_),
    .X(_03806_));
 sky130_fd_sc_hd__or3b_1 _12305_ (.A(_03801_),
    .B(_03804_),
    .C_N(_03805_),
    .X(_03807_));
 sky130_fd_sc_hd__xnor2_2 _12306_ (.A(_03801_),
    .B(_03806_),
    .Y(_03808_));
 sky130_fd_sc_hd__xnor2_2 _12307_ (.A(_03800_),
    .B(_03808_),
    .Y(_03809_));
 sky130_fd_sc_hd__o21ai_2 _12308_ (.A1(_03119_),
    .A2(_03167_),
    .B1(_03166_),
    .Y(_03810_));
 sky130_fd_sc_hd__nor2_1 _12309_ (.A(_03809_),
    .B(_03810_),
    .Y(_03811_));
 sky130_fd_sc_hd__xor2_2 _12310_ (.A(_03809_),
    .B(_03810_),
    .X(_03812_));
 sky130_fd_sc_hd__nand2_1 _12311_ (.A(net581),
    .B(net631),
    .Y(_03813_));
 sky130_fd_sc_hd__and3_1 _12312_ (.A(net581),
    .B(net631),
    .C(_03812_),
    .X(_03814_));
 sky130_fd_sc_hd__xnor2_2 _12313_ (.A(_03812_),
    .B(_03813_),
    .Y(_03815_));
 sky130_fd_sc_hd__and2b_1 _12314_ (.A_N(_03799_),
    .B(_03815_),
    .X(_03816_));
 sky130_fd_sc_hd__xnor2_2 _12315_ (.A(_03799_),
    .B(_03815_),
    .Y(_03817_));
 sky130_fd_sc_hd__or2_1 _12316_ (.A(_03122_),
    .B(_03169_),
    .X(_03818_));
 sky130_fd_sc_hd__xnor2_2 _12317_ (.A(_03817_),
    .B(_03818_),
    .Y(_03819_));
 sky130_fd_sc_hd__nand2_1 _12318_ (.A(_03200_),
    .B(_03202_),
    .Y(_03820_));
 sky130_fd_sc_hd__and4_1 _12319_ (.A(net554),
    .B(net560),
    .C(net396),
    .D(net390),
    .X(_03821_));
 sky130_fd_sc_hd__inv_2 _12320_ (.A(_03821_),
    .Y(_03822_));
 sky130_fd_sc_hd__a22o_1 _12321_ (.A1(net553),
    .A2(net396),
    .B1(net390),
    .B2(net560),
    .X(_03823_));
 sky130_fd_sc_hd__and4b_1 _12322_ (.A_N(_03821_),
    .B(_03823_),
    .C(net564),
    .D(net389),
    .X(_03824_));
 sky130_fd_sc_hd__a22oi_1 _12323_ (.A1(net564),
    .A2(net386),
    .B1(_03822_),
    .B2(_03823_),
    .Y(_03825_));
 sky130_fd_sc_hd__nor2_1 _12324_ (.A(_03824_),
    .B(_03825_),
    .Y(_03826_));
 sky130_fd_sc_hd__nand2_1 _12325_ (.A(net549),
    .B(net401),
    .Y(_03827_));
 sky130_fd_sc_hd__and4_1 _12326_ (.A(net541),
    .B(net545),
    .C(net409),
    .D(net404),
    .X(_03828_));
 sky130_fd_sc_hd__a22o_1 _12327_ (.A1(net541),
    .A2(net409),
    .B1(net404),
    .B2(net545),
    .X(_03829_));
 sky130_fd_sc_hd__and2b_1 _12328_ (.A_N(_03828_),
    .B(_03829_),
    .X(_03830_));
 sky130_fd_sc_hd__xnor2_1 _12329_ (.A(_03827_),
    .B(_03830_),
    .Y(_03831_));
 sky130_fd_sc_hd__and2_1 _12330_ (.A(_03195_),
    .B(_03197_),
    .X(_03832_));
 sky130_fd_sc_hd__and2b_1 _12331_ (.A_N(_03832_),
    .B(_03831_),
    .X(_03833_));
 sky130_fd_sc_hd__xnor2_1 _12332_ (.A(_03831_),
    .B(_03832_),
    .Y(_03834_));
 sky130_fd_sc_hd__and2_1 _12333_ (.A(_03826_),
    .B(_03834_),
    .X(_03835_));
 sky130_fd_sc_hd__xnor2_1 _12334_ (.A(_03826_),
    .B(_03834_),
    .Y(_03836_));
 sky130_fd_sc_hd__a21o_1 _12335_ (.A1(_03218_),
    .A2(_03220_),
    .B1(_03836_),
    .X(_03837_));
 sky130_fd_sc_hd__nand3_1 _12336_ (.A(_03218_),
    .B(_03220_),
    .C(_03836_),
    .Y(_03838_));
 sky130_fd_sc_hd__and3_1 _12337_ (.A(_03820_),
    .B(_03837_),
    .C(_03838_),
    .X(_03839_));
 sky130_fd_sc_hd__nand3_1 _12338_ (.A(_03820_),
    .B(_03837_),
    .C(_03838_),
    .Y(_03840_));
 sky130_fd_sc_hd__a21oi_2 _12339_ (.A1(_03837_),
    .A2(_03838_),
    .B1(_03820_),
    .Y(_03841_));
 sky130_fd_sc_hd__a31o_1 _12340_ (.A1(net414),
    .A2(net541),
    .A3(_03215_),
    .B1(_03214_),
    .X(_03842_));
 sky130_fd_sc_hd__o21ba_1 _12341_ (.A1(_03222_),
    .A2(_03223_),
    .B1_N(_03224_),
    .X(_03843_));
 sky130_fd_sc_hd__nand2_1 _12342_ (.A(net536),
    .B(net414),
    .Y(_03844_));
 sky130_fd_sc_hd__and4_1 _12343_ (.A(net525),
    .B(net531),
    .C(net422),
    .D(net418),
    .X(_03845_));
 sky130_fd_sc_hd__a22o_1 _12344_ (.A1(net525),
    .A2(net422),
    .B1(net418),
    .B2(net531),
    .X(_03846_));
 sky130_fd_sc_hd__and2b_1 _12345_ (.A_N(_03845_),
    .B(_03846_),
    .X(_03847_));
 sky130_fd_sc_hd__xnor2_2 _12346_ (.A(_03844_),
    .B(_03847_),
    .Y(_03848_));
 sky130_fd_sc_hd__nand2b_1 _12347_ (.A_N(_03843_),
    .B(_03848_),
    .Y(_03849_));
 sky130_fd_sc_hd__xnor2_2 _12348_ (.A(_03843_),
    .B(_03848_),
    .Y(_03850_));
 sky130_fd_sc_hd__nand2_1 _12349_ (.A(_03842_),
    .B(_03850_),
    .Y(_03851_));
 sky130_fd_sc_hd__xor2_2 _12350_ (.A(_03842_),
    .B(_03850_),
    .X(_03852_));
 sky130_fd_sc_hd__nand2_1 _12351_ (.A(net520),
    .B(net427),
    .Y(_03853_));
 sky130_fd_sc_hd__a22oi_2 _12352_ (.A1(net511),
    .A2(net437),
    .B1(net432),
    .B2(net515),
    .Y(_03854_));
 sky130_fd_sc_hd__and4_1 _12353_ (.A(net511),
    .B(net515),
    .C(net437),
    .D(net432),
    .X(_03855_));
 sky130_fd_sc_hd__nor2_1 _12354_ (.A(_03854_),
    .B(_03855_),
    .Y(_03856_));
 sky130_fd_sc_hd__xnor2_2 _12355_ (.A(_03853_),
    .B(_03856_),
    .Y(_03857_));
 sky130_fd_sc_hd__and2_1 _12356_ (.A(net507),
    .B(net441),
    .X(_03858_));
 sky130_fd_sc_hd__nand4_2 _12357_ (.A(net449),
    .B(net503),
    .C(net444),
    .D(net498),
    .Y(_03859_));
 sky130_fd_sc_hd__a22o_1 _12358_ (.A1(net503),
    .A2(net444),
    .B1(net498),
    .B2(net449),
    .X(_03860_));
 sky130_fd_sc_hd__nand3_1 _12359_ (.A(_03858_),
    .B(_03859_),
    .C(_03860_),
    .Y(_03861_));
 sky130_fd_sc_hd__a21o_1 _12360_ (.A1(_03859_),
    .A2(_03860_),
    .B1(_03858_),
    .X(_03862_));
 sky130_fd_sc_hd__a21bo_1 _12361_ (.A1(_03227_),
    .A2(_03229_),
    .B1_N(_03228_),
    .X(_03863_));
 sky130_fd_sc_hd__nand3_2 _12362_ (.A(_03861_),
    .B(_03862_),
    .C(_03863_),
    .Y(_03864_));
 sky130_fd_sc_hd__a21o_1 _12363_ (.A1(_03861_),
    .A2(_03862_),
    .B1(_03863_),
    .X(_03865_));
 sky130_fd_sc_hd__nand3_2 _12364_ (.A(_03857_),
    .B(_03864_),
    .C(_03865_),
    .Y(_03866_));
 sky130_fd_sc_hd__a21o_1 _12365_ (.A1(_03864_),
    .A2(_03865_),
    .B1(_03857_),
    .X(_03867_));
 sky130_fd_sc_hd__a21bo_1 _12366_ (.A1(_03226_),
    .A2(_03238_),
    .B1_N(_03237_),
    .X(_03868_));
 sky130_fd_sc_hd__nand3_4 _12367_ (.A(_03866_),
    .B(_03867_),
    .C(_03868_),
    .Y(_03869_));
 sky130_fd_sc_hd__a21o_1 _12368_ (.A1(_03866_),
    .A2(_03867_),
    .B1(_03868_),
    .X(_03870_));
 sky130_fd_sc_hd__and3_1 _12369_ (.A(_03852_),
    .B(_03869_),
    .C(_03870_),
    .X(_03871_));
 sky130_fd_sc_hd__nand3_2 _12370_ (.A(_03852_),
    .B(_03869_),
    .C(_03870_),
    .Y(_03872_));
 sky130_fd_sc_hd__a21oi_2 _12371_ (.A1(_03869_),
    .A2(_03870_),
    .B1(_03852_),
    .Y(_03873_));
 sky130_fd_sc_hd__a211oi_4 _12372_ (.A1(_03253_),
    .A2(_03256_),
    .B1(_03871_),
    .C1(_03873_),
    .Y(_03874_));
 sky130_fd_sc_hd__inv_2 _12373_ (.A(_03874_),
    .Y(_03875_));
 sky130_fd_sc_hd__o211a_1 _12374_ (.A1(_03871_),
    .A2(_03873_),
    .B1(_03253_),
    .C1(_03256_),
    .X(_03876_));
 sky130_fd_sc_hd__or4_4 _12375_ (.A(_03839_),
    .B(_03841_),
    .C(_03874_),
    .D(_03876_),
    .X(_03877_));
 sky130_fd_sc_hd__o22ai_4 _12376_ (.A1(_03839_),
    .A2(_03841_),
    .B1(_03874_),
    .B2(_03876_),
    .Y(_03878_));
 sky130_fd_sc_hd__o211ai_4 _12377_ (.A1(_03276_),
    .A2(_03278_),
    .B1(_03877_),
    .C1(_03878_),
    .Y(_03879_));
 sky130_fd_sc_hd__a211o_1 _12378_ (.A1(_03877_),
    .A2(_03878_),
    .B1(_03276_),
    .C1(_03278_),
    .X(_03880_));
 sky130_fd_sc_hd__nand3_4 _12379_ (.A(_03819_),
    .B(_03879_),
    .C(_03880_),
    .Y(_03881_));
 sky130_fd_sc_hd__a21o_1 _12380_ (.A1(_03879_),
    .A2(_03880_),
    .B1(_03819_),
    .X(_03882_));
 sky130_fd_sc_hd__o211ai_4 _12381_ (.A1(_03305_),
    .A2(_03308_),
    .B1(_03881_),
    .C1(_03882_),
    .Y(_03883_));
 sky130_fd_sc_hd__a211o_1 _12382_ (.A1(_03881_),
    .A2(_03882_),
    .B1(_03305_),
    .C1(_03308_),
    .X(_03884_));
 sky130_fd_sc_hd__o211ai_4 _12383_ (.A1(_03172_),
    .A2(_03174_),
    .B1(_03883_),
    .C1(_03884_),
    .Y(_03885_));
 sky130_fd_sc_hd__a211o_1 _12384_ (.A1(_03883_),
    .A2(_03884_),
    .B1(_03172_),
    .C1(_03174_),
    .X(_03886_));
 sky130_fd_sc_hd__o211ai_4 _12385_ (.A1(_03340_),
    .A2(_03342_),
    .B1(_03885_),
    .C1(_03886_),
    .Y(_03887_));
 sky130_fd_sc_hd__a211o_1 _12386_ (.A1(_03885_),
    .A2(_03886_),
    .B1(_03340_),
    .C1(_03342_),
    .X(_03888_));
 sky130_fd_sc_hd__nand2_2 _12387_ (.A(_03887_),
    .B(_03888_),
    .Y(_03889_));
 sky130_fd_sc_hd__nand2b_1 _12388_ (.A_N(_03412_),
    .B(_03481_),
    .Y(_03890_));
 sky130_fd_sc_hd__a21oi_2 _12389_ (.A1(_03411_),
    .A2(_03481_),
    .B1(_03409_),
    .Y(_03891_));
 sky130_fd_sc_hd__xnor2_4 _12390_ (.A(_03889_),
    .B(_03891_),
    .Y(_03892_));
 sky130_fd_sc_hd__xnor2_4 _12391_ (.A(_03797_),
    .B(_03892_),
    .Y(_03893_));
 sky130_fd_sc_hd__nor2_1 _12392_ (.A(net9),
    .B(_03893_),
    .Y(_03894_));
 sky130_fd_sc_hd__a221o_1 _12393_ (.A1(net599),
    .A2(net778),
    .B1(_02739_),
    .B2(net6),
    .C1(_03894_),
    .X(_03895_));
 sky130_fd_sc_hd__mux2_1 _12394_ (.A0(net852),
    .A1(_03895_),
    .S(net3),
    .X(_00268_));
 sky130_fd_sc_hd__a41o_1 _12395_ (.A1(_03121_),
    .A2(_03166_),
    .A3(_03168_),
    .A4(_03817_),
    .B1(_03816_),
    .X(_03896_));
 sky130_fd_sc_hd__a22o_1 _12396_ (.A1(net580),
    .A2(net631),
    .B1(net365),
    .B2(net581),
    .X(_03897_));
 sky130_fd_sc_hd__and4_1 _12397_ (.A(net578),
    .B(net583),
    .C(net631),
    .D(net365),
    .X(_03898_));
 sky130_fd_sc_hd__inv_2 _12398_ (.A(_03898_),
    .Y(_03899_));
 sky130_fd_sc_hd__and2_1 _12399_ (.A(_03897_),
    .B(_03899_),
    .X(_03900_));
 sky130_fd_sc_hd__a41o_1 _12400_ (.A1(net567),
    .A2(net572),
    .A3(net381),
    .A4(net375),
    .B1(_03804_),
    .X(_03901_));
 sky130_fd_sc_hd__or2_1 _12401_ (.A(_03821_),
    .B(_03824_),
    .X(_03902_));
 sky130_fd_sc_hd__nand2_1 _12402_ (.A(net572),
    .B(net371),
    .Y(_03903_));
 sky130_fd_sc_hd__and4_1 _12403_ (.A(net564),
    .B(net570),
    .C(net381),
    .D(net375),
    .X(_03904_));
 sky130_fd_sc_hd__a22o_1 _12404_ (.A1(net564),
    .A2(net381),
    .B1(net375),
    .B2(net570),
    .X(_03905_));
 sky130_fd_sc_hd__and2b_1 _12405_ (.A_N(_03904_),
    .B(_03905_),
    .X(_03906_));
 sky130_fd_sc_hd__xnor2_1 _12406_ (.A(_03903_),
    .B(_03906_),
    .Y(_03907_));
 sky130_fd_sc_hd__nand2_1 _12407_ (.A(_03902_),
    .B(_03907_),
    .Y(_03908_));
 sky130_fd_sc_hd__xor2_1 _12408_ (.A(_03902_),
    .B(_03907_),
    .X(_03909_));
 sky130_fd_sc_hd__nand2_1 _12409_ (.A(_03901_),
    .B(_03909_),
    .Y(_03910_));
 sky130_fd_sc_hd__xnor2_1 _12410_ (.A(_03901_),
    .B(_03909_),
    .Y(_03911_));
 sky130_fd_sc_hd__a21bo_1 _12411_ (.A1(_03800_),
    .A2(_03808_),
    .B1_N(_03807_),
    .X(_03912_));
 sky130_fd_sc_hd__and2b_1 _12412_ (.A_N(_03911_),
    .B(_03912_),
    .X(_03913_));
 sky130_fd_sc_hd__xnor2_1 _12413_ (.A(_03911_),
    .B(_03912_),
    .Y(_03914_));
 sky130_fd_sc_hd__xnor2_1 _12414_ (.A(_03900_),
    .B(_03914_),
    .Y(_03915_));
 sky130_fd_sc_hd__a21o_1 _12415_ (.A1(_03837_),
    .A2(_03840_),
    .B1(_03915_),
    .X(_03916_));
 sky130_fd_sc_hd__nand3_1 _12416_ (.A(_03837_),
    .B(_03840_),
    .C(_03915_),
    .Y(_03917_));
 sky130_fd_sc_hd__o211a_1 _12417_ (.A1(_03811_),
    .A2(_03814_),
    .B1(_03916_),
    .C1(_03917_),
    .X(_03918_));
 sky130_fd_sc_hd__inv_2 _12418_ (.A(_03918_),
    .Y(_03919_));
 sky130_fd_sc_hd__a211oi_2 _12419_ (.A1(_03916_),
    .A2(_03917_),
    .B1(_03811_),
    .C1(_03814_),
    .Y(_03920_));
 sky130_fd_sc_hd__and4_1 _12420_ (.A(net549),
    .B(net553),
    .C(net395),
    .D(net390),
    .X(_03921_));
 sky130_fd_sc_hd__inv_2 _12421_ (.A(_03921_),
    .Y(_03922_));
 sky130_fd_sc_hd__a22o_1 _12422_ (.A1(net549),
    .A2(net396),
    .B1(net390),
    .B2(net553),
    .X(_03923_));
 sky130_fd_sc_hd__and4b_1 _12423_ (.A_N(_03921_),
    .B(_03923_),
    .C(net557),
    .D(net389),
    .X(_03924_));
 sky130_fd_sc_hd__a22oi_1 _12424_ (.A1(net557),
    .A2(net389),
    .B1(_03922_),
    .B2(_03923_),
    .Y(_03925_));
 sky130_fd_sc_hd__nor2_1 _12425_ (.A(_03924_),
    .B(_03925_),
    .Y(_03926_));
 sky130_fd_sc_hd__nand2_1 _12426_ (.A(net545),
    .B(net400),
    .Y(_03927_));
 sky130_fd_sc_hd__and4_1 _12427_ (.A(net536),
    .B(net541),
    .C(net409),
    .D(net405),
    .X(_03928_));
 sky130_fd_sc_hd__a22o_1 _12428_ (.A1(net536),
    .A2(net412),
    .B1(net405),
    .B2(net541),
    .X(_03929_));
 sky130_fd_sc_hd__and2b_1 _12429_ (.A_N(_03928_),
    .B(_03929_),
    .X(_03930_));
 sky130_fd_sc_hd__xnor2_1 _12430_ (.A(_03927_),
    .B(_03930_),
    .Y(_03931_));
 sky130_fd_sc_hd__a31o_1 _12431_ (.A1(net548),
    .A2(net400),
    .A3(_03829_),
    .B1(_03828_),
    .X(_03932_));
 sky130_fd_sc_hd__and2_2 _12432_ (.A(_03931_),
    .B(_03932_),
    .X(_03933_));
 sky130_fd_sc_hd__xor2_1 _12433_ (.A(_03931_),
    .B(_03932_),
    .X(_03934_));
 sky130_fd_sc_hd__and2_2 _12434_ (.A(_03926_),
    .B(_03934_),
    .X(_03935_));
 sky130_fd_sc_hd__xnor2_1 _12435_ (.A(_03926_),
    .B(_03934_),
    .Y(_03936_));
 sky130_fd_sc_hd__a21o_2 _12436_ (.A1(_03849_),
    .A2(_03851_),
    .B1(_03936_),
    .X(_03937_));
 sky130_fd_sc_hd__nand3_2 _12437_ (.A(_03849_),
    .B(_03851_),
    .C(_03936_),
    .Y(_03938_));
 sky130_fd_sc_hd__o211a_1 _12438_ (.A1(_03833_),
    .A2(_03835_),
    .B1(_03937_),
    .C1(_03938_),
    .X(_03939_));
 sky130_fd_sc_hd__o211ai_2 _12439_ (.A1(_03833_),
    .A2(_03835_),
    .B1(_03937_),
    .C1(_03938_),
    .Y(_03940_));
 sky130_fd_sc_hd__a211oi_2 _12440_ (.A1(_03937_),
    .A2(_03938_),
    .B1(_03833_),
    .C1(_03835_),
    .Y(_03941_));
 sky130_fd_sc_hd__a31o_1 _12441_ (.A1(net535),
    .A2(net414),
    .A3(_03846_),
    .B1(_03845_),
    .X(_03942_));
 sky130_fd_sc_hd__o21ba_1 _12442_ (.A1(_03853_),
    .A2(_03854_),
    .B1_N(_03855_),
    .X(_03943_));
 sky130_fd_sc_hd__nand2_1 _12443_ (.A(net530),
    .B(net414),
    .Y(_03944_));
 sky130_fd_sc_hd__and4_1 _12444_ (.A(net520),
    .B(net525),
    .C(net425),
    .D(net418),
    .X(_03945_));
 sky130_fd_sc_hd__a22o_1 _12445_ (.A1(net520),
    .A2(net425),
    .B1(net418),
    .B2(net525),
    .X(_03946_));
 sky130_fd_sc_hd__and2b_1 _12446_ (.A_N(_03945_),
    .B(_03946_),
    .X(_03947_));
 sky130_fd_sc_hd__xnor2_2 _12447_ (.A(_03944_),
    .B(_03947_),
    .Y(_03948_));
 sky130_fd_sc_hd__nand2b_2 _12448_ (.A_N(_03943_),
    .B(_03948_),
    .Y(_03949_));
 sky130_fd_sc_hd__xnor2_2 _12449_ (.A(_03943_),
    .B(_03948_),
    .Y(_03950_));
 sky130_fd_sc_hd__nand2_1 _12450_ (.A(_03942_),
    .B(_03950_),
    .Y(_03951_));
 sky130_fd_sc_hd__xor2_2 _12451_ (.A(_03942_),
    .B(_03950_),
    .X(_03952_));
 sky130_fd_sc_hd__nand2_1 _12452_ (.A(net515),
    .B(net427),
    .Y(_03953_));
 sky130_fd_sc_hd__a22oi_2 _12453_ (.A1(net507),
    .A2(net437),
    .B1(net432),
    .B2(net511),
    .Y(_03954_));
 sky130_fd_sc_hd__and4_1 _12454_ (.A(net507),
    .B(net511),
    .C(net437),
    .D(net432),
    .X(_03955_));
 sky130_fd_sc_hd__nor2_1 _12455_ (.A(_03954_),
    .B(_03955_),
    .Y(_03956_));
 sky130_fd_sc_hd__xnor2_2 _12456_ (.A(_03953_),
    .B(_03956_),
    .Y(_03957_));
 sky130_fd_sc_hd__and2_1 _12457_ (.A(net503),
    .B(net441),
    .X(_03958_));
 sky130_fd_sc_hd__nand4_1 _12458_ (.A(net449),
    .B(net446),
    .C(net498),
    .D(net494),
    .Y(_03959_));
 sky130_fd_sc_hd__a22o_1 _12459_ (.A1(net444),
    .A2(net498),
    .B1(net494),
    .B2(net449),
    .X(_03960_));
 sky130_fd_sc_hd__nand3_1 _12460_ (.A(_03958_),
    .B(_03959_),
    .C(_03960_),
    .Y(_03961_));
 sky130_fd_sc_hd__a21o_1 _12461_ (.A1(_03959_),
    .A2(_03960_),
    .B1(_03958_),
    .X(_03962_));
 sky130_fd_sc_hd__a21bo_1 _12462_ (.A1(_03858_),
    .A2(_03860_),
    .B1_N(_03859_),
    .X(_03963_));
 sky130_fd_sc_hd__nand3_1 _12463_ (.A(_03961_),
    .B(_03962_),
    .C(_03963_),
    .Y(_03964_));
 sky130_fd_sc_hd__a21o_1 _12464_ (.A1(_03961_),
    .A2(_03962_),
    .B1(_03963_),
    .X(_03965_));
 sky130_fd_sc_hd__nand3_2 _12465_ (.A(_03957_),
    .B(_03964_),
    .C(_03965_),
    .Y(_03966_));
 sky130_fd_sc_hd__a21o_1 _12466_ (.A1(_03964_),
    .A2(_03965_),
    .B1(_03957_),
    .X(_03967_));
 sky130_fd_sc_hd__a21bo_1 _12467_ (.A1(_03857_),
    .A2(_03865_),
    .B1_N(_03864_),
    .X(_03968_));
 sky130_fd_sc_hd__nand3_4 _12468_ (.A(_03966_),
    .B(_03967_),
    .C(_03968_),
    .Y(_03969_));
 sky130_fd_sc_hd__a21o_1 _12469_ (.A1(_03966_),
    .A2(_03967_),
    .B1(_03968_),
    .X(_03970_));
 sky130_fd_sc_hd__and3_1 _12470_ (.A(_03952_),
    .B(_03969_),
    .C(_03970_),
    .X(_03971_));
 sky130_fd_sc_hd__nand3_2 _12471_ (.A(_03952_),
    .B(_03969_),
    .C(_03970_),
    .Y(_03972_));
 sky130_fd_sc_hd__a21oi_2 _12472_ (.A1(_03969_),
    .A2(_03970_),
    .B1(_03952_),
    .Y(_03973_));
 sky130_fd_sc_hd__a211oi_4 _12473_ (.A1(_03869_),
    .A2(_03872_),
    .B1(_03971_),
    .C1(_03973_),
    .Y(_03974_));
 sky130_fd_sc_hd__o211a_1 _12474_ (.A1(_03971_),
    .A2(_03973_),
    .B1(_03869_),
    .C1(_03872_),
    .X(_03975_));
 sky130_fd_sc_hd__nor4_4 _12475_ (.A(_03939_),
    .B(_03941_),
    .C(_03974_),
    .D(_03975_),
    .Y(_03976_));
 sky130_fd_sc_hd__o22a_1 _12476_ (.A1(_03939_),
    .A2(_03941_),
    .B1(_03974_),
    .B2(_03975_),
    .X(_03977_));
 sky130_fd_sc_hd__a211oi_4 _12477_ (.A1(_03875_),
    .A2(_03877_),
    .B1(_03976_),
    .C1(_03977_),
    .Y(_03978_));
 sky130_fd_sc_hd__o211a_1 _12478_ (.A1(_03976_),
    .A2(_03977_),
    .B1(_03875_),
    .C1(_03877_),
    .X(_03979_));
 sky130_fd_sc_hd__nor4_2 _12479_ (.A(_03918_),
    .B(_03920_),
    .C(_03978_),
    .D(_03979_),
    .Y(_03980_));
 sky130_fd_sc_hd__o22a_1 _12480_ (.A1(_03918_),
    .A2(_03920_),
    .B1(_03978_),
    .B2(_03979_),
    .X(_03981_));
 sky130_fd_sc_hd__a211oi_1 _12481_ (.A1(_03879_),
    .A2(_03881_),
    .B1(_03980_),
    .C1(_03981_),
    .Y(_03982_));
 sky130_fd_sc_hd__a211o_1 _12482_ (.A1(_03879_),
    .A2(_03881_),
    .B1(_03980_),
    .C1(_03981_),
    .X(_03983_));
 sky130_fd_sc_hd__o211ai_1 _12483_ (.A1(_03980_),
    .A2(_03981_),
    .B1(_03879_),
    .C1(_03881_),
    .Y(_03984_));
 sky130_fd_sc_hd__and3_1 _12484_ (.A(_03896_),
    .B(_03983_),
    .C(_03984_),
    .X(_03985_));
 sky130_fd_sc_hd__a21oi_1 _12485_ (.A1(_03983_),
    .A2(_03984_),
    .B1(_03896_),
    .Y(_03986_));
 sky130_fd_sc_hd__a211o_1 _12486_ (.A1(_03883_),
    .A2(_03885_),
    .B1(_03985_),
    .C1(_03986_),
    .X(_03987_));
 sky130_fd_sc_hd__o211ai_1 _12487_ (.A1(_03985_),
    .A2(_03986_),
    .B1(_03883_),
    .C1(_03885_),
    .Y(_03988_));
 sky130_fd_sc_hd__nand2_2 _12488_ (.A(_03987_),
    .B(_03988_),
    .Y(_03989_));
 sky130_fd_sc_hd__a21bo_1 _12489_ (.A1(_03409_),
    .A2(_03888_),
    .B1_N(_03887_),
    .X(_03990_));
 sky130_fd_sc_hd__xor2_4 _12490_ (.A(_03989_),
    .B(_03990_),
    .X(_03991_));
 sky130_fd_sc_hd__o22a_2 _12491_ (.A1(_03889_),
    .A2(_03890_),
    .B1(_03892_),
    .B2(_03797_),
    .X(_03992_));
 sky130_fd_sc_hd__xnor2_4 _12492_ (.A(_03991_),
    .B(_03992_),
    .Y(_03993_));
 sky130_fd_sc_hd__nor2_1 _12493_ (.A(net9),
    .B(_03993_),
    .Y(_03994_));
 sky130_fd_sc_hd__a221o_1 _12494_ (.A1(net599),
    .A2(\temp[2] ),
    .B1(_02741_),
    .B2(net6),
    .C1(_03994_),
    .X(_03995_));
 sky130_fd_sc_hd__mux2_1 _12495_ (.A0(net759),
    .A1(_03995_),
    .S(net3),
    .X(_00269_));
 sky130_fd_sc_hd__or3_1 _12496_ (.A(_03410_),
    .B(_03889_),
    .C(_03989_),
    .X(_03996_));
 sky130_fd_sc_hd__nor2_1 _12497_ (.A(_03892_),
    .B(_03991_),
    .Y(_03997_));
 sky130_fd_sc_hd__o31ai_1 _12498_ (.A1(_03889_),
    .A2(_03890_),
    .A3(_03991_),
    .B1(_03996_),
    .Y(_03998_));
 sky130_fd_sc_hd__a21o_2 _12499_ (.A1(_03798_),
    .A2(_03997_),
    .B1(_03998_),
    .X(_03999_));
 sky130_fd_sc_hd__a21oi_1 _12500_ (.A1(_03900_),
    .A2(_03914_),
    .B1(_03913_),
    .Y(_04000_));
 sky130_fd_sc_hd__nand4_1 _12501_ (.A(net574),
    .B(net578),
    .C(net631),
    .D(net365),
    .Y(_04001_));
 sky130_fd_sc_hd__a22o_1 _12502_ (.A1(net574),
    .A2(net631),
    .B1(net365),
    .B2(net578),
    .X(_04002_));
 sky130_fd_sc_hd__nand2_1 _12503_ (.A(_04001_),
    .B(_04002_),
    .Y(_04003_));
 sky130_fd_sc_hd__nand2_1 _12504_ (.A(net583),
    .B(net364),
    .Y(_04004_));
 sky130_fd_sc_hd__xnor2_1 _12505_ (.A(_04003_),
    .B(_04004_),
    .Y(_04005_));
 sky130_fd_sc_hd__nor2_1 _12506_ (.A(_03899_),
    .B(_04005_),
    .Y(_04006_));
 sky130_fd_sc_hd__and2_1 _12507_ (.A(_03899_),
    .B(_04005_),
    .X(_04007_));
 sky130_fd_sc_hd__or2_1 _12508_ (.A(_04006_),
    .B(_04007_),
    .X(_04008_));
 sky130_fd_sc_hd__a31o_1 _12509_ (.A1(net572),
    .A2(net371),
    .A3(_03905_),
    .B1(_03904_),
    .X(_04009_));
 sky130_fd_sc_hd__or2_1 _12510_ (.A(_03921_),
    .B(_03924_),
    .X(_04010_));
 sky130_fd_sc_hd__nand2_1 _12511_ (.A(net567),
    .B(net370),
    .Y(_04011_));
 sky130_fd_sc_hd__and4_1 _12512_ (.A(net557),
    .B(net565),
    .C(net381),
    .D(net375),
    .X(_04012_));
 sky130_fd_sc_hd__a22o_1 _12513_ (.A1(net557),
    .A2(net381),
    .B1(net375),
    .B2(net561),
    .X(_04013_));
 sky130_fd_sc_hd__and2b_1 _12514_ (.A_N(_04012_),
    .B(_04013_),
    .X(_04014_));
 sky130_fd_sc_hd__xnor2_2 _12515_ (.A(_04011_),
    .B(_04014_),
    .Y(_04015_));
 sky130_fd_sc_hd__nand2_1 _12516_ (.A(_04010_),
    .B(_04015_),
    .Y(_04016_));
 sky130_fd_sc_hd__xor2_2 _12517_ (.A(_04010_),
    .B(_04015_),
    .X(_04017_));
 sky130_fd_sc_hd__nand2_1 _12518_ (.A(_04009_),
    .B(_04017_),
    .Y(_04018_));
 sky130_fd_sc_hd__xnor2_2 _12519_ (.A(_04009_),
    .B(_04017_),
    .Y(_04019_));
 sky130_fd_sc_hd__a21oi_4 _12520_ (.A1(_03908_),
    .A2(_03910_),
    .B1(_04019_),
    .Y(_04020_));
 sky130_fd_sc_hd__and3_1 _12521_ (.A(_03908_),
    .B(_03910_),
    .C(_04019_),
    .X(_04021_));
 sky130_fd_sc_hd__nor3_2 _12522_ (.A(_04008_),
    .B(_04020_),
    .C(_04021_),
    .Y(_04022_));
 sky130_fd_sc_hd__o21a_1 _12523_ (.A1(_04020_),
    .A2(_04021_),
    .B1(_04008_),
    .X(_04023_));
 sky130_fd_sc_hd__a211oi_2 _12524_ (.A1(_03937_),
    .A2(_03940_),
    .B1(_04022_),
    .C1(_04023_),
    .Y(_04024_));
 sky130_fd_sc_hd__o211a_1 _12525_ (.A1(_04022_),
    .A2(_04023_),
    .B1(_03937_),
    .C1(_03940_),
    .X(_04025_));
 sky130_fd_sc_hd__nor3_1 _12526_ (.A(_04000_),
    .B(_04024_),
    .C(_04025_),
    .Y(_04026_));
 sky130_fd_sc_hd__o21a_1 _12527_ (.A1(_04024_),
    .A2(_04025_),
    .B1(_04000_),
    .X(_04027_));
 sky130_fd_sc_hd__nand4_2 _12528_ (.A(net545),
    .B(net548),
    .C(net395),
    .D(net391),
    .Y(_04028_));
 sky130_fd_sc_hd__a22o_1 _12529_ (.A1(net545),
    .A2(net395),
    .B1(net391),
    .B2(net548),
    .X(_04029_));
 sky130_fd_sc_hd__nand4_2 _12530_ (.A(net553),
    .B(net386),
    .C(_04028_),
    .D(_04029_),
    .Y(_04030_));
 sky130_fd_sc_hd__a22o_1 _12531_ (.A1(net553),
    .A2(net386),
    .B1(_04028_),
    .B2(_04029_),
    .X(_04031_));
 sky130_fd_sc_hd__and2_1 _12532_ (.A(_04030_),
    .B(_04031_),
    .X(_04032_));
 sky130_fd_sc_hd__nand2_1 _12533_ (.A(net541),
    .B(net401),
    .Y(_04033_));
 sky130_fd_sc_hd__and4_1 _12534_ (.A(net531),
    .B(net536),
    .C(net409),
    .D(net405),
    .X(_04034_));
 sky130_fd_sc_hd__a22o_1 _12535_ (.A1(net531),
    .A2(net409),
    .B1(net405),
    .B2(net536),
    .X(_04035_));
 sky130_fd_sc_hd__and2b_1 _12536_ (.A_N(_04034_),
    .B(_04035_),
    .X(_04036_));
 sky130_fd_sc_hd__xnor2_2 _12537_ (.A(_04033_),
    .B(_04036_),
    .Y(_04037_));
 sky130_fd_sc_hd__a31o_1 _12538_ (.A1(net545),
    .A2(net401),
    .A3(_03929_),
    .B1(_03928_),
    .X(_04038_));
 sky130_fd_sc_hd__and2_2 _12539_ (.A(_04037_),
    .B(_04038_),
    .X(_04039_));
 sky130_fd_sc_hd__xor2_2 _12540_ (.A(_04037_),
    .B(_04038_),
    .X(_04040_));
 sky130_fd_sc_hd__and2_2 _12541_ (.A(_04032_),
    .B(_04040_),
    .X(_04041_));
 sky130_fd_sc_hd__xnor2_2 _12542_ (.A(_04032_),
    .B(_04040_),
    .Y(_04042_));
 sky130_fd_sc_hd__a21o_4 _12543_ (.A1(_03949_),
    .A2(_03951_),
    .B1(_04042_),
    .X(_04043_));
 sky130_fd_sc_hd__nand3_4 _12544_ (.A(_03949_),
    .B(_03951_),
    .C(_04042_),
    .Y(_04044_));
 sky130_fd_sc_hd__o211a_1 _12545_ (.A1(_03933_),
    .A2(_03935_),
    .B1(_04043_),
    .C1(_04044_),
    .X(_04045_));
 sky130_fd_sc_hd__o211ai_4 _12546_ (.A1(_03933_),
    .A2(_03935_),
    .B1(_04043_),
    .C1(_04044_),
    .Y(_04046_));
 sky130_fd_sc_hd__a211oi_4 _12547_ (.A1(_04043_),
    .A2(_04044_),
    .B1(_03933_),
    .C1(_03935_),
    .Y(_04047_));
 sky130_fd_sc_hd__a31o_1 _12548_ (.A1(net530),
    .A2(net414),
    .A3(_03946_),
    .B1(_03945_),
    .X(_04048_));
 sky130_fd_sc_hd__o21ba_1 _12549_ (.A1(_03953_),
    .A2(_03954_),
    .B1_N(_03955_),
    .X(_04049_));
 sky130_fd_sc_hd__nand2_1 _12550_ (.A(net526),
    .B(net414),
    .Y(_04050_));
 sky130_fd_sc_hd__and4_1 _12551_ (.A(net515),
    .B(net520),
    .C(net422),
    .D(net418),
    .X(_04051_));
 sky130_fd_sc_hd__a22o_1 _12552_ (.A1(net515),
    .A2(net422),
    .B1(net418),
    .B2(net520),
    .X(_04052_));
 sky130_fd_sc_hd__and2b_1 _12553_ (.A_N(_04051_),
    .B(_04052_),
    .X(_04053_));
 sky130_fd_sc_hd__xnor2_2 _12554_ (.A(_04050_),
    .B(_04053_),
    .Y(_04054_));
 sky130_fd_sc_hd__nand2b_2 _12555_ (.A_N(_04049_),
    .B(_04054_),
    .Y(_04055_));
 sky130_fd_sc_hd__xnor2_2 _12556_ (.A(_04049_),
    .B(_04054_),
    .Y(_04056_));
 sky130_fd_sc_hd__nand2_2 _12557_ (.A(_04048_),
    .B(_04056_),
    .Y(_04057_));
 sky130_fd_sc_hd__xor2_2 _12558_ (.A(_04048_),
    .B(_04056_),
    .X(_04058_));
 sky130_fd_sc_hd__nand2_1 _12559_ (.A(net511),
    .B(net427),
    .Y(_04059_));
 sky130_fd_sc_hd__and4_1 _12560_ (.A(net503),
    .B(net507),
    .C(net437),
    .D(net432),
    .X(_04060_));
 sky130_fd_sc_hd__a22oi_1 _12561_ (.A1(net503),
    .A2(net437),
    .B1(net432),
    .B2(net507),
    .Y(_04061_));
 sky130_fd_sc_hd__nor2_1 _12562_ (.A(_04060_),
    .B(_04061_),
    .Y(_04062_));
 sky130_fd_sc_hd__xnor2_2 _12563_ (.A(_04059_),
    .B(_04062_),
    .Y(_04063_));
 sky130_fd_sc_hd__and2_1 _12564_ (.A(net441),
    .B(net498),
    .X(_04064_));
 sky130_fd_sc_hd__nand4_2 _12565_ (.A(net452),
    .B(net446),
    .C(net494),
    .D(net490),
    .Y(_04065_));
 sky130_fd_sc_hd__a22o_1 _12566_ (.A1(net446),
    .A2(net494),
    .B1(net490),
    .B2(net452),
    .X(_04066_));
 sky130_fd_sc_hd__nand3_1 _12567_ (.A(_04064_),
    .B(_04065_),
    .C(_04066_),
    .Y(_04067_));
 sky130_fd_sc_hd__a21o_1 _12568_ (.A1(_04065_),
    .A2(_04066_),
    .B1(_04064_),
    .X(_04068_));
 sky130_fd_sc_hd__a21bo_1 _12569_ (.A1(_03958_),
    .A2(_03960_),
    .B1_N(_03959_),
    .X(_04069_));
 sky130_fd_sc_hd__nand3_2 _12570_ (.A(_04067_),
    .B(_04068_),
    .C(_04069_),
    .Y(_04070_));
 sky130_fd_sc_hd__a21o_1 _12571_ (.A1(_04067_),
    .A2(_04068_),
    .B1(_04069_),
    .X(_04071_));
 sky130_fd_sc_hd__nand3_2 _12572_ (.A(_04063_),
    .B(_04070_),
    .C(_04071_),
    .Y(_04072_));
 sky130_fd_sc_hd__a21o_1 _12573_ (.A1(_04070_),
    .A2(_04071_),
    .B1(_04063_),
    .X(_04073_));
 sky130_fd_sc_hd__a21bo_1 _12574_ (.A1(_03957_),
    .A2(_03965_),
    .B1_N(_03964_),
    .X(_04074_));
 sky130_fd_sc_hd__nand3_4 _12575_ (.A(_04072_),
    .B(_04073_),
    .C(_04074_),
    .Y(_04075_));
 sky130_fd_sc_hd__a21o_1 _12576_ (.A1(_04072_),
    .A2(_04073_),
    .B1(_04074_),
    .X(_04076_));
 sky130_fd_sc_hd__and3_1 _12577_ (.A(_04058_),
    .B(_04075_),
    .C(_04076_),
    .X(_04077_));
 sky130_fd_sc_hd__nand3_2 _12578_ (.A(_04058_),
    .B(_04075_),
    .C(_04076_),
    .Y(_04078_));
 sky130_fd_sc_hd__a21oi_2 _12579_ (.A1(_04075_),
    .A2(_04076_),
    .B1(_04058_),
    .Y(_04079_));
 sky130_fd_sc_hd__a211oi_4 _12580_ (.A1(_03969_),
    .A2(_03972_),
    .B1(_04077_),
    .C1(_04079_),
    .Y(_04080_));
 sky130_fd_sc_hd__o211a_1 _12581_ (.A1(_04077_),
    .A2(_04079_),
    .B1(_03969_),
    .C1(_03972_),
    .X(_04081_));
 sky130_fd_sc_hd__nor4_2 _12582_ (.A(_04045_),
    .B(_04047_),
    .C(_04080_),
    .D(_04081_),
    .Y(_04082_));
 sky130_fd_sc_hd__or4_2 _12583_ (.A(_04045_),
    .B(_04047_),
    .C(_04080_),
    .D(_04081_),
    .X(_04083_));
 sky130_fd_sc_hd__o22ai_4 _12584_ (.A1(_04045_),
    .A2(_04047_),
    .B1(_04080_),
    .B2(_04081_),
    .Y(_04084_));
 sky130_fd_sc_hd__o211ai_4 _12585_ (.A1(_03974_),
    .A2(_03976_),
    .B1(_04083_),
    .C1(_04084_),
    .Y(_04085_));
 sky130_fd_sc_hd__a211o_1 _12586_ (.A1(_04083_),
    .A2(_04084_),
    .B1(_03974_),
    .C1(_03976_),
    .X(_04086_));
 sky130_fd_sc_hd__or4bb_4 _12587_ (.A(_04026_),
    .B(_04027_),
    .C_N(_04085_),
    .D_N(_04086_),
    .X(_04087_));
 sky130_fd_sc_hd__a2bb2o_1 _12588_ (.A1_N(_04026_),
    .A2_N(_04027_),
    .B1(_04085_),
    .B2(_04086_),
    .X(_04088_));
 sky130_fd_sc_hd__o211a_1 _12589_ (.A1(_03978_),
    .A2(_03980_),
    .B1(_04087_),
    .C1(_04088_),
    .X(_04089_));
 sky130_fd_sc_hd__a211oi_2 _12590_ (.A1(_04087_),
    .A2(_04088_),
    .B1(_03978_),
    .C1(_03980_),
    .Y(_04090_));
 sky130_fd_sc_hd__a211oi_1 _12591_ (.A1(_03916_),
    .A2(_03919_),
    .B1(_04089_),
    .C1(_04090_),
    .Y(_04091_));
 sky130_fd_sc_hd__a211o_1 _12592_ (.A1(_03916_),
    .A2(_03919_),
    .B1(_04089_),
    .C1(_04090_),
    .X(_04092_));
 sky130_fd_sc_hd__o211ai_1 _12593_ (.A1(_04089_),
    .A2(_04090_),
    .B1(_03916_),
    .C1(_03919_),
    .Y(_04093_));
 sky130_fd_sc_hd__o211a_1 _12594_ (.A1(_03982_),
    .A2(_03985_),
    .B1(_04092_),
    .C1(_04093_),
    .X(_04094_));
 sky130_fd_sc_hd__a211oi_1 _12595_ (.A1(_04092_),
    .A2(_04093_),
    .B1(_03982_),
    .C1(_03985_),
    .Y(_04095_));
 sky130_fd_sc_hd__or2_1 _12596_ (.A(_04094_),
    .B(_04095_),
    .X(_04096_));
 sky130_fd_sc_hd__o21a_1 _12597_ (.A1(_03887_),
    .A2(_03989_),
    .B1(_03987_),
    .X(_04097_));
 sky130_fd_sc_hd__xnor2_1 _12598_ (.A(_04096_),
    .B(_04097_),
    .Y(_04098_));
 sky130_fd_sc_hd__inv_2 _12599_ (.A(_04098_),
    .Y(_04099_));
 sky130_fd_sc_hd__xnor2_4 _12600_ (.A(_03999_),
    .B(_04099_),
    .Y(_04100_));
 sky130_fd_sc_hd__nor2_1 _12601_ (.A(net9),
    .B(_04100_),
    .Y(_04101_));
 sky130_fd_sc_hd__a221o_1 _12602_ (.A1(net599),
    .A2(\temp[3] ),
    .B1(_02743_),
    .B2(net6),
    .C1(_04101_),
    .X(_04102_));
 sky130_fd_sc_hd__mux2_1 _12603_ (.A0(net720),
    .A1(_04102_),
    .S(net3),
    .X(_00270_));
 sky130_fd_sc_hd__nor2_1 _12604_ (.A(_04024_),
    .B(_04026_),
    .Y(_04103_));
 sky130_fd_sc_hd__or3_2 _12605_ (.A(_03899_),
    .B(_04005_),
    .C(_04103_),
    .X(_04104_));
 sky130_fd_sc_hd__xnor2_1 _12606_ (.A(_04006_),
    .B(_04103_),
    .Y(_04105_));
 sky130_fd_sc_hd__and4_1 _12607_ (.A(net568),
    .B(net573),
    .C(\mul0.b[18] ),
    .D(net365),
    .X(_04106_));
 sky130_fd_sc_hd__inv_2 _12608_ (.A(_04106_),
    .Y(_04107_));
 sky130_fd_sc_hd__a22o_1 _12609_ (.A1(net568),
    .A2(net631),
    .B1(net365),
    .B2(net573),
    .X(_04108_));
 sky130_fd_sc_hd__and4_1 _12610_ (.A(net578),
    .B(net364),
    .C(_04107_),
    .D(_04108_),
    .X(_04109_));
 sky130_fd_sc_hd__a22oi_1 _12611_ (.A1(net578),
    .A2(net364),
    .B1(_04107_),
    .B2(_04108_),
    .Y(_04110_));
 sky130_fd_sc_hd__or2_1 _12612_ (.A(_04109_),
    .B(_04110_),
    .X(_04111_));
 sky130_fd_sc_hd__o21ai_2 _12613_ (.A1(_04003_),
    .A2(_04004_),
    .B1(_04001_),
    .Y(_04112_));
 sky130_fd_sc_hd__and2b_1 _12614_ (.A_N(_04111_),
    .B(_04112_),
    .X(_04113_));
 sky130_fd_sc_hd__xnor2_2 _12615_ (.A(_04111_),
    .B(_04112_),
    .Y(_04114_));
 sky130_fd_sc_hd__nand2_1 _12616_ (.A(net583),
    .B(net360),
    .Y(_04115_));
 sky130_fd_sc_hd__xnor2_1 _12617_ (.A(_04114_),
    .B(_04115_),
    .Y(_04116_));
 sky130_fd_sc_hd__a31o_1 _12618_ (.A1(net568),
    .A2(net370),
    .A3(_04013_),
    .B1(_04012_),
    .X(_04117_));
 sky130_fd_sc_hd__and4_1 _12619_ (.A(net552),
    .B(net558),
    .C(net382),
    .D(net375),
    .X(_04118_));
 sky130_fd_sc_hd__a22oi_1 _12620_ (.A1(net552),
    .A2(net382),
    .B1(net375),
    .B2(net558),
    .Y(_04119_));
 sky130_fd_sc_hd__and4bb_1 _12621_ (.A_N(_04118_),
    .B_N(_04119_),
    .C(net565),
    .D(net370),
    .X(_04120_));
 sky130_fd_sc_hd__o2bb2a_1 _12622_ (.A1_N(net565),
    .A2_N(net370),
    .B1(_04118_),
    .B2(_04119_),
    .X(_04121_));
 sky130_fd_sc_hd__a211o_1 _12623_ (.A1(_04028_),
    .A2(_04030_),
    .B1(_04120_),
    .C1(_04121_),
    .X(_04122_));
 sky130_fd_sc_hd__o211ai_1 _12624_ (.A1(_04120_),
    .A2(_04121_),
    .B1(_04028_),
    .C1(_04030_),
    .Y(_04123_));
 sky130_fd_sc_hd__and2_1 _12625_ (.A(_04122_),
    .B(_04123_),
    .X(_04124_));
 sky130_fd_sc_hd__nand2_1 _12626_ (.A(_04117_),
    .B(_04124_),
    .Y(_04125_));
 sky130_fd_sc_hd__xnor2_1 _12627_ (.A(_04117_),
    .B(_04124_),
    .Y(_04126_));
 sky130_fd_sc_hd__a21o_1 _12628_ (.A1(_04016_),
    .A2(_04018_),
    .B1(_04126_),
    .X(_04127_));
 sky130_fd_sc_hd__nand3_1 _12629_ (.A(_04016_),
    .B(_04018_),
    .C(_04126_),
    .Y(_04128_));
 sky130_fd_sc_hd__and3_2 _12630_ (.A(_04116_),
    .B(_04127_),
    .C(_04128_),
    .X(_04129_));
 sky130_fd_sc_hd__inv_2 _12631_ (.A(_04129_),
    .Y(_04130_));
 sky130_fd_sc_hd__a21oi_2 _12632_ (.A1(_04127_),
    .A2(_04128_),
    .B1(_04116_),
    .Y(_04131_));
 sky130_fd_sc_hd__a211o_2 _12633_ (.A1(_04043_),
    .A2(_04046_),
    .B1(_04129_),
    .C1(_04131_),
    .X(_04132_));
 sky130_fd_sc_hd__o211ai_4 _12634_ (.A1(_04129_),
    .A2(_04131_),
    .B1(_04043_),
    .C1(_04046_),
    .Y(_04133_));
 sky130_fd_sc_hd__o211ai_4 _12635_ (.A1(_04020_),
    .A2(_04022_),
    .B1(_04132_),
    .C1(_04133_),
    .Y(_04134_));
 sky130_fd_sc_hd__a211o_1 _12636_ (.A1(_04132_),
    .A2(_04133_),
    .B1(_04020_),
    .C1(_04022_),
    .X(_04135_));
 sky130_fd_sc_hd__nand4_2 _12637_ (.A(net541),
    .B(net544),
    .C(net395),
    .D(net391),
    .Y(_04136_));
 sky130_fd_sc_hd__a22o_1 _12638_ (.A1(net541),
    .A2(net395),
    .B1(net391),
    .B2(net545),
    .X(_04137_));
 sky130_fd_sc_hd__nand4_2 _12639_ (.A(net549),
    .B(net386),
    .C(_04136_),
    .D(_04137_),
    .Y(_04138_));
 sky130_fd_sc_hd__a22o_1 _12640_ (.A1(net548),
    .A2(net389),
    .B1(_04136_),
    .B2(_04137_),
    .X(_04139_));
 sky130_fd_sc_hd__and2_1 _12641_ (.A(_04138_),
    .B(_04139_),
    .X(_04140_));
 sky130_fd_sc_hd__nand2_1 _12642_ (.A(net536),
    .B(net401),
    .Y(_04141_));
 sky130_fd_sc_hd__and4_1 _12643_ (.A(net526),
    .B(net531),
    .C(net409),
    .D(net405),
    .X(_04142_));
 sky130_fd_sc_hd__a22o_1 _12644_ (.A1(net526),
    .A2(net409),
    .B1(net405),
    .B2(net531),
    .X(_04143_));
 sky130_fd_sc_hd__and2b_1 _12645_ (.A_N(_04142_),
    .B(_04143_),
    .X(_04144_));
 sky130_fd_sc_hd__xnor2_2 _12646_ (.A(_04141_),
    .B(_04144_),
    .Y(_04145_));
 sky130_fd_sc_hd__a31o_1 _12647_ (.A1(net541),
    .A2(net401),
    .A3(_04035_),
    .B1(_04034_),
    .X(_04146_));
 sky130_fd_sc_hd__and2_2 _12648_ (.A(_04145_),
    .B(_04146_),
    .X(_04147_));
 sky130_fd_sc_hd__xor2_2 _12649_ (.A(_04145_),
    .B(_04146_),
    .X(_04148_));
 sky130_fd_sc_hd__and2_2 _12650_ (.A(_04140_),
    .B(_04148_),
    .X(_04149_));
 sky130_fd_sc_hd__xnor2_2 _12651_ (.A(_04140_),
    .B(_04148_),
    .Y(_04150_));
 sky130_fd_sc_hd__a21o_4 _12652_ (.A1(_04055_),
    .A2(_04057_),
    .B1(_04150_),
    .X(_04151_));
 sky130_fd_sc_hd__nand3_4 _12653_ (.A(_04055_),
    .B(_04057_),
    .C(_04150_),
    .Y(_04152_));
 sky130_fd_sc_hd__o211a_2 _12654_ (.A1(_04039_),
    .A2(_04041_),
    .B1(_04151_),
    .C1(_04152_),
    .X(_04153_));
 sky130_fd_sc_hd__o211ai_4 _12655_ (.A1(_04039_),
    .A2(_04041_),
    .B1(_04151_),
    .C1(_04152_),
    .Y(_04154_));
 sky130_fd_sc_hd__a211oi_4 _12656_ (.A1(_04151_),
    .A2(_04152_),
    .B1(_04039_),
    .C1(_04041_),
    .Y(_04155_));
 sky130_fd_sc_hd__a31o_1 _12657_ (.A1(net526),
    .A2(net414),
    .A3(_04052_),
    .B1(_04051_),
    .X(_04156_));
 sky130_fd_sc_hd__o21ba_1 _12658_ (.A1(_04059_),
    .A2(_04061_),
    .B1_N(_04060_),
    .X(_04157_));
 sky130_fd_sc_hd__nand2_1 _12659_ (.A(net521),
    .B(net414),
    .Y(_04158_));
 sky130_fd_sc_hd__and3_1 _12660_ (.A(net512),
    .B(net516),
    .C(\mul0.b[7] ),
    .X(_04159_));
 sky130_fd_sc_hd__a22o_1 _12661_ (.A1(net511),
    .A2(net425),
    .B1(\mul0.b[7] ),
    .B2(net516),
    .X(_04160_));
 sky130_fd_sc_hd__a21bo_1 _12662_ (.A1(net422),
    .A2(_04159_),
    .B1_N(_04160_),
    .X(_04161_));
 sky130_fd_sc_hd__xor2_2 _12663_ (.A(_04158_),
    .B(_04161_),
    .X(_04162_));
 sky130_fd_sc_hd__nand2b_2 _12664_ (.A_N(_04157_),
    .B(_04162_),
    .Y(_04163_));
 sky130_fd_sc_hd__xnor2_2 _12665_ (.A(_04157_),
    .B(_04162_),
    .Y(_04164_));
 sky130_fd_sc_hd__nand2_2 _12666_ (.A(_04156_),
    .B(_04164_),
    .Y(_04165_));
 sky130_fd_sc_hd__xor2_2 _12667_ (.A(_04156_),
    .B(_04164_),
    .X(_04166_));
 sky130_fd_sc_hd__a22oi_1 _12668_ (.A1(net503),
    .A2(net432),
    .B1(net498),
    .B2(net437),
    .Y(_04167_));
 sky130_fd_sc_hd__and4_1 _12669_ (.A(net503),
    .B(net437),
    .C(net432),
    .D(net498),
    .X(_04168_));
 sky130_fd_sc_hd__and4bb_1 _12670_ (.A_N(_04167_),
    .B_N(_04168_),
    .C(net507),
    .D(net427),
    .X(_04169_));
 sky130_fd_sc_hd__o2bb2a_1 _12671_ (.A1_N(net507),
    .A2_N(net427),
    .B1(_04167_),
    .B2(_04168_),
    .X(_04170_));
 sky130_fd_sc_hd__nor2_1 _12672_ (.A(_04169_),
    .B(_04170_),
    .Y(_04171_));
 sky130_fd_sc_hd__and2_1 _12673_ (.A(net441),
    .B(net494),
    .X(_04172_));
 sky130_fd_sc_hd__nand4_2 _12674_ (.A(net452),
    .B(net446),
    .C(net490),
    .D(net486),
    .Y(_04173_));
 sky130_fd_sc_hd__a22o_1 _12675_ (.A1(net446),
    .A2(net490),
    .B1(net486),
    .B2(net452),
    .X(_04174_));
 sky130_fd_sc_hd__nand3_1 _12676_ (.A(_04172_),
    .B(_04173_),
    .C(_04174_),
    .Y(_04175_));
 sky130_fd_sc_hd__a21o_1 _12677_ (.A1(_04173_),
    .A2(_04174_),
    .B1(_04172_),
    .X(_04176_));
 sky130_fd_sc_hd__a21bo_1 _12678_ (.A1(_04064_),
    .A2(_04066_),
    .B1_N(_04065_),
    .X(_04177_));
 sky130_fd_sc_hd__nand3_1 _12679_ (.A(_04175_),
    .B(_04176_),
    .C(_04177_),
    .Y(_04178_));
 sky130_fd_sc_hd__a21o_1 _12680_ (.A1(_04175_),
    .A2(_04176_),
    .B1(_04177_),
    .X(_04179_));
 sky130_fd_sc_hd__nand3_2 _12681_ (.A(_04171_),
    .B(_04178_),
    .C(_04179_),
    .Y(_04180_));
 sky130_fd_sc_hd__a21o_1 _12682_ (.A1(_04178_),
    .A2(_04179_),
    .B1(_04171_),
    .X(_04181_));
 sky130_fd_sc_hd__a21bo_1 _12683_ (.A1(_04063_),
    .A2(_04071_),
    .B1_N(_04070_),
    .X(_04182_));
 sky130_fd_sc_hd__nand3_4 _12684_ (.A(_04180_),
    .B(_04181_),
    .C(_04182_),
    .Y(_04183_));
 sky130_fd_sc_hd__a21o_1 _12685_ (.A1(_04180_),
    .A2(_04181_),
    .B1(_04182_),
    .X(_04184_));
 sky130_fd_sc_hd__and3_1 _12686_ (.A(_04166_),
    .B(_04183_),
    .C(_04184_),
    .X(_04185_));
 sky130_fd_sc_hd__nand3_2 _12687_ (.A(_04166_),
    .B(_04183_),
    .C(_04184_),
    .Y(_04186_));
 sky130_fd_sc_hd__a21oi_2 _12688_ (.A1(_04183_),
    .A2(_04184_),
    .B1(_04166_),
    .Y(_04187_));
 sky130_fd_sc_hd__a211oi_4 _12689_ (.A1(_04075_),
    .A2(_04078_),
    .B1(_04185_),
    .C1(_04187_),
    .Y(_04188_));
 sky130_fd_sc_hd__o211a_2 _12690_ (.A1(_04185_),
    .A2(_04187_),
    .B1(_04075_),
    .C1(_04078_),
    .X(_04189_));
 sky130_fd_sc_hd__nor4_2 _12691_ (.A(_04153_),
    .B(_04155_),
    .C(_04188_),
    .D(_04189_),
    .Y(_04190_));
 sky130_fd_sc_hd__or4_2 _12692_ (.A(_04153_),
    .B(_04155_),
    .C(_04188_),
    .D(_04189_),
    .X(_04191_));
 sky130_fd_sc_hd__o22ai_4 _12693_ (.A1(_04153_),
    .A2(_04155_),
    .B1(_04188_),
    .B2(_04189_),
    .Y(_04192_));
 sky130_fd_sc_hd__o211ai_4 _12694_ (.A1(_04080_),
    .A2(_04082_),
    .B1(_04191_),
    .C1(_04192_),
    .Y(_04193_));
 sky130_fd_sc_hd__a211o_2 _12695_ (.A1(_04191_),
    .A2(_04192_),
    .B1(_04080_),
    .C1(_04082_),
    .X(_04194_));
 sky130_fd_sc_hd__and4_1 _12696_ (.A(_04134_),
    .B(_04135_),
    .C(_04193_),
    .D(_04194_),
    .X(_04195_));
 sky130_fd_sc_hd__nand4_2 _12697_ (.A(_04134_),
    .B(_04135_),
    .C(_04193_),
    .D(_04194_),
    .Y(_04196_));
 sky130_fd_sc_hd__a22oi_2 _12698_ (.A1(_04134_),
    .A2(_04135_),
    .B1(_04193_),
    .B2(_04194_),
    .Y(_04197_));
 sky130_fd_sc_hd__a211o_1 _12699_ (.A1(_04085_),
    .A2(_04087_),
    .B1(_04195_),
    .C1(_04197_),
    .X(_04198_));
 sky130_fd_sc_hd__o211ai_2 _12700_ (.A1(_04195_),
    .A2(_04197_),
    .B1(_04085_),
    .C1(_04087_),
    .Y(_04199_));
 sky130_fd_sc_hd__nand3_1 _12701_ (.A(_04105_),
    .B(_04198_),
    .C(_04199_),
    .Y(_04200_));
 sky130_fd_sc_hd__a21o_1 _12702_ (.A1(_04198_),
    .A2(_04199_),
    .B1(_04105_),
    .X(_04201_));
 sky130_fd_sc_hd__o211a_1 _12703_ (.A1(_04089_),
    .A2(_04091_),
    .B1(_04200_),
    .C1(_04201_),
    .X(_04202_));
 sky130_fd_sc_hd__a211o_1 _12704_ (.A1(_04200_),
    .A2(_04201_),
    .B1(_04089_),
    .C1(_04091_),
    .X(_04203_));
 sky130_fd_sc_hd__nand2b_2 _12705_ (.A_N(_04202_),
    .B(_04203_),
    .Y(_04204_));
 sky130_fd_sc_hd__o21ba_1 _12706_ (.A1(_03987_),
    .A2(_04095_),
    .B1_N(_04094_),
    .X(_04205_));
 sky130_fd_sc_hd__xnor2_4 _12707_ (.A(_04204_),
    .B(_04205_),
    .Y(_04206_));
 sky130_fd_sc_hd__or3_1 _12708_ (.A(_03887_),
    .B(_03989_),
    .C(_04096_),
    .X(_04207_));
 sky130_fd_sc_hd__a21boi_4 _12709_ (.A1(_03999_),
    .A2(_04099_),
    .B1_N(_04207_),
    .Y(_04208_));
 sky130_fd_sc_hd__xnor2_4 _12710_ (.A(_04206_),
    .B(_04208_),
    .Y(_04209_));
 sky130_fd_sc_hd__nor2_1 _12711_ (.A(net9),
    .B(_04209_),
    .Y(_04210_));
 sky130_fd_sc_hd__a221o_1 _12712_ (.A1(net599),
    .A2(net706),
    .B1(_02744_),
    .B2(net6),
    .C1(_04210_),
    .X(_04211_));
 sky130_fd_sc_hd__mux2_1 _12713_ (.A0(net849),
    .A1(_04211_),
    .S(net3),
    .X(_00271_));
 sky130_fd_sc_hd__a31oi_2 _12714_ (.A1(net583),
    .A2(net360),
    .A3(_04114_),
    .B1(_04113_),
    .Y(_04212_));
 sky130_fd_sc_hd__a21oi_2 _12715_ (.A1(_04132_),
    .A2(_04134_),
    .B1(_04212_),
    .Y(_04213_));
 sky130_fd_sc_hd__and3_1 _12716_ (.A(_04132_),
    .B(_04134_),
    .C(_04212_),
    .X(_04214_));
 sky130_fd_sc_hd__or2_1 _12717_ (.A(_04213_),
    .B(_04214_),
    .X(_04215_));
 sky130_fd_sc_hd__a22o_1 _12718_ (.A1(net578),
    .A2(net360),
    .B1(net355),
    .B2(net583),
    .X(_04216_));
 sky130_fd_sc_hd__inv_2 _12719_ (.A(_04216_),
    .Y(_04217_));
 sky130_fd_sc_hd__and4_2 _12720_ (.A(net578),
    .B(net583),
    .C(net360),
    .D(net355),
    .X(_04218_));
 sky130_fd_sc_hd__nor2_1 _12721_ (.A(_04217_),
    .B(_04218_),
    .Y(_04219_));
 sky130_fd_sc_hd__and4_1 _12722_ (.A(net562),
    .B(net568),
    .C(net631),
    .D(net365),
    .X(_04220_));
 sky130_fd_sc_hd__inv_2 _12723_ (.A(_04220_),
    .Y(_04221_));
 sky130_fd_sc_hd__a22o_1 _12724_ (.A1(net562),
    .A2(net631),
    .B1(net365),
    .B2(net568),
    .X(_04222_));
 sky130_fd_sc_hd__and4_1 _12725_ (.A(net573),
    .B(net364),
    .C(_04221_),
    .D(_04222_),
    .X(_04223_));
 sky130_fd_sc_hd__a22oi_1 _12726_ (.A1(net573),
    .A2(net364),
    .B1(_04221_),
    .B2(_04222_),
    .Y(_04224_));
 sky130_fd_sc_hd__or2_2 _12727_ (.A(_04223_),
    .B(_04224_),
    .X(_04225_));
 sky130_fd_sc_hd__or2_2 _12728_ (.A(_04106_),
    .B(_04109_),
    .X(_04226_));
 sky130_fd_sc_hd__and2b_1 _12729_ (.A_N(_04225_),
    .B(_04226_),
    .X(_04227_));
 sky130_fd_sc_hd__xor2_4 _12730_ (.A(_04225_),
    .B(_04226_),
    .X(_04228_));
 sky130_fd_sc_hd__xor2_2 _12731_ (.A(_04219_),
    .B(_04228_),
    .X(_04229_));
 sky130_fd_sc_hd__or2_1 _12732_ (.A(_04118_),
    .B(_04120_),
    .X(_04230_));
 sky130_fd_sc_hd__and4_1 _12733_ (.A(net550),
    .B(net554),
    .C(net381),
    .D(net376),
    .X(_04231_));
 sky130_fd_sc_hd__a22oi_1 _12734_ (.A1(net550),
    .A2(net382),
    .B1(net376),
    .B2(net554),
    .Y(_04232_));
 sky130_fd_sc_hd__and4bb_1 _12735_ (.A_N(_04231_),
    .B_N(_04232_),
    .C(net558),
    .D(net370),
    .X(_04233_));
 sky130_fd_sc_hd__o2bb2a_1 _12736_ (.A1_N(net558),
    .A2_N(net370),
    .B1(_04231_),
    .B2(_04232_),
    .X(_04234_));
 sky130_fd_sc_hd__a211o_1 _12737_ (.A1(_04136_),
    .A2(_04138_),
    .B1(_04233_),
    .C1(_04234_),
    .X(_04235_));
 sky130_fd_sc_hd__o211ai_1 _12738_ (.A1(_04233_),
    .A2(_04234_),
    .B1(_04136_),
    .C1(_04138_),
    .Y(_04236_));
 sky130_fd_sc_hd__and2_1 _12739_ (.A(_04235_),
    .B(_04236_),
    .X(_04237_));
 sky130_fd_sc_hd__nand2_1 _12740_ (.A(_04230_),
    .B(_04237_),
    .Y(_04238_));
 sky130_fd_sc_hd__xnor2_2 _12741_ (.A(_04230_),
    .B(_04237_),
    .Y(_04239_));
 sky130_fd_sc_hd__a21oi_4 _12742_ (.A1(_04122_),
    .A2(_04125_),
    .B1(_04239_),
    .Y(_04240_));
 sky130_fd_sc_hd__and3_1 _12743_ (.A(_04122_),
    .B(_04125_),
    .C(_04239_),
    .X(_04241_));
 sky130_fd_sc_hd__nor3_4 _12744_ (.A(_04229_),
    .B(_04240_),
    .C(_04241_),
    .Y(_04242_));
 sky130_fd_sc_hd__o21a_1 _12745_ (.A1(_04240_),
    .A2(_04241_),
    .B1(_04229_),
    .X(_04243_));
 sky130_fd_sc_hd__a211oi_4 _12746_ (.A1(_04151_),
    .A2(_04154_),
    .B1(_04242_),
    .C1(_04243_),
    .Y(_04244_));
 sky130_fd_sc_hd__o211a_1 _12747_ (.A1(_04242_),
    .A2(_04243_),
    .B1(_04151_),
    .C1(_04154_),
    .X(_04245_));
 sky130_fd_sc_hd__a211oi_4 _12748_ (.A1(_04127_),
    .A2(_04130_),
    .B1(_04244_),
    .C1(_04245_),
    .Y(_04246_));
 sky130_fd_sc_hd__o211a_1 _12749_ (.A1(_04244_),
    .A2(_04245_),
    .B1(_04127_),
    .C1(_04130_),
    .X(_04247_));
 sky130_fd_sc_hd__nand2_1 _12750_ (.A(net545),
    .B(net389),
    .Y(_04248_));
 sky130_fd_sc_hd__and3_1 _12751_ (.A(net535),
    .B(net540),
    .C(net391),
    .X(_04249_));
 sky130_fd_sc_hd__a22o_1 _12752_ (.A1(net535),
    .A2(net395),
    .B1(net391),
    .B2(net541),
    .X(_04250_));
 sky130_fd_sc_hd__a21bo_1 _12753_ (.A1(net395),
    .A2(_04249_),
    .B1_N(_04250_),
    .X(_04251_));
 sky130_fd_sc_hd__xor2_2 _12754_ (.A(_04248_),
    .B(_04251_),
    .X(_04252_));
 sky130_fd_sc_hd__nand2_1 _12755_ (.A(net531),
    .B(net401),
    .Y(_04253_));
 sky130_fd_sc_hd__and3_1 _12756_ (.A(net521),
    .B(net526),
    .C(net405),
    .X(_04254_));
 sky130_fd_sc_hd__a22o_1 _12757_ (.A1(net521),
    .A2(net409),
    .B1(net405),
    .B2(net526),
    .X(_04255_));
 sky130_fd_sc_hd__a21bo_1 _12758_ (.A1(net409),
    .A2(_04254_),
    .B1_N(_04255_),
    .X(_04256_));
 sky130_fd_sc_hd__xor2_2 _12759_ (.A(_04253_),
    .B(_04256_),
    .X(_04257_));
 sky130_fd_sc_hd__a31o_1 _12760_ (.A1(net536),
    .A2(net401),
    .A3(_04143_),
    .B1(_04142_),
    .X(_04258_));
 sky130_fd_sc_hd__and2_1 _12761_ (.A(_04257_),
    .B(_04258_),
    .X(_04259_));
 sky130_fd_sc_hd__xor2_2 _12762_ (.A(_04257_),
    .B(_04258_),
    .X(_04260_));
 sky130_fd_sc_hd__and2_1 _12763_ (.A(_04252_),
    .B(_04260_),
    .X(_04261_));
 sky130_fd_sc_hd__xnor2_2 _12764_ (.A(_04252_),
    .B(_04260_),
    .Y(_04262_));
 sky130_fd_sc_hd__a21o_4 _12765_ (.A1(_04163_),
    .A2(_04165_),
    .B1(_04262_),
    .X(_04263_));
 sky130_fd_sc_hd__nand3_4 _12766_ (.A(_04163_),
    .B(_04165_),
    .C(_04262_),
    .Y(_04264_));
 sky130_fd_sc_hd__o211a_1 _12767_ (.A1(_04147_),
    .A2(_04149_),
    .B1(_04263_),
    .C1(_04264_),
    .X(_04265_));
 sky130_fd_sc_hd__o211ai_4 _12768_ (.A1(_04147_),
    .A2(_04149_),
    .B1(_04263_),
    .C1(_04264_),
    .Y(_04266_));
 sky130_fd_sc_hd__a211oi_4 _12769_ (.A1(_04263_),
    .A2(_04264_),
    .B1(_04147_),
    .C1(_04149_),
    .Y(_04267_));
 sky130_fd_sc_hd__a32o_1 _12770_ (.A1(net521),
    .A2(net414),
    .A3(_04160_),
    .B1(_04159_),
    .B2(net425),
    .X(_04268_));
 sky130_fd_sc_hd__nand4_2 _12771_ (.A(net507),
    .B(net512),
    .C(net425),
    .D(\mul0.b[7] ),
    .Y(_04269_));
 sky130_fd_sc_hd__a22o_1 _12772_ (.A1(net507),
    .A2(net425),
    .B1(\mul0.b[7] ),
    .B2(net512),
    .X(_04270_));
 sky130_fd_sc_hd__nand4_2 _12773_ (.A(net516),
    .B(\mul0.b[8] ),
    .C(_04269_),
    .D(_04270_),
    .Y(_04271_));
 sky130_fd_sc_hd__a22o_1 _12774_ (.A1(net516),
    .A2(\mul0.b[8] ),
    .B1(_04269_),
    .B2(_04270_),
    .X(_04272_));
 sky130_fd_sc_hd__o211a_1 _12775_ (.A1(_04168_),
    .A2(_04169_),
    .B1(_04271_),
    .C1(_04272_),
    .X(_04273_));
 sky130_fd_sc_hd__a211o_1 _12776_ (.A1(_04271_),
    .A2(_04272_),
    .B1(_04168_),
    .C1(_04169_),
    .X(_04274_));
 sky130_fd_sc_hd__nand2b_1 _12777_ (.A_N(_04273_),
    .B(_04274_),
    .Y(_04275_));
 sky130_fd_sc_hd__xnor2_2 _12778_ (.A(_04268_),
    .B(_04275_),
    .Y(_04276_));
 sky130_fd_sc_hd__a22oi_1 _12779_ (.A1(net432),
    .A2(net498),
    .B1(net494),
    .B2(net437),
    .Y(_04277_));
 sky130_fd_sc_hd__and4_1 _12780_ (.A(net437),
    .B(net432),
    .C(net498),
    .D(net494),
    .X(_04278_));
 sky130_fd_sc_hd__and4bb_1 _12781_ (.A_N(_04277_),
    .B_N(_04278_),
    .C(net503),
    .D(net427),
    .X(_04279_));
 sky130_fd_sc_hd__o2bb2a_1 _12782_ (.A1_N(net503),
    .A2_N(net427),
    .B1(_04277_),
    .B2(_04278_),
    .X(_04280_));
 sky130_fd_sc_hd__nor2_1 _12783_ (.A(_04279_),
    .B(_04280_),
    .Y(_04281_));
 sky130_fd_sc_hd__and2_1 _12784_ (.A(net441),
    .B(net490),
    .X(_04282_));
 sky130_fd_sc_hd__nand4_2 _12785_ (.A(net452),
    .B(net446),
    .C(net486),
    .D(net482),
    .Y(_04283_));
 sky130_fd_sc_hd__a22o_1 _12786_ (.A1(net446),
    .A2(net486),
    .B1(net482),
    .B2(net452),
    .X(_04284_));
 sky130_fd_sc_hd__nand3_1 _12787_ (.A(_04282_),
    .B(_04283_),
    .C(_04284_),
    .Y(_04285_));
 sky130_fd_sc_hd__a21o_1 _12788_ (.A1(_04283_),
    .A2(_04284_),
    .B1(_04282_),
    .X(_04286_));
 sky130_fd_sc_hd__a21bo_1 _12789_ (.A1(_04172_),
    .A2(_04174_),
    .B1_N(_04173_),
    .X(_04287_));
 sky130_fd_sc_hd__nand3_1 _12790_ (.A(_04285_),
    .B(_04286_),
    .C(_04287_),
    .Y(_04288_));
 sky130_fd_sc_hd__a21o_1 _12791_ (.A1(_04285_),
    .A2(_04286_),
    .B1(_04287_),
    .X(_04289_));
 sky130_fd_sc_hd__nand3_2 _12792_ (.A(_04281_),
    .B(_04288_),
    .C(_04289_),
    .Y(_04290_));
 sky130_fd_sc_hd__a21o_1 _12793_ (.A1(_04288_),
    .A2(_04289_),
    .B1(_04281_),
    .X(_04291_));
 sky130_fd_sc_hd__a21bo_1 _12794_ (.A1(_04171_),
    .A2(_04179_),
    .B1_N(_04178_),
    .X(_04292_));
 sky130_fd_sc_hd__nand3_4 _12795_ (.A(_04290_),
    .B(_04291_),
    .C(_04292_),
    .Y(_04293_));
 sky130_fd_sc_hd__a21o_1 _12796_ (.A1(_04290_),
    .A2(_04291_),
    .B1(_04292_),
    .X(_04294_));
 sky130_fd_sc_hd__and3_1 _12797_ (.A(_04276_),
    .B(_04293_),
    .C(_04294_),
    .X(_04295_));
 sky130_fd_sc_hd__nand3_2 _12798_ (.A(_04276_),
    .B(_04293_),
    .C(_04294_),
    .Y(_04296_));
 sky130_fd_sc_hd__a21oi_2 _12799_ (.A1(_04293_),
    .A2(_04294_),
    .B1(_04276_),
    .Y(_04297_));
 sky130_fd_sc_hd__a211oi_4 _12800_ (.A1(_04183_),
    .A2(_04186_),
    .B1(_04295_),
    .C1(_04297_),
    .Y(_04298_));
 sky130_fd_sc_hd__o211a_2 _12801_ (.A1(_04295_),
    .A2(_04297_),
    .B1(_04183_),
    .C1(_04186_),
    .X(_04299_));
 sky130_fd_sc_hd__nor4_2 _12802_ (.A(_04265_),
    .B(_04267_),
    .C(_04298_),
    .D(_04299_),
    .Y(_04300_));
 sky130_fd_sc_hd__or4_2 _12803_ (.A(_04265_),
    .B(_04267_),
    .C(_04298_),
    .D(_04299_),
    .X(_04301_));
 sky130_fd_sc_hd__o22ai_4 _12804_ (.A1(_04265_),
    .A2(_04267_),
    .B1(_04298_),
    .B2(_04299_),
    .Y(_04302_));
 sky130_fd_sc_hd__o211ai_4 _12805_ (.A1(_04188_),
    .A2(_04190_),
    .B1(_04301_),
    .C1(_04302_),
    .Y(_04303_));
 sky130_fd_sc_hd__a211o_1 _12806_ (.A1(_04301_),
    .A2(_04302_),
    .B1(_04188_),
    .C1(_04190_),
    .X(_04304_));
 sky130_fd_sc_hd__and4bb_2 _12807_ (.A_N(_04246_),
    .B_N(_04247_),
    .C(_04303_),
    .D(_04304_),
    .X(_04305_));
 sky130_fd_sc_hd__or4bb_2 _12808_ (.A(_04246_),
    .B(_04247_),
    .C_N(_04303_),
    .D_N(_04304_),
    .X(_04306_));
 sky130_fd_sc_hd__a2bb2oi_2 _12809_ (.A1_N(_04246_),
    .A2_N(_04247_),
    .B1(_04303_),
    .B2(_04304_),
    .Y(_04307_));
 sky130_fd_sc_hd__a211oi_4 _12810_ (.A1(_04193_),
    .A2(_04196_),
    .B1(_04305_),
    .C1(_04307_),
    .Y(_04308_));
 sky130_fd_sc_hd__o211a_1 _12811_ (.A1(_04305_),
    .A2(_04307_),
    .B1(_04193_),
    .C1(_04196_),
    .X(_04309_));
 sky130_fd_sc_hd__nor3_2 _12812_ (.A(_04215_),
    .B(_04308_),
    .C(_04309_),
    .Y(_04310_));
 sky130_fd_sc_hd__or3_1 _12813_ (.A(_04215_),
    .B(_04308_),
    .C(_04309_),
    .X(_04311_));
 sky130_fd_sc_hd__o21ai_1 _12814_ (.A1(_04308_),
    .A2(_04309_),
    .B1(_04215_),
    .Y(_04312_));
 sky130_fd_sc_hd__a21bo_1 _12815_ (.A1(_04105_),
    .A2(_04199_),
    .B1_N(_04198_),
    .X(_04313_));
 sky130_fd_sc_hd__and3_1 _12816_ (.A(_04311_),
    .B(_04312_),
    .C(_04313_),
    .X(_04314_));
 sky130_fd_sc_hd__a21oi_2 _12817_ (.A1(_04311_),
    .A2(_04312_),
    .B1(_04313_),
    .Y(_04315_));
 sky130_fd_sc_hd__or3_1 _12818_ (.A(_04104_),
    .B(_04314_),
    .C(_04315_),
    .X(_04316_));
 sky130_fd_sc_hd__o21ai_2 _12819_ (.A1(_04314_),
    .A2(_04315_),
    .B1(_04104_),
    .Y(_04317_));
 sky130_fd_sc_hd__nand2_1 _12820_ (.A(_04316_),
    .B(_04317_),
    .Y(_04318_));
 sky130_fd_sc_hd__a21oi_1 _12821_ (.A1(_04094_),
    .A2(_04203_),
    .B1(_04202_),
    .Y(_04319_));
 sky130_fd_sc_hd__and3_1 _12822_ (.A(_04316_),
    .B(_04317_),
    .C(_04319_),
    .X(_04320_));
 sky130_fd_sc_hd__a21oi_1 _12823_ (.A1(_04316_),
    .A2(_04317_),
    .B1(_04319_),
    .Y(_04321_));
 sky130_fd_sc_hd__nor2_2 _12824_ (.A(_04320_),
    .B(_04321_),
    .Y(_04322_));
 sky130_fd_sc_hd__or3_1 _12825_ (.A(_03987_),
    .B(_04096_),
    .C(_04204_),
    .X(_04323_));
 sky130_fd_sc_hd__o21a_2 _12826_ (.A1(_04206_),
    .A2(_04208_),
    .B1(_04323_),
    .X(_04324_));
 sky130_fd_sc_hd__xnor2_4 _12827_ (.A(_04322_),
    .B(_04324_),
    .Y(_04325_));
 sky130_fd_sc_hd__nor2_1 _12828_ (.A(net9),
    .B(_04325_),
    .Y(_04326_));
 sky130_fd_sc_hd__a221o_1 _12829_ (.A1(net599),
    .A2(net809),
    .B1(_02745_),
    .B2(net6),
    .C1(_04326_),
    .X(_04327_));
 sky130_fd_sc_hd__mux2_1 _12830_ (.A0(net873),
    .A1(_04327_),
    .S(_03055_),
    .X(_00272_));
 sky130_fd_sc_hd__and4bb_1 _12831_ (.A_N(_04202_),
    .B_N(_04318_),
    .C(_04203_),
    .D(_04094_),
    .X(_04328_));
 sky130_fd_sc_hd__o21ba_2 _12832_ (.A1(_04322_),
    .A2(_04324_),
    .B1_N(_04328_),
    .X(_04329_));
 sky130_fd_sc_hd__and2_2 _12833_ (.A(_04218_),
    .B(_04227_),
    .X(_04330_));
 sky130_fd_sc_hd__nor2_1 _12834_ (.A(_04218_),
    .B(_04227_),
    .Y(_04331_));
 sky130_fd_sc_hd__o32ai_4 _12835_ (.A1(_04217_),
    .A2(_04218_),
    .A3(_04228_),
    .B1(_04330_),
    .B2(_04331_),
    .Y(_04332_));
 sky130_fd_sc_hd__o21ai_2 _12836_ (.A1(_04244_),
    .A2(_04246_),
    .B1(_04332_),
    .Y(_04333_));
 sky130_fd_sc_hd__or3_1 _12837_ (.A(_04244_),
    .B(_04246_),
    .C(_04332_),
    .X(_04334_));
 sky130_fd_sc_hd__and2_1 _12838_ (.A(_04333_),
    .B(_04334_),
    .X(_04335_));
 sky130_fd_sc_hd__and4_1 _12839_ (.A(net573),
    .B(net578),
    .C(net360),
    .D(net355),
    .X(_04336_));
 sky130_fd_sc_hd__a22o_1 _12840_ (.A1(net573),
    .A2(net360),
    .B1(net355),
    .B2(net578),
    .X(_04337_));
 sky130_fd_sc_hd__inv_2 _12841_ (.A(_04337_),
    .Y(_04338_));
 sky130_fd_sc_hd__and4b_1 _12842_ (.A_N(_04336_),
    .B(_04337_),
    .C(net583),
    .D(net348),
    .X(_04339_));
 sky130_fd_sc_hd__o2bb2a_1 _12843_ (.A1_N(net583),
    .A2_N(net348),
    .B1(_04336_),
    .B2(_04338_),
    .X(_04340_));
 sky130_fd_sc_hd__or2_1 _12844_ (.A(_04339_),
    .B(_04340_),
    .X(_04341_));
 sky130_fd_sc_hd__and4_1 _12845_ (.A(net559),
    .B(net562),
    .C(net631),
    .D(net365),
    .X(_04342_));
 sky130_fd_sc_hd__a22o_1 _12846_ (.A1(net559),
    .A2(net631),
    .B1(net365),
    .B2(net562),
    .X(_04343_));
 sky130_fd_sc_hd__inv_2 _12847_ (.A(_04343_),
    .Y(_04344_));
 sky130_fd_sc_hd__and4b_1 _12848_ (.A_N(_04342_),
    .B(_04343_),
    .C(net568),
    .D(net364),
    .X(_04345_));
 sky130_fd_sc_hd__o2bb2a_1 _12849_ (.A1_N(net568),
    .A2_N(net364),
    .B1(_04342_),
    .B2(_04344_),
    .X(_04346_));
 sky130_fd_sc_hd__or2_1 _12850_ (.A(_04345_),
    .B(_04346_),
    .X(_04347_));
 sky130_fd_sc_hd__or2_1 _12851_ (.A(_04220_),
    .B(_04223_),
    .X(_04348_));
 sky130_fd_sc_hd__nand2b_1 _12852_ (.A_N(_04347_),
    .B(_04348_),
    .Y(_04349_));
 sky130_fd_sc_hd__xor2_2 _12853_ (.A(_04347_),
    .B(_04348_),
    .X(_04350_));
 sky130_fd_sc_hd__or2_1 _12854_ (.A(_04341_),
    .B(_04350_),
    .X(_04351_));
 sky130_fd_sc_hd__xor2_2 _12855_ (.A(_04341_),
    .B(_04350_),
    .X(_04352_));
 sky130_fd_sc_hd__or2_1 _12856_ (.A(_04231_),
    .B(_04233_),
    .X(_04353_));
 sky130_fd_sc_hd__a32o_1 _12857_ (.A1(net546),
    .A2(net389),
    .A3(_04250_),
    .B1(_04249_),
    .B2(net395),
    .X(_04354_));
 sky130_fd_sc_hd__nand4_2 _12858_ (.A(net546),
    .B(net550),
    .C(net381),
    .D(net376),
    .Y(_04355_));
 sky130_fd_sc_hd__a22o_1 _12859_ (.A1(net546),
    .A2(net382),
    .B1(net376),
    .B2(net550),
    .X(_04356_));
 sky130_fd_sc_hd__nand4_2 _12860_ (.A(net554),
    .B(net370),
    .C(_04355_),
    .D(_04356_),
    .Y(_04357_));
 sky130_fd_sc_hd__a22o_1 _12861_ (.A1(net554),
    .A2(net371),
    .B1(_04355_),
    .B2(_04356_),
    .X(_04358_));
 sky130_fd_sc_hd__and3_1 _12862_ (.A(_04354_),
    .B(_04357_),
    .C(_04358_),
    .X(_04359_));
 sky130_fd_sc_hd__a21o_1 _12863_ (.A1(_04357_),
    .A2(_04358_),
    .B1(_04354_),
    .X(_04360_));
 sky130_fd_sc_hd__and2b_1 _12864_ (.A_N(_04359_),
    .B(_04360_),
    .X(_04361_));
 sky130_fd_sc_hd__xnor2_2 _12865_ (.A(_04353_),
    .B(_04361_),
    .Y(_04362_));
 sky130_fd_sc_hd__a21oi_1 _12866_ (.A1(_04235_),
    .A2(_04238_),
    .B1(_04362_),
    .Y(_04363_));
 sky130_fd_sc_hd__a21o_1 _12867_ (.A1(_04235_),
    .A2(_04238_),
    .B1(_04362_),
    .X(_04364_));
 sky130_fd_sc_hd__nand3_1 _12868_ (.A(_04235_),
    .B(_04238_),
    .C(_04362_),
    .Y(_04365_));
 sky130_fd_sc_hd__and3_2 _12869_ (.A(_04352_),
    .B(_04364_),
    .C(_04365_),
    .X(_04366_));
 sky130_fd_sc_hd__a21oi_2 _12870_ (.A1(_04364_),
    .A2(_04365_),
    .B1(_04352_),
    .Y(_04367_));
 sky130_fd_sc_hd__a211o_2 _12871_ (.A1(_04263_),
    .A2(_04266_),
    .B1(_04366_),
    .C1(_04367_),
    .X(_04368_));
 sky130_fd_sc_hd__o211ai_4 _12872_ (.A1(_04366_),
    .A2(_04367_),
    .B1(_04263_),
    .C1(_04266_),
    .Y(_04369_));
 sky130_fd_sc_hd__o211ai_4 _12873_ (.A1(_04240_),
    .A2(_04242_),
    .B1(_04368_),
    .C1(_04369_),
    .Y(_04370_));
 sky130_fd_sc_hd__a211o_1 _12874_ (.A1(_04368_),
    .A2(_04369_),
    .B1(_04240_),
    .C1(_04242_),
    .X(_04371_));
 sky130_fd_sc_hd__a21o_1 _12875_ (.A1(_04268_),
    .A2(_04274_),
    .B1(_04273_),
    .X(_04372_));
 sky130_fd_sc_hd__nand2_1 _12876_ (.A(net542),
    .B(net386),
    .Y(_04373_));
 sky130_fd_sc_hd__and3_1 _12877_ (.A(net531),
    .B(net535),
    .C(net391),
    .X(_04374_));
 sky130_fd_sc_hd__a22o_1 _12878_ (.A1(net531),
    .A2(net395),
    .B1(net391),
    .B2(net535),
    .X(_04375_));
 sky130_fd_sc_hd__a21bo_1 _12879_ (.A1(net395),
    .A2(_04374_),
    .B1_N(_04375_),
    .X(_04376_));
 sky130_fd_sc_hd__xor2_1 _12880_ (.A(_04373_),
    .B(_04376_),
    .X(_04377_));
 sky130_fd_sc_hd__and2_1 _12881_ (.A(net526),
    .B(net401),
    .X(_04378_));
 sky130_fd_sc_hd__nand4_2 _12882_ (.A(net515),
    .B(net521),
    .C(net409),
    .D(net405),
    .Y(_04379_));
 sky130_fd_sc_hd__a22o_1 _12883_ (.A1(net515),
    .A2(net409),
    .B1(net405),
    .B2(net521),
    .X(_04380_));
 sky130_fd_sc_hd__nand3_1 _12884_ (.A(_04378_),
    .B(_04379_),
    .C(_04380_),
    .Y(_04381_));
 sky130_fd_sc_hd__a21o_1 _12885_ (.A1(_04379_),
    .A2(_04380_),
    .B1(_04378_),
    .X(_04382_));
 sky130_fd_sc_hd__a32o_1 _12886_ (.A1(net531),
    .A2(net401),
    .A3(_04255_),
    .B1(_04254_),
    .B2(net409),
    .X(_04383_));
 sky130_fd_sc_hd__nand3_1 _12887_ (.A(_04381_),
    .B(_04382_),
    .C(_04383_),
    .Y(_04384_));
 sky130_fd_sc_hd__a21o_1 _12888_ (.A1(_04381_),
    .A2(_04382_),
    .B1(_04383_),
    .X(_04385_));
 sky130_fd_sc_hd__nand3_2 _12889_ (.A(_04377_),
    .B(_04384_),
    .C(_04385_),
    .Y(_04386_));
 sky130_fd_sc_hd__a21o_1 _12890_ (.A1(_04384_),
    .A2(_04385_),
    .B1(_04377_),
    .X(_04387_));
 sky130_fd_sc_hd__nand3_2 _12891_ (.A(_04372_),
    .B(_04386_),
    .C(_04387_),
    .Y(_04388_));
 sky130_fd_sc_hd__a21o_1 _12892_ (.A1(_04386_),
    .A2(_04387_),
    .B1(_04372_),
    .X(_04389_));
 sky130_fd_sc_hd__o211ai_2 _12893_ (.A1(_04259_),
    .A2(_04261_),
    .B1(_04388_),
    .C1(_04389_),
    .Y(_04390_));
 sky130_fd_sc_hd__a211o_1 _12894_ (.A1(_04388_),
    .A2(_04389_),
    .B1(_04259_),
    .C1(_04261_),
    .X(_04391_));
 sky130_fd_sc_hd__nand2_1 _12895_ (.A(_04390_),
    .B(_04391_),
    .Y(_04392_));
 sky130_fd_sc_hd__nand2_1 _12896_ (.A(_04269_),
    .B(_04271_),
    .Y(_04393_));
 sky130_fd_sc_hd__nand4_2 _12897_ (.A(\mul0.a[17] ),
    .B(net508),
    .C(net422),
    .D(net418),
    .Y(_04394_));
 sky130_fd_sc_hd__a22o_1 _12898_ (.A1(\mul0.a[17] ),
    .A2(net422),
    .B1(net418),
    .B2(net508),
    .X(_04395_));
 sky130_fd_sc_hd__nand4_1 _12899_ (.A(net512),
    .B(net414),
    .C(_04394_),
    .D(_04395_),
    .Y(_04396_));
 sky130_fd_sc_hd__a22o_1 _12900_ (.A1(net512),
    .A2(net414),
    .B1(_04394_),
    .B2(_04395_),
    .X(_04397_));
 sky130_fd_sc_hd__o211a_1 _12901_ (.A1(_04278_),
    .A2(_04279_),
    .B1(_04396_),
    .C1(_04397_),
    .X(_04398_));
 sky130_fd_sc_hd__a211o_1 _12902_ (.A1(_04396_),
    .A2(_04397_),
    .B1(_04278_),
    .C1(_04279_),
    .X(_04399_));
 sky130_fd_sc_hd__nand2b_1 _12903_ (.A_N(_04398_),
    .B(_04399_),
    .Y(_04400_));
 sky130_fd_sc_hd__xnor2_2 _12904_ (.A(_04393_),
    .B(_04400_),
    .Y(_04401_));
 sky130_fd_sc_hd__nand2_1 _12905_ (.A(net429),
    .B(net498),
    .Y(_04402_));
 sky130_fd_sc_hd__a22o_1 _12906_ (.A1(net434),
    .A2(net494),
    .B1(net490),
    .B2(net439),
    .X(_04403_));
 sky130_fd_sc_hd__and3_1 _12907_ (.A(net439),
    .B(net434),
    .C(net494),
    .X(_04404_));
 sky130_fd_sc_hd__a21bo_1 _12908_ (.A1(net490),
    .A2(_04404_),
    .B1_N(_04403_),
    .X(_04405_));
 sky130_fd_sc_hd__xor2_2 _12909_ (.A(_04402_),
    .B(_04405_),
    .X(_04406_));
 sky130_fd_sc_hd__and2_1 _12910_ (.A(net442),
    .B(net486),
    .X(_04407_));
 sky130_fd_sc_hd__nand4_1 _12911_ (.A(net451),
    .B(net447),
    .C(net482),
    .D(net478),
    .Y(_04408_));
 sky130_fd_sc_hd__a22o_1 _12912_ (.A1(net447),
    .A2(net482),
    .B1(net478),
    .B2(net451),
    .X(_04409_));
 sky130_fd_sc_hd__nand3_1 _12913_ (.A(_04407_),
    .B(_04408_),
    .C(_04409_),
    .Y(_04410_));
 sky130_fd_sc_hd__a21o_1 _12914_ (.A1(_04408_),
    .A2(_04409_),
    .B1(_04407_),
    .X(_04411_));
 sky130_fd_sc_hd__a21bo_1 _12915_ (.A1(_04282_),
    .A2(_04284_),
    .B1_N(_04283_),
    .X(_04412_));
 sky130_fd_sc_hd__nand3_1 _12916_ (.A(_04410_),
    .B(_04411_),
    .C(_04412_),
    .Y(_04413_));
 sky130_fd_sc_hd__a21o_1 _12917_ (.A1(_04410_),
    .A2(_04411_),
    .B1(_04412_),
    .X(_04414_));
 sky130_fd_sc_hd__nand3_2 _12918_ (.A(_04406_),
    .B(_04413_),
    .C(_04414_),
    .Y(_04415_));
 sky130_fd_sc_hd__a21o_1 _12919_ (.A1(_04413_),
    .A2(_04414_),
    .B1(_04406_),
    .X(_04416_));
 sky130_fd_sc_hd__a21bo_1 _12920_ (.A1(_04281_),
    .A2(_04289_),
    .B1_N(_04288_),
    .X(_04417_));
 sky130_fd_sc_hd__nand3_4 _12921_ (.A(_04415_),
    .B(_04416_),
    .C(_04417_),
    .Y(_04418_));
 sky130_fd_sc_hd__a21o_1 _12922_ (.A1(_04415_),
    .A2(_04416_),
    .B1(_04417_),
    .X(_04419_));
 sky130_fd_sc_hd__and3_1 _12923_ (.A(_04401_),
    .B(_04418_),
    .C(_04419_),
    .X(_04420_));
 sky130_fd_sc_hd__nand3_2 _12924_ (.A(_04401_),
    .B(_04418_),
    .C(_04419_),
    .Y(_04421_));
 sky130_fd_sc_hd__a21oi_2 _12925_ (.A1(_04418_),
    .A2(_04419_),
    .B1(_04401_),
    .Y(_04422_));
 sky130_fd_sc_hd__a211oi_4 _12926_ (.A1(_04293_),
    .A2(_04296_),
    .B1(_04420_),
    .C1(_04422_),
    .Y(_04423_));
 sky130_fd_sc_hd__o211a_1 _12927_ (.A1(_04420_),
    .A2(_04422_),
    .B1(_04293_),
    .C1(_04296_),
    .X(_04424_));
 sky130_fd_sc_hd__nor3_1 _12928_ (.A(_04392_),
    .B(_04423_),
    .C(_04424_),
    .Y(_04425_));
 sky130_fd_sc_hd__or3_2 _12929_ (.A(_04392_),
    .B(_04423_),
    .C(_04424_),
    .X(_04426_));
 sky130_fd_sc_hd__o21ai_2 _12930_ (.A1(_04423_),
    .A2(_04424_),
    .B1(_04392_),
    .Y(_04427_));
 sky130_fd_sc_hd__o211a_1 _12931_ (.A1(_04298_),
    .A2(_04300_),
    .B1(_04426_),
    .C1(_04427_),
    .X(_04428_));
 sky130_fd_sc_hd__o211ai_4 _12932_ (.A1(_04298_),
    .A2(_04300_),
    .B1(_04426_),
    .C1(_04427_),
    .Y(_04429_));
 sky130_fd_sc_hd__a211o_1 _12933_ (.A1(_04426_),
    .A2(_04427_),
    .B1(_04298_),
    .C1(_04300_),
    .X(_04430_));
 sky130_fd_sc_hd__and4_2 _12934_ (.A(_04370_),
    .B(_04371_),
    .C(_04429_),
    .D(_04430_),
    .X(_04431_));
 sky130_fd_sc_hd__a22oi_4 _12935_ (.A1(_04370_),
    .A2(_04371_),
    .B1(_04429_),
    .B2(_04430_),
    .Y(_04432_));
 sky130_fd_sc_hd__a211o_2 _12936_ (.A1(_04303_),
    .A2(_04306_),
    .B1(_04431_),
    .C1(_04432_),
    .X(_04433_));
 sky130_fd_sc_hd__o211ai_4 _12937_ (.A1(_04431_),
    .A2(_04432_),
    .B1(_04303_),
    .C1(_04306_),
    .Y(_04434_));
 sky130_fd_sc_hd__nand3_4 _12938_ (.A(_04335_),
    .B(_04433_),
    .C(_04434_),
    .Y(_04435_));
 sky130_fd_sc_hd__a21o_1 _12939_ (.A1(_04433_),
    .A2(_04434_),
    .B1(_04335_),
    .X(_04436_));
 sky130_fd_sc_hd__o211ai_4 _12940_ (.A1(_04308_),
    .A2(_04310_),
    .B1(_04435_),
    .C1(_04436_),
    .Y(_04437_));
 sky130_fd_sc_hd__a211o_1 _12941_ (.A1(_04435_),
    .A2(_04436_),
    .B1(_04308_),
    .C1(_04310_),
    .X(_04438_));
 sky130_fd_sc_hd__nand3_4 _12942_ (.A(_04213_),
    .B(_04437_),
    .C(_04438_),
    .Y(_04439_));
 sky130_fd_sc_hd__a21o_1 _12943_ (.A1(_04437_),
    .A2(_04438_),
    .B1(_04213_),
    .X(_04440_));
 sky130_fd_sc_hd__o21bai_2 _12944_ (.A1(_04104_),
    .A2(_04315_),
    .B1_N(_04314_),
    .Y(_04441_));
 sky130_fd_sc_hd__nand3_4 _12945_ (.A(_04439_),
    .B(_04440_),
    .C(_04441_),
    .Y(_04442_));
 sky130_fd_sc_hd__a21o_1 _12946_ (.A1(_04439_),
    .A2(_04440_),
    .B1(_04441_),
    .X(_04443_));
 sky130_fd_sc_hd__and3_1 _12947_ (.A(_04202_),
    .B(_04316_),
    .C(_04317_),
    .X(_04444_));
 sky130_fd_sc_hd__a21oi_1 _12948_ (.A1(_04442_),
    .A2(_04443_),
    .B1(_04444_),
    .Y(_04445_));
 sky130_fd_sc_hd__a21o_1 _12949_ (.A1(_04442_),
    .A2(_04443_),
    .B1(_04444_),
    .X(_04446_));
 sky130_fd_sc_hd__and3_1 _12950_ (.A(_04442_),
    .B(_04443_),
    .C(_04444_),
    .X(_04447_));
 sky130_fd_sc_hd__nor2_2 _12951_ (.A(_04445_),
    .B(_04447_),
    .Y(_04448_));
 sky130_fd_sc_hd__xor2_4 _12952_ (.A(_04329_),
    .B(_04448_),
    .X(_04449_));
 sky130_fd_sc_hd__nor2_1 _12953_ (.A(net9),
    .B(_04449_),
    .Y(_04450_));
 sky130_fd_sc_hd__a221o_1 _12954_ (.A1(net599),
    .A2(net742),
    .B1(_02746_),
    .B2(net6),
    .C1(_04450_),
    .X(_04451_));
 sky130_fd_sc_hd__mux2_1 _12955_ (.A0(net867),
    .A1(_04451_),
    .S(net3),
    .X(_00273_));
 sky130_fd_sc_hd__o211a_1 _12956_ (.A1(_04320_),
    .A2(_04321_),
    .B1(_04442_),
    .C1(_04443_),
    .X(_04452_));
 sky130_fd_sc_hd__nor2_1 _12957_ (.A(_04098_),
    .B(_04206_),
    .Y(_04453_));
 sky130_fd_sc_hd__o21ai_1 _12958_ (.A1(_04206_),
    .A2(_04207_),
    .B1(_04323_),
    .Y(_04454_));
 sky130_fd_sc_hd__a221o_1 _12959_ (.A1(_04328_),
    .A2(_04446_),
    .B1(_04452_),
    .B2(_04454_),
    .C1(_04447_),
    .X(_04455_));
 sky130_fd_sc_hd__a31o_4 _12960_ (.A1(_03999_),
    .A2(_04452_),
    .A3(_04453_),
    .B1(_04455_),
    .X(_04456_));
 sky130_fd_sc_hd__nand2_2 _12961_ (.A(_04437_),
    .B(_04439_),
    .Y(_04457_));
 sky130_fd_sc_hd__o211a_1 _12962_ (.A1(_04336_),
    .A2(_04339_),
    .B1(net583),
    .C1(net344),
    .X(_04458_));
 sky130_fd_sc_hd__a211oi_1 _12963_ (.A1(net583),
    .A2(net344),
    .B1(_04336_),
    .C1(_04339_),
    .Y(_04459_));
 sky130_fd_sc_hd__or2_1 _12964_ (.A(_04458_),
    .B(_04459_),
    .X(_04460_));
 sky130_fd_sc_hd__a21oi_1 _12965_ (.A1(_04349_),
    .A2(_04351_),
    .B1(_04460_),
    .Y(_04461_));
 sky130_fd_sc_hd__and3_1 _12966_ (.A(_04349_),
    .B(_04351_),
    .C(_04460_),
    .X(_04462_));
 sky130_fd_sc_hd__nor2_1 _12967_ (.A(_04461_),
    .B(_04462_),
    .Y(_04463_));
 sky130_fd_sc_hd__nand2_1 _12968_ (.A(_04330_),
    .B(_04463_),
    .Y(_04464_));
 sky130_fd_sc_hd__xnor2_1 _12969_ (.A(_04330_),
    .B(_04463_),
    .Y(_04465_));
 sky130_fd_sc_hd__a21oi_2 _12970_ (.A1(_04368_),
    .A2(_04370_),
    .B1(_04465_),
    .Y(_04466_));
 sky130_fd_sc_hd__and3_1 _12971_ (.A(_04368_),
    .B(_04370_),
    .C(_04465_),
    .X(_04467_));
 sky130_fd_sc_hd__nor2_1 _12972_ (.A(_04466_),
    .B(_04467_),
    .Y(_04468_));
 sky130_fd_sc_hd__and4_1 _12973_ (.A(net569),
    .B(net573),
    .C(net360),
    .D(net355),
    .X(_04469_));
 sky130_fd_sc_hd__inv_2 _12974_ (.A(_04469_),
    .Y(_04470_));
 sky130_fd_sc_hd__a22o_1 _12975_ (.A1(net568),
    .A2(net360),
    .B1(net355),
    .B2(net573),
    .X(_04471_));
 sky130_fd_sc_hd__and4_1 _12976_ (.A(net580),
    .B(net348),
    .C(_04470_),
    .D(_04471_),
    .X(_04472_));
 sky130_fd_sc_hd__a22oi_1 _12977_ (.A1(net579),
    .A2(net348),
    .B1(_04470_),
    .B2(_04471_),
    .Y(_04473_));
 sky130_fd_sc_hd__or2_1 _12978_ (.A(_04472_),
    .B(_04473_),
    .X(_04474_));
 sky130_fd_sc_hd__nand2_1 _12979_ (.A(net562),
    .B(net364),
    .Y(_04475_));
 sky130_fd_sc_hd__and4_1 _12980_ (.A(net555),
    .B(net559),
    .C(net631),
    .D(net365),
    .X(_04476_));
 sky130_fd_sc_hd__a22o_1 _12981_ (.A1(net555),
    .A2(net631),
    .B1(net365),
    .B2(net559),
    .X(_04477_));
 sky130_fd_sc_hd__and2b_1 _12982_ (.A_N(_04476_),
    .B(_04477_),
    .X(_04478_));
 sky130_fd_sc_hd__xnor2_1 _12983_ (.A(_04475_),
    .B(_04478_),
    .Y(_04479_));
 sky130_fd_sc_hd__nor2_1 _12984_ (.A(_04342_),
    .B(_04345_),
    .Y(_04480_));
 sky130_fd_sc_hd__nand2b_1 _12985_ (.A_N(_04480_),
    .B(_04479_),
    .Y(_04481_));
 sky130_fd_sc_hd__xnor2_1 _12986_ (.A(_04479_),
    .B(_04480_),
    .Y(_04482_));
 sky130_fd_sc_hd__nand2b_1 _12987_ (.A_N(_04474_),
    .B(_04482_),
    .Y(_04483_));
 sky130_fd_sc_hd__xnor2_1 _12988_ (.A(_04474_),
    .B(_04482_),
    .Y(_04484_));
 sky130_fd_sc_hd__nand2_1 _12989_ (.A(_04355_),
    .B(_04357_),
    .Y(_04485_));
 sky130_fd_sc_hd__a32o_1 _12990_ (.A1(net542),
    .A2(net386),
    .A3(_04375_),
    .B1(_04374_),
    .B2(net395),
    .X(_04486_));
 sky130_fd_sc_hd__nand4_2 _12991_ (.A(net542),
    .B(net546),
    .C(net382),
    .D(net375),
    .Y(_04487_));
 sky130_fd_sc_hd__a22o_1 _12992_ (.A1(\mul0.a[9] ),
    .A2(net382),
    .B1(net376),
    .B2(net546),
    .X(_04488_));
 sky130_fd_sc_hd__nand4_2 _12993_ (.A(net550),
    .B(net370),
    .C(_04487_),
    .D(_04488_),
    .Y(_04489_));
 sky130_fd_sc_hd__a22o_1 _12994_ (.A1(net550),
    .A2(net370),
    .B1(_04487_),
    .B2(_04488_),
    .X(_04490_));
 sky130_fd_sc_hd__nand3_1 _12995_ (.A(_04486_),
    .B(_04489_),
    .C(_04490_),
    .Y(_04491_));
 sky130_fd_sc_hd__a21o_1 _12996_ (.A1(_04489_),
    .A2(_04490_),
    .B1(_04486_),
    .X(_04492_));
 sky130_fd_sc_hd__nand3_1 _12997_ (.A(_04485_),
    .B(_04491_),
    .C(_04492_),
    .Y(_04493_));
 sky130_fd_sc_hd__a21o_1 _12998_ (.A1(_04491_),
    .A2(_04492_),
    .B1(_04485_),
    .X(_04494_));
 sky130_fd_sc_hd__a21o_1 _12999_ (.A1(_04353_),
    .A2(_04360_),
    .B1(_04359_),
    .X(_04495_));
 sky130_fd_sc_hd__nand3_2 _13000_ (.A(_04493_),
    .B(_04494_),
    .C(_04495_),
    .Y(_04496_));
 sky130_fd_sc_hd__a21o_1 _13001_ (.A1(_04493_),
    .A2(_04494_),
    .B1(_04495_),
    .X(_04497_));
 sky130_fd_sc_hd__and3_1 _13002_ (.A(_04484_),
    .B(_04496_),
    .C(_04497_),
    .X(_04498_));
 sky130_fd_sc_hd__inv_2 _13003_ (.A(_04498_),
    .Y(_04499_));
 sky130_fd_sc_hd__a21oi_1 _13004_ (.A1(_04496_),
    .A2(_04497_),
    .B1(_04484_),
    .Y(_04500_));
 sky130_fd_sc_hd__a211o_1 _13005_ (.A1(_04388_),
    .A2(_04390_),
    .B1(_04498_),
    .C1(_04500_),
    .X(_04501_));
 sky130_fd_sc_hd__o211ai_1 _13006_ (.A1(_04498_),
    .A2(_04500_),
    .B1(_04388_),
    .C1(_04390_),
    .Y(_04502_));
 sky130_fd_sc_hd__o211ai_1 _13007_ (.A1(_04363_),
    .A2(_04366_),
    .B1(_04501_),
    .C1(_04502_),
    .Y(_04503_));
 sky130_fd_sc_hd__a211o_1 _13008_ (.A1(_04501_),
    .A2(_04502_),
    .B1(_04363_),
    .C1(_04366_),
    .X(_04504_));
 sky130_fd_sc_hd__nand2_1 _13009_ (.A(_04503_),
    .B(_04504_),
    .Y(_04505_));
 sky130_fd_sc_hd__nand2_1 _13010_ (.A(_04384_),
    .B(_04386_),
    .Y(_04506_));
 sky130_fd_sc_hd__a21o_1 _13011_ (.A1(_04393_),
    .A2(_04399_),
    .B1(_04398_),
    .X(_04507_));
 sky130_fd_sc_hd__nand2_1 _13012_ (.A(net537),
    .B(net386),
    .Y(_04508_));
 sky130_fd_sc_hd__and3_1 _13013_ (.A(net526),
    .B(net532),
    .C(net391),
    .X(_04509_));
 sky130_fd_sc_hd__a22o_1 _13014_ (.A1(net525),
    .A2(net395),
    .B1(net391),
    .B2(net532),
    .X(_04510_));
 sky130_fd_sc_hd__a21bo_1 _13015_ (.A1(net395),
    .A2(_04509_),
    .B1_N(_04510_),
    .X(_04511_));
 sky130_fd_sc_hd__xor2_1 _13016_ (.A(_04508_),
    .B(_04511_),
    .X(_04512_));
 sky130_fd_sc_hd__and2_1 _13017_ (.A(net520),
    .B(net401),
    .X(_04513_));
 sky130_fd_sc_hd__nand4_1 _13018_ (.A(net511),
    .B(net516),
    .C(net409),
    .D(\mul0.b[10] ),
    .Y(_04514_));
 sky130_fd_sc_hd__a22o_1 _13019_ (.A1(net511),
    .A2(net409),
    .B1(\mul0.b[10] ),
    .B2(net516),
    .X(_04515_));
 sky130_fd_sc_hd__nand3_1 _13020_ (.A(_04513_),
    .B(_04514_),
    .C(_04515_),
    .Y(_04516_));
 sky130_fd_sc_hd__a21o_1 _13021_ (.A1(_04514_),
    .A2(_04515_),
    .B1(_04513_),
    .X(_04517_));
 sky130_fd_sc_hd__a21bo_1 _13022_ (.A1(_04378_),
    .A2(_04380_),
    .B1_N(_04379_),
    .X(_04518_));
 sky130_fd_sc_hd__nand3_2 _13023_ (.A(_04516_),
    .B(_04517_),
    .C(_04518_),
    .Y(_04519_));
 sky130_fd_sc_hd__a21o_1 _13024_ (.A1(_04516_),
    .A2(_04517_),
    .B1(_04518_),
    .X(_04520_));
 sky130_fd_sc_hd__nand3_2 _13025_ (.A(_04512_),
    .B(_04519_),
    .C(_04520_),
    .Y(_04521_));
 sky130_fd_sc_hd__a21o_1 _13026_ (.A1(_04519_),
    .A2(_04520_),
    .B1(_04512_),
    .X(_04522_));
 sky130_fd_sc_hd__nand3_4 _13027_ (.A(_04507_),
    .B(_04521_),
    .C(_04522_),
    .Y(_04523_));
 sky130_fd_sc_hd__a21o_1 _13028_ (.A1(_04521_),
    .A2(_04522_),
    .B1(_04507_),
    .X(_04524_));
 sky130_fd_sc_hd__nand3_2 _13029_ (.A(_04506_),
    .B(_04523_),
    .C(_04524_),
    .Y(_04525_));
 sky130_fd_sc_hd__a21o_1 _13030_ (.A1(_04523_),
    .A2(_04524_),
    .B1(_04506_),
    .X(_04526_));
 sky130_fd_sc_hd__nand2_1 _13031_ (.A(_04525_),
    .B(_04526_),
    .Y(_04527_));
 sky130_fd_sc_hd__nand2_1 _13032_ (.A(_04394_),
    .B(_04396_),
    .Y(_04528_));
 sky130_fd_sc_hd__a32o_1 _13033_ (.A1(net429),
    .A2(net498),
    .A3(_04403_),
    .B1(_04404_),
    .B2(net490),
    .X(_04529_));
 sky130_fd_sc_hd__nand4_2 _13034_ (.A(net503),
    .B(net424),
    .C(net420),
    .D(net498),
    .Y(_04530_));
 sky130_fd_sc_hd__a22o_1 _13035_ (.A1(net503),
    .A2(net420),
    .B1(net498),
    .B2(net424),
    .X(_04531_));
 sky130_fd_sc_hd__nand4_2 _13036_ (.A(net508),
    .B(net416),
    .C(_04530_),
    .D(_04531_),
    .Y(_04532_));
 sky130_fd_sc_hd__a22o_1 _13037_ (.A1(net508),
    .A2(net416),
    .B1(_04530_),
    .B2(_04531_),
    .X(_04533_));
 sky130_fd_sc_hd__nand3_1 _13038_ (.A(_04529_),
    .B(_04532_),
    .C(_04533_),
    .Y(_04534_));
 sky130_fd_sc_hd__a21o_1 _13039_ (.A1(_04532_),
    .A2(_04533_),
    .B1(_04529_),
    .X(_04535_));
 sky130_fd_sc_hd__and3_1 _13040_ (.A(_04528_),
    .B(_04534_),
    .C(_04535_),
    .X(_04536_));
 sky130_fd_sc_hd__a21oi_1 _13041_ (.A1(_04534_),
    .A2(_04535_),
    .B1(_04528_),
    .Y(_04537_));
 sky130_fd_sc_hd__nor2_1 _13042_ (.A(_04536_),
    .B(_04537_),
    .Y(_04538_));
 sky130_fd_sc_hd__nand2_1 _13043_ (.A(net429),
    .B(net494),
    .Y(_04539_));
 sky130_fd_sc_hd__and4_1 _13044_ (.A(net439),
    .B(net434),
    .C(net490),
    .D(net486),
    .X(_04540_));
 sky130_fd_sc_hd__a22oi_2 _13045_ (.A1(net434),
    .A2(net490),
    .B1(net486),
    .B2(net439),
    .Y(_04541_));
 sky130_fd_sc_hd__nor2_1 _13046_ (.A(_04540_),
    .B(_04541_),
    .Y(_04542_));
 sky130_fd_sc_hd__xnor2_2 _13047_ (.A(_04539_),
    .B(_04542_),
    .Y(_04543_));
 sky130_fd_sc_hd__and2_1 _13048_ (.A(net442),
    .B(net482),
    .X(_04544_));
 sky130_fd_sc_hd__nand4_1 _13049_ (.A(net451),
    .B(net447),
    .C(net478),
    .D(net474),
    .Y(_04545_));
 sky130_fd_sc_hd__a22o_1 _13050_ (.A1(net447),
    .A2(net478),
    .B1(net474),
    .B2(net451),
    .X(_04546_));
 sky130_fd_sc_hd__nand3_1 _13051_ (.A(_04544_),
    .B(_04545_),
    .C(_04546_),
    .Y(_04547_));
 sky130_fd_sc_hd__a21o_1 _13052_ (.A1(_04545_),
    .A2(_04546_),
    .B1(_04544_),
    .X(_04548_));
 sky130_fd_sc_hd__a21bo_1 _13053_ (.A1(_04407_),
    .A2(_04409_),
    .B1_N(_04408_),
    .X(_04549_));
 sky130_fd_sc_hd__nand3_1 _13054_ (.A(_04547_),
    .B(_04548_),
    .C(_04549_),
    .Y(_04550_));
 sky130_fd_sc_hd__a21o_1 _13055_ (.A1(_04547_),
    .A2(_04548_),
    .B1(_04549_),
    .X(_04551_));
 sky130_fd_sc_hd__nand3_2 _13056_ (.A(_04543_),
    .B(_04550_),
    .C(_04551_),
    .Y(_04552_));
 sky130_fd_sc_hd__a21o_1 _13057_ (.A1(_04550_),
    .A2(_04551_),
    .B1(_04543_),
    .X(_04553_));
 sky130_fd_sc_hd__a21bo_1 _13058_ (.A1(_04406_),
    .A2(_04414_),
    .B1_N(_04413_),
    .X(_04554_));
 sky130_fd_sc_hd__nand3_4 _13059_ (.A(_04552_),
    .B(_04553_),
    .C(_04554_),
    .Y(_04555_));
 sky130_fd_sc_hd__a21o_1 _13060_ (.A1(_04552_),
    .A2(_04553_),
    .B1(_04554_),
    .X(_04556_));
 sky130_fd_sc_hd__and3_1 _13061_ (.A(_04538_),
    .B(_04555_),
    .C(_04556_),
    .X(_04557_));
 sky130_fd_sc_hd__nand3_2 _13062_ (.A(_04538_),
    .B(_04555_),
    .C(_04556_),
    .Y(_04558_));
 sky130_fd_sc_hd__a21oi_2 _13063_ (.A1(_04555_),
    .A2(_04556_),
    .B1(_04538_),
    .Y(_04559_));
 sky130_fd_sc_hd__a211oi_4 _13064_ (.A1(_04418_),
    .A2(_04421_),
    .B1(_04557_),
    .C1(_04559_),
    .Y(_04560_));
 sky130_fd_sc_hd__o211a_1 _13065_ (.A1(_04557_),
    .A2(_04559_),
    .B1(_04418_),
    .C1(_04421_),
    .X(_04561_));
 sky130_fd_sc_hd__nor3_2 _13066_ (.A(_04527_),
    .B(_04560_),
    .C(_04561_),
    .Y(_04562_));
 sky130_fd_sc_hd__or3_1 _13067_ (.A(_04527_),
    .B(_04560_),
    .C(_04561_),
    .X(_04563_));
 sky130_fd_sc_hd__o21ai_1 _13068_ (.A1(_04560_),
    .A2(_04561_),
    .B1(_04527_),
    .Y(_04564_));
 sky130_fd_sc_hd__o211a_2 _13069_ (.A1(_04423_),
    .A2(_04425_),
    .B1(_04563_),
    .C1(_04564_),
    .X(_04565_));
 sky130_fd_sc_hd__a211oi_2 _13070_ (.A1(_04563_),
    .A2(_04564_),
    .B1(_04423_),
    .C1(_04425_),
    .Y(_04566_));
 sky130_fd_sc_hd__nor3_1 _13071_ (.A(_04505_),
    .B(_04565_),
    .C(_04566_),
    .Y(_04567_));
 sky130_fd_sc_hd__or3_1 _13072_ (.A(_04505_),
    .B(_04565_),
    .C(_04566_),
    .X(_04568_));
 sky130_fd_sc_hd__o21ai_2 _13073_ (.A1(_04565_),
    .A2(_04566_),
    .B1(_04505_),
    .Y(_04569_));
 sky130_fd_sc_hd__o211a_1 _13074_ (.A1(_04428_),
    .A2(_04431_),
    .B1(_04568_),
    .C1(_04569_),
    .X(_04570_));
 sky130_fd_sc_hd__o211ai_1 _13075_ (.A1(_04428_),
    .A2(_04431_),
    .B1(_04568_),
    .C1(_04569_),
    .Y(_04571_));
 sky130_fd_sc_hd__a211o_1 _13076_ (.A1(_04568_),
    .A2(_04569_),
    .B1(_04428_),
    .C1(_04431_),
    .X(_04572_));
 sky130_fd_sc_hd__and3_2 _13077_ (.A(_04468_),
    .B(_04571_),
    .C(_04572_),
    .X(_04573_));
 sky130_fd_sc_hd__a21oi_1 _13078_ (.A1(_04571_),
    .A2(_04572_),
    .B1(_04468_),
    .Y(_04574_));
 sky130_fd_sc_hd__a211oi_2 _13079_ (.A1(_04433_),
    .A2(_04435_),
    .B1(_04573_),
    .C1(_04574_),
    .Y(_04575_));
 sky130_fd_sc_hd__inv_2 _13080_ (.A(_04575_),
    .Y(_04576_));
 sky130_fd_sc_hd__o211a_1 _13081_ (.A1(_04573_),
    .A2(_04574_),
    .B1(_04433_),
    .C1(_04435_),
    .X(_04577_));
 sky130_fd_sc_hd__nor3_1 _13082_ (.A(_04333_),
    .B(_04575_),
    .C(_04577_),
    .Y(_04578_));
 sky130_fd_sc_hd__or3_1 _13083_ (.A(_04333_),
    .B(_04575_),
    .C(_04577_),
    .X(_04579_));
 sky130_fd_sc_hd__o21a_1 _13084_ (.A1(_04575_),
    .A2(_04577_),
    .B1(_04333_),
    .X(_04580_));
 sky130_fd_sc_hd__nor2_2 _13085_ (.A(_04578_),
    .B(_04580_),
    .Y(_04581_));
 sky130_fd_sc_hd__a211o_2 _13086_ (.A1(_04437_),
    .A2(_04439_),
    .B1(_04578_),
    .C1(_04580_),
    .X(_04582_));
 sky130_fd_sc_hd__o211a_1 _13087_ (.A1(_04578_),
    .A2(_04580_),
    .B1(_04437_),
    .C1(_04439_),
    .X(_04583_));
 sky130_fd_sc_hd__xor2_4 _13088_ (.A(_04457_),
    .B(_04581_),
    .X(_04584_));
 sky130_fd_sc_hd__and2b_1 _13089_ (.A_N(_04442_),
    .B(_04584_),
    .X(_04585_));
 sky130_fd_sc_hd__xnor2_4 _13090_ (.A(_04442_),
    .B(_04584_),
    .Y(_04586_));
 sky130_fd_sc_hd__xor2_1 _13091_ (.A(_04442_),
    .B(_04584_),
    .X(_04587_));
 sky130_fd_sc_hd__xnor2_4 _13092_ (.A(_04456_),
    .B(_04586_),
    .Y(_04588_));
 sky130_fd_sc_hd__nor2_1 _13093_ (.A(net9),
    .B(_04588_),
    .Y(_04589_));
 sky130_fd_sc_hd__a221o_1 _13094_ (.A1(net600),
    .A2(\temp[7] ),
    .B1(_02747_),
    .B2(net6),
    .C1(_04589_),
    .X(_04590_));
 sky130_fd_sc_hd__mux2_1 _13095_ (.A0(net753),
    .A1(_04590_),
    .S(net2),
    .X(_00274_));
 sky130_fd_sc_hd__a21oi_2 _13096_ (.A1(_04456_),
    .A2(_04586_),
    .B1(_04585_),
    .Y(_04591_));
 sky130_fd_sc_hd__and2_1 _13097_ (.A(_04501_),
    .B(_04503_),
    .X(_04592_));
 sky130_fd_sc_hd__a22oi_1 _13098_ (.A1(net579),
    .A2(net344),
    .B1(net340),
    .B2(net583),
    .Y(_04593_));
 sky130_fd_sc_hd__and4_2 _13099_ (.A(net579),
    .B(net583),
    .C(net344),
    .D(net340),
    .X(_04594_));
 sky130_fd_sc_hd__nor2_1 _13100_ (.A(_04593_),
    .B(_04594_),
    .Y(_04595_));
 sky130_fd_sc_hd__o21ai_2 _13101_ (.A1(_04469_),
    .A2(_04472_),
    .B1(_04595_),
    .Y(_04596_));
 sky130_fd_sc_hd__or3_1 _13102_ (.A(_04469_),
    .B(_04472_),
    .C(_04595_),
    .X(_04597_));
 sky130_fd_sc_hd__nand2_1 _13103_ (.A(_04596_),
    .B(_04597_),
    .Y(_04598_));
 sky130_fd_sc_hd__nand3_2 _13104_ (.A(_04481_),
    .B(_04483_),
    .C(_04598_),
    .Y(_04599_));
 sky130_fd_sc_hd__inv_2 _13105_ (.A(_04599_),
    .Y(_04600_));
 sky130_fd_sc_hd__a21oi_1 _13106_ (.A1(_04481_),
    .A2(_04483_),
    .B1(_04598_),
    .Y(_04601_));
 sky130_fd_sc_hd__or2_1 _13107_ (.A(_04600_),
    .B(_04601_),
    .X(_04602_));
 sky130_fd_sc_hd__nor2_1 _13108_ (.A(_04458_),
    .B(_04461_),
    .Y(_04603_));
 sky130_fd_sc_hd__xnor2_2 _13109_ (.A(_04602_),
    .B(_04603_),
    .Y(_04604_));
 sky130_fd_sc_hd__nor2_1 _13110_ (.A(_04592_),
    .B(_04604_),
    .Y(_04605_));
 sky130_fd_sc_hd__xor2_2 _13111_ (.A(_04592_),
    .B(_04604_),
    .X(_04606_));
 sky130_fd_sc_hd__xnor2_2 _13112_ (.A(_04464_),
    .B(_04606_),
    .Y(_04607_));
 sky130_fd_sc_hd__and4_1 _13113_ (.A(net562),
    .B(net569),
    .C(net356),
    .D(net355),
    .X(_04608_));
 sky130_fd_sc_hd__a22o_1 _13114_ (.A1(net562),
    .A2(net356),
    .B1(net355),
    .B2(net569),
    .X(_04609_));
 sky130_fd_sc_hd__nand2b_1 _13115_ (.A_N(_04608_),
    .B(_04609_),
    .Y(_04610_));
 sky130_fd_sc_hd__nand2_1 _13116_ (.A(net574),
    .B(net348),
    .Y(_04611_));
 sky130_fd_sc_hd__xnor2_2 _13117_ (.A(_04610_),
    .B(_04611_),
    .Y(_04612_));
 sky130_fd_sc_hd__and2_1 _13118_ (.A(net559),
    .B(net364),
    .X(_04613_));
 sky130_fd_sc_hd__nand4_2 _13119_ (.A(net551),
    .B(net555),
    .C(\mul0.b[18] ),
    .D(\mul0.b[19] ),
    .Y(_04614_));
 sky130_fd_sc_hd__a22o_1 _13120_ (.A1(net551),
    .A2(\mul0.b[18] ),
    .B1(net365),
    .B2(net555),
    .X(_04615_));
 sky130_fd_sc_hd__nand3_1 _13121_ (.A(_04613_),
    .B(_04614_),
    .C(_04615_),
    .Y(_04616_));
 sky130_fd_sc_hd__a21o_1 _13122_ (.A1(_04614_),
    .A2(_04615_),
    .B1(_04613_),
    .X(_04617_));
 sky130_fd_sc_hd__a31o_1 _13123_ (.A1(net562),
    .A2(net364),
    .A3(_04477_),
    .B1(_04476_),
    .X(_04618_));
 sky130_fd_sc_hd__and3_1 _13124_ (.A(_04616_),
    .B(_04617_),
    .C(_04618_),
    .X(_04619_));
 sky130_fd_sc_hd__a21oi_1 _13125_ (.A1(_04616_),
    .A2(_04617_),
    .B1(_04618_),
    .Y(_04620_));
 sky130_fd_sc_hd__nor2_1 _13126_ (.A(_04619_),
    .B(_04620_),
    .Y(_04621_));
 sky130_fd_sc_hd__xnor2_2 _13127_ (.A(_04612_),
    .B(_04621_),
    .Y(_04622_));
 sky130_fd_sc_hd__nand2_1 _13128_ (.A(_04487_),
    .B(_04489_),
    .Y(_04623_));
 sky130_fd_sc_hd__a32o_1 _13129_ (.A1(net537),
    .A2(net389),
    .A3(_04510_),
    .B1(_04509_),
    .B2(net395),
    .X(_04624_));
 sky130_fd_sc_hd__nand4_2 _13130_ (.A(net537),
    .B(net542),
    .C(net382),
    .D(net376),
    .Y(_04625_));
 sky130_fd_sc_hd__a22o_1 _13131_ (.A1(net537),
    .A2(net382),
    .B1(net376),
    .B2(net542),
    .X(_04626_));
 sky130_fd_sc_hd__nand4_2 _13132_ (.A(net546),
    .B(net370),
    .C(_04625_),
    .D(_04626_),
    .Y(_04627_));
 sky130_fd_sc_hd__a22o_1 _13133_ (.A1(net546),
    .A2(net370),
    .B1(_04625_),
    .B2(_04626_),
    .X(_04628_));
 sky130_fd_sc_hd__nand3_1 _13134_ (.A(_04624_),
    .B(_04627_),
    .C(_04628_),
    .Y(_04629_));
 sky130_fd_sc_hd__a21o_1 _13135_ (.A1(_04627_),
    .A2(_04628_),
    .B1(_04624_),
    .X(_04630_));
 sky130_fd_sc_hd__nand3_1 _13136_ (.A(_04623_),
    .B(_04629_),
    .C(_04630_),
    .Y(_04631_));
 sky130_fd_sc_hd__a21o_1 _13137_ (.A1(_04629_),
    .A2(_04630_),
    .B1(_04623_),
    .X(_04632_));
 sky130_fd_sc_hd__a21bo_1 _13138_ (.A1(_04485_),
    .A2(_04492_),
    .B1_N(_04491_),
    .X(_04633_));
 sky130_fd_sc_hd__and3_1 _13139_ (.A(_04631_),
    .B(_04632_),
    .C(_04633_),
    .X(_04634_));
 sky130_fd_sc_hd__nand3_1 _13140_ (.A(_04631_),
    .B(_04632_),
    .C(_04633_),
    .Y(_04635_));
 sky130_fd_sc_hd__a21o_1 _13141_ (.A1(_04631_),
    .A2(_04632_),
    .B1(_04633_),
    .X(_04636_));
 sky130_fd_sc_hd__and3_2 _13142_ (.A(_04622_),
    .B(_04635_),
    .C(_04636_),
    .X(_04637_));
 sky130_fd_sc_hd__a21oi_2 _13143_ (.A1(_04635_),
    .A2(_04636_),
    .B1(_04622_),
    .Y(_04638_));
 sky130_fd_sc_hd__a211oi_4 _13144_ (.A1(_04523_),
    .A2(_04525_),
    .B1(_04637_),
    .C1(_04638_),
    .Y(_04639_));
 sky130_fd_sc_hd__o211a_1 _13145_ (.A1(_04637_),
    .A2(_04638_),
    .B1(_04523_),
    .C1(_04525_),
    .X(_04640_));
 sky130_fd_sc_hd__a211oi_4 _13146_ (.A1(_04496_),
    .A2(_04499_),
    .B1(_04639_),
    .C1(_04640_),
    .Y(_04641_));
 sky130_fd_sc_hd__o211a_1 _13147_ (.A1(_04639_),
    .A2(_04640_),
    .B1(_04496_),
    .C1(_04499_),
    .X(_04642_));
 sky130_fd_sc_hd__nand2_1 _13148_ (.A(_04519_),
    .B(_04521_),
    .Y(_04643_));
 sky130_fd_sc_hd__a21bo_1 _13149_ (.A1(_04528_),
    .A2(_04535_),
    .B1_N(_04534_),
    .X(_04644_));
 sky130_fd_sc_hd__and2_1 _13150_ (.A(net532),
    .B(net387),
    .X(_04645_));
 sky130_fd_sc_hd__a22o_1 _13151_ (.A1(net521),
    .A2(net395),
    .B1(net390),
    .B2(net527),
    .X(_04646_));
 sky130_fd_sc_hd__nand4_1 _13152_ (.A(net521),
    .B(net527),
    .C(net395),
    .D(net391),
    .Y(_04647_));
 sky130_fd_sc_hd__nand2_1 _13153_ (.A(_04646_),
    .B(_04647_),
    .Y(_04648_));
 sky130_fd_sc_hd__xnor2_1 _13154_ (.A(_04645_),
    .B(_04648_),
    .Y(_04649_));
 sky130_fd_sc_hd__nand4_2 _13155_ (.A(net507),
    .B(net511),
    .C(net409),
    .D(net405),
    .Y(_04650_));
 sky130_fd_sc_hd__a22o_1 _13156_ (.A1(net507),
    .A2(net409),
    .B1(net405),
    .B2(net511),
    .X(_04651_));
 sky130_fd_sc_hd__nand4_2 _13157_ (.A(net515),
    .B(net401),
    .C(_04650_),
    .D(_04651_),
    .Y(_04652_));
 sky130_fd_sc_hd__a22o_1 _13158_ (.A1(net515),
    .A2(net401),
    .B1(_04650_),
    .B2(_04651_),
    .X(_04653_));
 sky130_fd_sc_hd__a21bo_1 _13159_ (.A1(_04513_),
    .A2(_04515_),
    .B1_N(_04514_),
    .X(_04654_));
 sky130_fd_sc_hd__nand3_1 _13160_ (.A(_04652_),
    .B(_04653_),
    .C(_04654_),
    .Y(_04655_));
 sky130_fd_sc_hd__a21o_1 _13161_ (.A1(_04652_),
    .A2(_04653_),
    .B1(_04654_),
    .X(_04656_));
 sky130_fd_sc_hd__nand3_1 _13162_ (.A(_04649_),
    .B(_04655_),
    .C(_04656_),
    .Y(_04657_));
 sky130_fd_sc_hd__a21o_1 _13163_ (.A1(_04655_),
    .A2(_04656_),
    .B1(_04649_),
    .X(_04658_));
 sky130_fd_sc_hd__nand3_2 _13164_ (.A(_04644_),
    .B(_04657_),
    .C(_04658_),
    .Y(_04659_));
 sky130_fd_sc_hd__a21o_1 _13165_ (.A1(_04657_),
    .A2(_04658_),
    .B1(_04644_),
    .X(_04660_));
 sky130_fd_sc_hd__nand3_2 _13166_ (.A(_04643_),
    .B(_04659_),
    .C(_04660_),
    .Y(_04661_));
 sky130_fd_sc_hd__a21o_1 _13167_ (.A1(_04659_),
    .A2(_04660_),
    .B1(_04643_),
    .X(_04662_));
 sky130_fd_sc_hd__nand2_1 _13168_ (.A(_04661_),
    .B(_04662_),
    .Y(_04663_));
 sky130_fd_sc_hd__nand2_1 _13169_ (.A(_04530_),
    .B(_04532_),
    .Y(_04664_));
 sky130_fd_sc_hd__o21ba_1 _13170_ (.A1(_04539_),
    .A2(_04541_),
    .B1_N(_04540_),
    .X(_04665_));
 sky130_fd_sc_hd__a22oi_1 _13171_ (.A1(net420),
    .A2(net498),
    .B1(net494),
    .B2(net424),
    .Y(_04666_));
 sky130_fd_sc_hd__and4_1 _13172_ (.A(net424),
    .B(net420),
    .C(net499),
    .D(net494),
    .X(_04667_));
 sky130_fd_sc_hd__and4bb_1 _13173_ (.A_N(_04666_),
    .B_N(_04667_),
    .C(net503),
    .D(net416),
    .X(_04668_));
 sky130_fd_sc_hd__o2bb2a_1 _13174_ (.A1_N(net503),
    .A2_N(net416),
    .B1(_04666_),
    .B2(_04667_),
    .X(_04669_));
 sky130_fd_sc_hd__nor2_1 _13175_ (.A(_04668_),
    .B(_04669_),
    .Y(_04670_));
 sky130_fd_sc_hd__or3_1 _13176_ (.A(_04665_),
    .B(_04668_),
    .C(_04669_),
    .X(_04671_));
 sky130_fd_sc_hd__xnor2_2 _13177_ (.A(_04665_),
    .B(_04670_),
    .Y(_04672_));
 sky130_fd_sc_hd__nand2_1 _13178_ (.A(_04664_),
    .B(_04672_),
    .Y(_04673_));
 sky130_fd_sc_hd__xor2_2 _13179_ (.A(_04664_),
    .B(_04672_),
    .X(_04674_));
 sky130_fd_sc_hd__nand2_1 _13180_ (.A(net429),
    .B(net490),
    .Y(_04675_));
 sky130_fd_sc_hd__and4_1 _13181_ (.A(net439),
    .B(net434),
    .C(net486),
    .D(net482),
    .X(_04676_));
 sky130_fd_sc_hd__a22oi_2 _13182_ (.A1(net434),
    .A2(net486),
    .B1(net482),
    .B2(net439),
    .Y(_04677_));
 sky130_fd_sc_hd__nor2_1 _13183_ (.A(_04676_),
    .B(_04677_),
    .Y(_04678_));
 sky130_fd_sc_hd__xnor2_2 _13184_ (.A(_04675_),
    .B(_04678_),
    .Y(_04679_));
 sky130_fd_sc_hd__and2_1 _13185_ (.A(net442),
    .B(net478),
    .X(_04680_));
 sky130_fd_sc_hd__nand4_1 _13186_ (.A(net451),
    .B(net447),
    .C(net474),
    .D(net470),
    .Y(_04681_));
 sky130_fd_sc_hd__a22o_1 _13187_ (.A1(net447),
    .A2(net474),
    .B1(net470),
    .B2(net451),
    .X(_04682_));
 sky130_fd_sc_hd__nand3_1 _13188_ (.A(_04680_),
    .B(_04681_),
    .C(_04682_),
    .Y(_04683_));
 sky130_fd_sc_hd__a21o_1 _13189_ (.A1(_04681_),
    .A2(_04682_),
    .B1(_04680_),
    .X(_04684_));
 sky130_fd_sc_hd__a21bo_1 _13190_ (.A1(_04544_),
    .A2(_04546_),
    .B1_N(_04545_),
    .X(_04685_));
 sky130_fd_sc_hd__nand3_1 _13191_ (.A(_04683_),
    .B(_04684_),
    .C(_04685_),
    .Y(_04686_));
 sky130_fd_sc_hd__a21o_1 _13192_ (.A1(_04683_),
    .A2(_04684_),
    .B1(_04685_),
    .X(_04687_));
 sky130_fd_sc_hd__nand3_2 _13193_ (.A(_04679_),
    .B(_04686_),
    .C(_04687_),
    .Y(_04688_));
 sky130_fd_sc_hd__a21o_1 _13194_ (.A1(_04686_),
    .A2(_04687_),
    .B1(_04679_),
    .X(_04689_));
 sky130_fd_sc_hd__a21bo_1 _13195_ (.A1(_04543_),
    .A2(_04551_),
    .B1_N(_04550_),
    .X(_04690_));
 sky130_fd_sc_hd__nand3_4 _13196_ (.A(_04688_),
    .B(_04689_),
    .C(_04690_),
    .Y(_04691_));
 sky130_fd_sc_hd__a21o_1 _13197_ (.A1(_04688_),
    .A2(_04689_),
    .B1(_04690_),
    .X(_04692_));
 sky130_fd_sc_hd__and3_1 _13198_ (.A(_04674_),
    .B(_04691_),
    .C(_04692_),
    .X(_04693_));
 sky130_fd_sc_hd__nand3_2 _13199_ (.A(_04674_),
    .B(_04691_),
    .C(_04692_),
    .Y(_04694_));
 sky130_fd_sc_hd__a21oi_2 _13200_ (.A1(_04691_),
    .A2(_04692_),
    .B1(_04674_),
    .Y(_04695_));
 sky130_fd_sc_hd__a211oi_4 _13201_ (.A1(_04555_),
    .A2(_04558_),
    .B1(_04693_),
    .C1(_04695_),
    .Y(_04696_));
 sky130_fd_sc_hd__o211a_1 _13202_ (.A1(_04693_),
    .A2(_04695_),
    .B1(_04555_),
    .C1(_04558_),
    .X(_04697_));
 sky130_fd_sc_hd__nor3_2 _13203_ (.A(_04663_),
    .B(_04696_),
    .C(_04697_),
    .Y(_04698_));
 sky130_fd_sc_hd__or3_2 _13204_ (.A(_04663_),
    .B(_04696_),
    .C(_04697_),
    .X(_04699_));
 sky130_fd_sc_hd__o21ai_2 _13205_ (.A1(_04696_),
    .A2(_04697_),
    .B1(_04663_),
    .Y(_04700_));
 sky130_fd_sc_hd__o211a_4 _13206_ (.A1(_04560_),
    .A2(_04562_),
    .B1(_04699_),
    .C1(_04700_),
    .X(_04701_));
 sky130_fd_sc_hd__a211oi_4 _13207_ (.A1(_04699_),
    .A2(_04700_),
    .B1(_04560_),
    .C1(_04562_),
    .Y(_04702_));
 sky130_fd_sc_hd__nor4_2 _13208_ (.A(_04641_),
    .B(_04642_),
    .C(_04701_),
    .D(_04702_),
    .Y(_04703_));
 sky130_fd_sc_hd__or4_2 _13209_ (.A(_04641_),
    .B(_04642_),
    .C(_04701_),
    .D(_04702_),
    .X(_04704_));
 sky130_fd_sc_hd__o22ai_4 _13210_ (.A1(_04641_),
    .A2(_04642_),
    .B1(_04701_),
    .B2(_04702_),
    .Y(_04705_));
 sky130_fd_sc_hd__o211ai_4 _13211_ (.A1(_04565_),
    .A2(_04567_),
    .B1(_04704_),
    .C1(_04705_),
    .Y(_04706_));
 sky130_fd_sc_hd__a211o_1 _13212_ (.A1(_04704_),
    .A2(_04705_),
    .B1(_04565_),
    .C1(_04567_),
    .X(_04707_));
 sky130_fd_sc_hd__nand3_4 _13213_ (.A(_04607_),
    .B(_04706_),
    .C(_04707_),
    .Y(_04708_));
 sky130_fd_sc_hd__a21o_1 _13214_ (.A1(_04706_),
    .A2(_04707_),
    .B1(_04607_),
    .X(_04709_));
 sky130_fd_sc_hd__o211ai_4 _13215_ (.A1(_04570_),
    .A2(_04573_),
    .B1(_04708_),
    .C1(_04709_),
    .Y(_04710_));
 sky130_fd_sc_hd__a211o_1 _13216_ (.A1(_04708_),
    .A2(_04709_),
    .B1(_04570_),
    .C1(_04573_),
    .X(_04711_));
 sky130_fd_sc_hd__and3_1 _13217_ (.A(_04466_),
    .B(_04710_),
    .C(_04711_),
    .X(_04712_));
 sky130_fd_sc_hd__nand3_2 _13218_ (.A(_04466_),
    .B(_04710_),
    .C(_04711_),
    .Y(_04713_));
 sky130_fd_sc_hd__a21oi_1 _13219_ (.A1(_04710_),
    .A2(_04711_),
    .B1(_04466_),
    .Y(_04714_));
 sky130_fd_sc_hd__a211o_2 _13220_ (.A1(_04576_),
    .A2(_04579_),
    .B1(_04712_),
    .C1(_04714_),
    .X(_04715_));
 sky130_fd_sc_hd__o211ai_1 _13221_ (.A1(_04712_),
    .A2(_04714_),
    .B1(_04576_),
    .C1(_04579_),
    .Y(_04716_));
 sky130_fd_sc_hd__nand2_2 _13222_ (.A(_04715_),
    .B(_04716_),
    .Y(_04717_));
 sky130_fd_sc_hd__xnor2_4 _13223_ (.A(_04582_),
    .B(_04717_),
    .Y(_04718_));
 sky130_fd_sc_hd__xnor2_4 _13224_ (.A(_04591_),
    .B(_04718_),
    .Y(_04719_));
 sky130_fd_sc_hd__nor2_1 _13225_ (.A(net9),
    .B(_04719_),
    .Y(_04720_));
 sky130_fd_sc_hd__a221o_1 _13226_ (.A1(net599),
    .A2(net709),
    .B1(_02748_),
    .B2(net6),
    .C1(_04720_),
    .X(_04721_));
 sky130_fd_sc_hd__mux2_1 _13227_ (.A0(net865),
    .A1(_04721_),
    .S(net3),
    .X(_00275_));
 sky130_fd_sc_hd__a31o_1 _13228_ (.A1(_04330_),
    .A2(_04463_),
    .A3(_04606_),
    .B1(_04605_),
    .X(_04722_));
 sky130_fd_sc_hd__inv_2 _13229_ (.A(_04722_),
    .Y(_04723_));
 sky130_fd_sc_hd__or2_1 _13230_ (.A(_04639_),
    .B(_04641_),
    .X(_04724_));
 sky130_fd_sc_hd__o21ba_1 _13231_ (.A1(_04612_),
    .A2(_04620_),
    .B1_N(_04619_),
    .X(_04725_));
 sky130_fd_sc_hd__a31oi_2 _13232_ (.A1(net573),
    .A2(net348),
    .A3(_04609_),
    .B1(_04608_),
    .Y(_04726_));
 sky130_fd_sc_hd__and4_1 _13233_ (.A(net573),
    .B(net579),
    .C(net344),
    .D(net340),
    .X(_04727_));
 sky130_fd_sc_hd__a22oi_1 _13234_ (.A1(net573),
    .A2(net344),
    .B1(net340),
    .B2(net579),
    .Y(_04728_));
 sky130_fd_sc_hd__and4bb_1 _13235_ (.A_N(_04727_),
    .B_N(_04728_),
    .C(net583),
    .D(net337),
    .X(_04729_));
 sky130_fd_sc_hd__o2bb2a_1 _13236_ (.A1_N(net583),
    .A2_N(net337),
    .B1(_04727_),
    .B2(_04728_),
    .X(_04730_));
 sky130_fd_sc_hd__nor3_1 _13237_ (.A(_04726_),
    .B(_04729_),
    .C(_04730_),
    .Y(_04731_));
 sky130_fd_sc_hd__o21ai_1 _13238_ (.A1(_04729_),
    .A2(_04730_),
    .B1(_04726_),
    .Y(_04732_));
 sky130_fd_sc_hd__and2b_1 _13239_ (.A_N(_04731_),
    .B(_04732_),
    .X(_04733_));
 sky130_fd_sc_hd__xnor2_2 _13240_ (.A(_04594_),
    .B(_04733_),
    .Y(_04734_));
 sky130_fd_sc_hd__or2_1 _13241_ (.A(_04725_),
    .B(_04734_),
    .X(_04735_));
 sky130_fd_sc_hd__xnor2_2 _13242_ (.A(_04725_),
    .B(_04734_),
    .Y(_04736_));
 sky130_fd_sc_hd__xor2_1 _13243_ (.A(_04596_),
    .B(_04736_),
    .X(_04737_));
 sky130_fd_sc_hd__or2_1 _13244_ (.A(_04458_),
    .B(_04601_),
    .X(_04738_));
 sky130_fd_sc_hd__and3_1 _13245_ (.A(_04599_),
    .B(_04737_),
    .C(_04738_),
    .X(_04739_));
 sky130_fd_sc_hd__a21oi_1 _13246_ (.A1(_04599_),
    .A2(_04738_),
    .B1(_04737_),
    .Y(_04740_));
 sky130_fd_sc_hd__nor2_1 _13247_ (.A(_04739_),
    .B(_04740_),
    .Y(_04741_));
 sky130_fd_sc_hd__nand2_1 _13248_ (.A(_04724_),
    .B(_04741_),
    .Y(_04742_));
 sky130_fd_sc_hd__xor2_1 _13249_ (.A(_04724_),
    .B(_04741_),
    .X(_04743_));
 sky130_fd_sc_hd__and3b_1 _13250_ (.A_N(_04601_),
    .B(_04461_),
    .C(_04599_),
    .X(_04744_));
 sky130_fd_sc_hd__nand2_1 _13251_ (.A(_04743_),
    .B(_04744_),
    .Y(_04745_));
 sky130_fd_sc_hd__xor2_1 _13252_ (.A(_04743_),
    .B(_04744_),
    .X(_04746_));
 sky130_fd_sc_hd__a22o_1 _13253_ (.A1(net559),
    .A2(net356),
    .B1(net355),
    .B2(net563),
    .X(_04747_));
 sky130_fd_sc_hd__and3_1 _13254_ (.A(net559),
    .B(net563),
    .C(net355),
    .X(_04748_));
 sky130_fd_sc_hd__a21bo_1 _13255_ (.A1(net356),
    .A2(_04748_),
    .B1_N(_04747_),
    .X(_04749_));
 sky130_fd_sc_hd__nand2_1 _13256_ (.A(net569),
    .B(net348),
    .Y(_04750_));
 sky130_fd_sc_hd__xnor2_1 _13257_ (.A(_04749_),
    .B(_04750_),
    .Y(_04751_));
 sky130_fd_sc_hd__nand4_2 _13258_ (.A(net546),
    .B(net550),
    .C(net631),
    .D(net365),
    .Y(_04752_));
 sky130_fd_sc_hd__a22o_1 _13259_ (.A1(net546),
    .A2(net631),
    .B1(net365),
    .B2(net550),
    .X(_04753_));
 sky130_fd_sc_hd__nand4_2 _13260_ (.A(net554),
    .B(net364),
    .C(_04752_),
    .D(_04753_),
    .Y(_04754_));
 sky130_fd_sc_hd__a22o_1 _13261_ (.A1(net554),
    .A2(net364),
    .B1(_04752_),
    .B2(_04753_),
    .X(_04755_));
 sky130_fd_sc_hd__a21bo_1 _13262_ (.A1(_04613_),
    .A2(_04615_),
    .B1_N(_04614_),
    .X(_04756_));
 sky130_fd_sc_hd__and3_1 _13263_ (.A(_04754_),
    .B(_04755_),
    .C(_04756_),
    .X(_04757_));
 sky130_fd_sc_hd__a21oi_1 _13264_ (.A1(_04754_),
    .A2(_04755_),
    .B1(_04756_),
    .Y(_04758_));
 sky130_fd_sc_hd__nor2_1 _13265_ (.A(_04757_),
    .B(_04758_),
    .Y(_04759_));
 sky130_fd_sc_hd__xnor2_1 _13266_ (.A(_04751_),
    .B(_04759_),
    .Y(_04760_));
 sky130_fd_sc_hd__nand2_1 _13267_ (.A(_04625_),
    .B(_04627_),
    .Y(_04761_));
 sky130_fd_sc_hd__a21boi_1 _13268_ (.A1(_04645_),
    .A2(_04646_),
    .B1_N(_04647_),
    .Y(_04762_));
 sky130_fd_sc_hd__and4_1 _13269_ (.A(net532),
    .B(net537),
    .C(net382),
    .D(net376),
    .X(_04763_));
 sky130_fd_sc_hd__a22oi_1 _13270_ (.A1(net532),
    .A2(net382),
    .B1(net376),
    .B2(net537),
    .Y(_04764_));
 sky130_fd_sc_hd__and4bb_1 _13271_ (.A_N(_04763_),
    .B_N(_04764_),
    .C(net542),
    .D(net370),
    .X(_04765_));
 sky130_fd_sc_hd__o2bb2a_1 _13272_ (.A1_N(net542),
    .A2_N(net370),
    .B1(_04763_),
    .B2(_04764_),
    .X(_04766_));
 sky130_fd_sc_hd__or3_2 _13273_ (.A(_04762_),
    .B(_04765_),
    .C(_04766_),
    .X(_04767_));
 sky130_fd_sc_hd__o21ai_1 _13274_ (.A1(_04765_),
    .A2(_04766_),
    .B1(_04762_),
    .Y(_04768_));
 sky130_fd_sc_hd__nand3_2 _13275_ (.A(_04761_),
    .B(_04767_),
    .C(_04768_),
    .Y(_04769_));
 sky130_fd_sc_hd__a21o_1 _13276_ (.A1(_04767_),
    .A2(_04768_),
    .B1(_04761_),
    .X(_04770_));
 sky130_fd_sc_hd__a21bo_1 _13277_ (.A1(_04623_),
    .A2(_04630_),
    .B1_N(_04629_),
    .X(_04771_));
 sky130_fd_sc_hd__and3_2 _13278_ (.A(_04769_),
    .B(_04770_),
    .C(_04771_),
    .X(_04772_));
 sky130_fd_sc_hd__a21oi_2 _13279_ (.A1(_04769_),
    .A2(_04770_),
    .B1(_04771_),
    .Y(_04773_));
 sky130_fd_sc_hd__nor3b_4 _13280_ (.A(_04772_),
    .B(_04773_),
    .C_N(_04760_),
    .Y(_04774_));
 sky130_fd_sc_hd__o21ba_1 _13281_ (.A1(_04772_),
    .A2(_04773_),
    .B1_N(_04760_),
    .X(_04775_));
 sky130_fd_sc_hd__a211o_1 _13282_ (.A1(_04659_),
    .A2(_04661_),
    .B1(_04774_),
    .C1(_04775_),
    .X(_04776_));
 sky130_fd_sc_hd__o211ai_2 _13283_ (.A1(_04774_),
    .A2(_04775_),
    .B1(_04659_),
    .C1(_04661_),
    .Y(_04777_));
 sky130_fd_sc_hd__o211ai_2 _13284_ (.A1(_04634_),
    .A2(_04637_),
    .B1(_04776_),
    .C1(_04777_),
    .Y(_04778_));
 sky130_fd_sc_hd__a211o_1 _13285_ (.A1(_04776_),
    .A2(_04777_),
    .B1(_04634_),
    .C1(_04637_),
    .X(_04779_));
 sky130_fd_sc_hd__nand2_1 _13286_ (.A(_04778_),
    .B(_04779_),
    .Y(_04780_));
 sky130_fd_sc_hd__nand2_1 _13287_ (.A(_04655_),
    .B(_04657_),
    .Y(_04781_));
 sky130_fd_sc_hd__a22o_1 _13288_ (.A1(net517),
    .A2(net397),
    .B1(net392),
    .B2(net524),
    .X(_04782_));
 sky130_fd_sc_hd__nand4_2 _13289_ (.A(net517),
    .B(net521),
    .C(net397),
    .D(net392),
    .Y(_04783_));
 sky130_fd_sc_hd__nand4_2 _13290_ (.A(net527),
    .B(net387),
    .C(_04782_),
    .D(_04783_),
    .Y(_04784_));
 sky130_fd_sc_hd__a22o_1 _13291_ (.A1(net527),
    .A2(net387),
    .B1(_04782_),
    .B2(_04783_),
    .X(_04785_));
 sky130_fd_sc_hd__and2_1 _13292_ (.A(_04784_),
    .B(_04785_),
    .X(_04786_));
 sky130_fd_sc_hd__a22oi_1 _13293_ (.A1(net504),
    .A2(net411),
    .B1(net407),
    .B2(net508),
    .Y(_04787_));
 sky130_fd_sc_hd__and4_1 _13294_ (.A(net504),
    .B(net508),
    .C(net411),
    .D(net407),
    .X(_04788_));
 sky130_fd_sc_hd__and4bb_1 _13295_ (.A_N(_04787_),
    .B_N(_04788_),
    .C(net512),
    .D(net403),
    .X(_04789_));
 sky130_fd_sc_hd__o2bb2a_1 _13296_ (.A1_N(net512),
    .A2_N(net403),
    .B1(_04787_),
    .B2(_04788_),
    .X(_04790_));
 sky130_fd_sc_hd__nor2_1 _13297_ (.A(_04789_),
    .B(_04790_),
    .Y(_04791_));
 sky130_fd_sc_hd__and2_1 _13298_ (.A(_04650_),
    .B(_04652_),
    .X(_04792_));
 sky130_fd_sc_hd__and2b_2 _13299_ (.A_N(_04792_),
    .B(_04791_),
    .X(_04793_));
 sky130_fd_sc_hd__xnor2_1 _13300_ (.A(_04791_),
    .B(_04792_),
    .Y(_04794_));
 sky130_fd_sc_hd__and2_2 _13301_ (.A(_04786_),
    .B(_04794_),
    .X(_04795_));
 sky130_fd_sc_hd__xnor2_1 _13302_ (.A(_04786_),
    .B(_04794_),
    .Y(_04796_));
 sky130_fd_sc_hd__a21o_2 _13303_ (.A1(_04671_),
    .A2(_04673_),
    .B1(_04796_),
    .X(_04797_));
 sky130_fd_sc_hd__nand3_2 _13304_ (.A(_04671_),
    .B(_04673_),
    .C(_04796_),
    .Y(_04798_));
 sky130_fd_sc_hd__and3_2 _13305_ (.A(_04781_),
    .B(_04797_),
    .C(_04798_),
    .X(_04799_));
 sky130_fd_sc_hd__nand3_2 _13306_ (.A(_04781_),
    .B(_04797_),
    .C(_04798_),
    .Y(_04800_));
 sky130_fd_sc_hd__a21oi_2 _13307_ (.A1(_04797_),
    .A2(_04798_),
    .B1(_04781_),
    .Y(_04801_));
 sky130_fd_sc_hd__or2_2 _13308_ (.A(_04667_),
    .B(_04668_),
    .X(_04802_));
 sky130_fd_sc_hd__o21ba_1 _13309_ (.A1(_04675_),
    .A2(_04677_),
    .B1_N(_04676_),
    .X(_04803_));
 sky130_fd_sc_hd__a22oi_1 _13310_ (.A1(net420),
    .A2(net494),
    .B1(net490),
    .B2(net424),
    .Y(_04804_));
 sky130_fd_sc_hd__and4_1 _13311_ (.A(net424),
    .B(net420),
    .C(net494),
    .D(net490),
    .X(_04805_));
 sky130_fd_sc_hd__and4bb_1 _13312_ (.A_N(_04804_),
    .B_N(_04805_),
    .C(net416),
    .D(net499),
    .X(_04806_));
 sky130_fd_sc_hd__o2bb2a_1 _13313_ (.A1_N(net416),
    .A2_N(net498),
    .B1(_04804_),
    .B2(_04805_),
    .X(_04807_));
 sky130_fd_sc_hd__nor2_1 _13314_ (.A(_04806_),
    .B(_04807_),
    .Y(_04808_));
 sky130_fd_sc_hd__or3_2 _13315_ (.A(_04803_),
    .B(_04806_),
    .C(_04807_),
    .X(_04809_));
 sky130_fd_sc_hd__xnor2_2 _13316_ (.A(_04803_),
    .B(_04808_),
    .Y(_04810_));
 sky130_fd_sc_hd__nand2_2 _13317_ (.A(_04802_),
    .B(_04810_),
    .Y(_04811_));
 sky130_fd_sc_hd__xor2_2 _13318_ (.A(_04802_),
    .B(_04810_),
    .X(_04812_));
 sky130_fd_sc_hd__nand2_1 _13319_ (.A(net429),
    .B(net486),
    .Y(_04813_));
 sky130_fd_sc_hd__and4_1 _13320_ (.A(net439),
    .B(net434),
    .C(net482),
    .D(net478),
    .X(_04814_));
 sky130_fd_sc_hd__a22o_1 _13321_ (.A1(net434),
    .A2(net482),
    .B1(net478),
    .B2(net439),
    .X(_04815_));
 sky130_fd_sc_hd__and2b_1 _13322_ (.A_N(_04814_),
    .B(_04815_),
    .X(_04816_));
 sky130_fd_sc_hd__xnor2_2 _13323_ (.A(_04813_),
    .B(_04816_),
    .Y(_04817_));
 sky130_fd_sc_hd__and2_1 _13324_ (.A(net442),
    .B(net474),
    .X(_04818_));
 sky130_fd_sc_hd__nand4_1 _13325_ (.A(net451),
    .B(net447),
    .C(net470),
    .D(net466),
    .Y(_04819_));
 sky130_fd_sc_hd__a22o_1 _13326_ (.A1(net447),
    .A2(net470),
    .B1(net466),
    .B2(net451),
    .X(_04820_));
 sky130_fd_sc_hd__nand3_1 _13327_ (.A(_04818_),
    .B(_04819_),
    .C(_04820_),
    .Y(_04821_));
 sky130_fd_sc_hd__a21o_1 _13328_ (.A1(_04819_),
    .A2(_04820_),
    .B1(_04818_),
    .X(_04822_));
 sky130_fd_sc_hd__a21bo_1 _13329_ (.A1(_04680_),
    .A2(_04682_),
    .B1_N(_04681_),
    .X(_04823_));
 sky130_fd_sc_hd__nand3_1 _13330_ (.A(_04821_),
    .B(_04822_),
    .C(_04823_),
    .Y(_04824_));
 sky130_fd_sc_hd__a21o_1 _13331_ (.A1(_04821_),
    .A2(_04822_),
    .B1(_04823_),
    .X(_04825_));
 sky130_fd_sc_hd__nand3_2 _13332_ (.A(_04817_),
    .B(_04824_),
    .C(_04825_),
    .Y(_04826_));
 sky130_fd_sc_hd__a21o_1 _13333_ (.A1(_04824_),
    .A2(_04825_),
    .B1(_04817_),
    .X(_04827_));
 sky130_fd_sc_hd__a21bo_1 _13334_ (.A1(_04679_),
    .A2(_04687_),
    .B1_N(_04686_),
    .X(_04828_));
 sky130_fd_sc_hd__nand3_4 _13335_ (.A(_04826_),
    .B(_04827_),
    .C(_04828_),
    .Y(_04829_));
 sky130_fd_sc_hd__a21o_1 _13336_ (.A1(_04826_),
    .A2(_04827_),
    .B1(_04828_),
    .X(_04830_));
 sky130_fd_sc_hd__and3_1 _13337_ (.A(_04812_),
    .B(_04829_),
    .C(_04830_),
    .X(_04831_));
 sky130_fd_sc_hd__nand3_2 _13338_ (.A(_04812_),
    .B(_04829_),
    .C(_04830_),
    .Y(_04832_));
 sky130_fd_sc_hd__a21oi_2 _13339_ (.A1(_04829_),
    .A2(_04830_),
    .B1(_04812_),
    .Y(_04833_));
 sky130_fd_sc_hd__a211oi_4 _13340_ (.A1(_04691_),
    .A2(_04694_),
    .B1(_04831_),
    .C1(_04833_),
    .Y(_04834_));
 sky130_fd_sc_hd__o211a_1 _13341_ (.A1(_04831_),
    .A2(_04833_),
    .B1(_04691_),
    .C1(_04694_),
    .X(_04835_));
 sky130_fd_sc_hd__nor4_2 _13342_ (.A(_04799_),
    .B(_04801_),
    .C(_04834_),
    .D(_04835_),
    .Y(_04836_));
 sky130_fd_sc_hd__or4_2 _13343_ (.A(_04799_),
    .B(_04801_),
    .C(_04834_),
    .D(_04835_),
    .X(_04837_));
 sky130_fd_sc_hd__o22ai_4 _13344_ (.A1(_04799_),
    .A2(_04801_),
    .B1(_04834_),
    .B2(_04835_),
    .Y(_04838_));
 sky130_fd_sc_hd__o211a_2 _13345_ (.A1(_04696_),
    .A2(_04698_),
    .B1(_04837_),
    .C1(_04838_),
    .X(_04839_));
 sky130_fd_sc_hd__a211oi_4 _13346_ (.A1(_04837_),
    .A2(_04838_),
    .B1(_04696_),
    .C1(_04698_),
    .Y(_04840_));
 sky130_fd_sc_hd__nor3_2 _13347_ (.A(_04780_),
    .B(_04839_),
    .C(_04840_),
    .Y(_04841_));
 sky130_fd_sc_hd__or3_2 _13348_ (.A(_04780_),
    .B(_04839_),
    .C(_04840_),
    .X(_04842_));
 sky130_fd_sc_hd__o21ai_2 _13349_ (.A1(_04839_),
    .A2(_04840_),
    .B1(_04780_),
    .Y(_04843_));
 sky130_fd_sc_hd__o211ai_4 _13350_ (.A1(_04701_),
    .A2(_04703_),
    .B1(_04842_),
    .C1(_04843_),
    .Y(_04844_));
 sky130_fd_sc_hd__a211o_1 _13351_ (.A1(_04842_),
    .A2(_04843_),
    .B1(_04701_),
    .C1(_04703_),
    .X(_04845_));
 sky130_fd_sc_hd__and3_1 _13352_ (.A(_04746_),
    .B(_04844_),
    .C(_04845_),
    .X(_04846_));
 sky130_fd_sc_hd__nand3_1 _13353_ (.A(_04746_),
    .B(_04844_),
    .C(_04845_),
    .Y(_04847_));
 sky130_fd_sc_hd__a21oi_1 _13354_ (.A1(_04844_),
    .A2(_04845_),
    .B1(_04746_),
    .Y(_04848_));
 sky130_fd_sc_hd__a211oi_2 _13355_ (.A1(_04706_),
    .A2(_04708_),
    .B1(_04846_),
    .C1(_04848_),
    .Y(_04849_));
 sky130_fd_sc_hd__o211a_1 _13356_ (.A1(_04846_),
    .A2(_04848_),
    .B1(_04706_),
    .C1(_04708_),
    .X(_04850_));
 sky130_fd_sc_hd__nor3_2 _13357_ (.A(_04723_),
    .B(_04849_),
    .C(_04850_),
    .Y(_04851_));
 sky130_fd_sc_hd__o21a_1 _13358_ (.A1(_04849_),
    .A2(_04850_),
    .B1(_04723_),
    .X(_04852_));
 sky130_fd_sc_hd__a211oi_4 _13359_ (.A1(_04710_),
    .A2(_04713_),
    .B1(_04851_),
    .C1(_04852_),
    .Y(_04853_));
 sky130_fd_sc_hd__o211a_1 _13360_ (.A1(_04851_),
    .A2(_04852_),
    .B1(_04710_),
    .C1(_04713_),
    .X(_04854_));
 sky130_fd_sc_hd__or3_1 _13361_ (.A(_04715_),
    .B(_04853_),
    .C(_04854_),
    .X(_04855_));
 sky130_fd_sc_hd__o21ai_2 _13362_ (.A1(_04853_),
    .A2(_04854_),
    .B1(_04715_),
    .Y(_04856_));
 sky130_fd_sc_hd__nand2_4 _13363_ (.A(_04855_),
    .B(_04856_),
    .Y(_04857_));
 sky130_fd_sc_hd__o21a_1 _13364_ (.A1(_04442_),
    .A2(_04583_),
    .B1(_04582_),
    .X(_04858_));
 sky130_fd_sc_hd__or2_1 _13365_ (.A(_04717_),
    .B(_04858_),
    .X(_04859_));
 sky130_fd_sc_hd__nor2_2 _13366_ (.A(_04587_),
    .B(_04718_),
    .Y(_04860_));
 sky130_fd_sc_hd__a21boi_4 _13367_ (.A1(_04456_),
    .A2(_04860_),
    .B1_N(_04859_),
    .Y(_04861_));
 sky130_fd_sc_hd__xnor2_4 _13368_ (.A(_04857_),
    .B(_04861_),
    .Y(_04862_));
 sky130_fd_sc_hd__nor2_1 _13369_ (.A(net9),
    .B(_04862_),
    .Y(_04863_));
 sky130_fd_sc_hd__a221o_1 _13370_ (.A1(net600),
    .A2(net836),
    .B1(_02749_),
    .B2(net6),
    .C1(_04863_),
    .X(_04864_));
 sky130_fd_sc_hd__mux2_1 _13371_ (.A0(net961),
    .A1(_04864_),
    .S(net1),
    .X(_00276_));
 sky130_fd_sc_hd__o32a_2 _13372_ (.A1(_04715_),
    .A2(_04853_),
    .A3(_04854_),
    .B1(_04857_),
    .B2(_04861_),
    .X(_04865_));
 sky130_fd_sc_hd__nand2_1 _13373_ (.A(_04776_),
    .B(_04778_),
    .Y(_04866_));
 sky130_fd_sc_hd__a21o_1 _13374_ (.A1(_04594_),
    .A2(_04732_),
    .B1(_04731_),
    .X(_04867_));
 sky130_fd_sc_hd__o21ba_1 _13375_ (.A1(_04751_),
    .A2(_04758_),
    .B1_N(_04757_),
    .X(_04868_));
 sky130_fd_sc_hd__or2_1 _13376_ (.A(_04727_),
    .B(_04729_),
    .X(_04869_));
 sky130_fd_sc_hd__a32oi_4 _13377_ (.A1(net568),
    .A2(net348),
    .A3(_04747_),
    .B1(_04748_),
    .B2(net356),
    .Y(_04870_));
 sky130_fd_sc_hd__a22oi_1 _13378_ (.A1(net568),
    .A2(net344),
    .B1(net340),
    .B2(net573),
    .Y(_04871_));
 sky130_fd_sc_hd__and4_1 _13379_ (.A(net568),
    .B(net573),
    .C(net344),
    .D(net340),
    .X(_04872_));
 sky130_fd_sc_hd__o2bb2a_1 _13380_ (.A1_N(net579),
    .A2_N(net337),
    .B1(_04871_),
    .B2(_04872_),
    .X(_04873_));
 sky130_fd_sc_hd__and4bb_1 _13381_ (.A_N(_04871_),
    .B_N(_04872_),
    .C(net579),
    .D(net337),
    .X(_04874_));
 sky130_fd_sc_hd__or2_1 _13382_ (.A(_04873_),
    .B(_04874_),
    .X(_04875_));
 sky130_fd_sc_hd__or2_1 _13383_ (.A(_04870_),
    .B(_04875_),
    .X(_04876_));
 sky130_fd_sc_hd__xor2_1 _13384_ (.A(_04870_),
    .B(_04875_),
    .X(_04877_));
 sky130_fd_sc_hd__nand2_1 _13385_ (.A(_04869_),
    .B(_04877_),
    .Y(_04878_));
 sky130_fd_sc_hd__xnor2_1 _13386_ (.A(_04869_),
    .B(_04877_),
    .Y(_04879_));
 sky130_fd_sc_hd__or2_1 _13387_ (.A(_04868_),
    .B(_04879_),
    .X(_04880_));
 sky130_fd_sc_hd__xor2_1 _13388_ (.A(_04868_),
    .B(_04879_),
    .X(_04881_));
 sky130_fd_sc_hd__nand2_1 _13389_ (.A(_04867_),
    .B(_04881_),
    .Y(_04882_));
 sky130_fd_sc_hd__xor2_1 _13390_ (.A(_04867_),
    .B(_04881_),
    .X(_04883_));
 sky130_fd_sc_hd__o21ai_2 _13391_ (.A1(_04596_),
    .A2(_04736_),
    .B1(_04735_),
    .Y(_04884_));
 sky130_fd_sc_hd__nand2_1 _13392_ (.A(_04883_),
    .B(_04884_),
    .Y(_04885_));
 sky130_fd_sc_hd__xnor2_1 _13393_ (.A(_04883_),
    .B(_04884_),
    .Y(_04886_));
 sky130_fd_sc_hd__nand2_1 _13394_ (.A(net583),
    .B(net336),
    .Y(_04887_));
 sky130_fd_sc_hd__or2_1 _13395_ (.A(_04886_),
    .B(_04887_),
    .X(_04888_));
 sky130_fd_sc_hd__xnor2_1 _13396_ (.A(_04886_),
    .B(_04887_),
    .Y(_04889_));
 sky130_fd_sc_hd__and2b_1 _13397_ (.A_N(_04889_),
    .B(_04866_),
    .X(_04890_));
 sky130_fd_sc_hd__xnor2_1 _13398_ (.A(_04866_),
    .B(_04889_),
    .Y(_04891_));
 sky130_fd_sc_hd__and2_1 _13399_ (.A(_04739_),
    .B(_04891_),
    .X(_04892_));
 sky130_fd_sc_hd__nor2_1 _13400_ (.A(_04739_),
    .B(_04891_),
    .Y(_04893_));
 sky130_fd_sc_hd__a22o_1 _13401_ (.A1(net554),
    .A2(net356),
    .B1(net355),
    .B2(net558),
    .X(_04894_));
 sky130_fd_sc_hd__nand4_2 _13402_ (.A(net554),
    .B(net558),
    .C(net356),
    .D(net355),
    .Y(_04895_));
 sky130_fd_sc_hd__a22o_1 _13403_ (.A1(net563),
    .A2(\mul0.b[23] ),
    .B1(_04894_),
    .B2(_04895_),
    .X(_04896_));
 sky130_fd_sc_hd__nand4_1 _13404_ (.A(net563),
    .B(net348),
    .C(_04894_),
    .D(_04895_),
    .Y(_04897_));
 sky130_fd_sc_hd__nand2_1 _13405_ (.A(_04896_),
    .B(_04897_),
    .Y(_04898_));
 sky130_fd_sc_hd__nand2_1 _13406_ (.A(net550),
    .B(net364),
    .Y(_04899_));
 sky130_fd_sc_hd__a22o_1 _13407_ (.A1(net542),
    .A2(net632),
    .B1(net367),
    .B2(\mul0.a[8] ),
    .X(_04900_));
 sky130_fd_sc_hd__nand4_1 _13408_ (.A(net542),
    .B(net546),
    .C(net632),
    .D(net367),
    .Y(_04901_));
 sky130_fd_sc_hd__nand2_1 _13409_ (.A(_04900_),
    .B(_04901_),
    .Y(_04902_));
 sky130_fd_sc_hd__xor2_2 _13410_ (.A(_04899_),
    .B(_04902_),
    .X(_04903_));
 sky130_fd_sc_hd__and2_1 _13411_ (.A(_04752_),
    .B(_04754_),
    .X(_04904_));
 sky130_fd_sc_hd__nand2b_1 _13412_ (.A_N(_04904_),
    .B(_04903_),
    .Y(_04905_));
 sky130_fd_sc_hd__xnor2_1 _13413_ (.A(_04903_),
    .B(_04904_),
    .Y(_04906_));
 sky130_fd_sc_hd__nand2b_1 _13414_ (.A_N(_04898_),
    .B(_04906_),
    .Y(_04907_));
 sky130_fd_sc_hd__xnor2_1 _13415_ (.A(_04898_),
    .B(_04906_),
    .Y(_04908_));
 sky130_fd_sc_hd__or2_1 _13416_ (.A(_04763_),
    .B(_04765_),
    .X(_04909_));
 sky130_fd_sc_hd__a22oi_1 _13417_ (.A1(net527),
    .A2(net383),
    .B1(net377),
    .B2(net532),
    .Y(_04910_));
 sky130_fd_sc_hd__and4_1 _13418_ (.A(net527),
    .B(net532),
    .C(net383),
    .D(net377),
    .X(_04911_));
 sky130_fd_sc_hd__o2bb2a_1 _13419_ (.A1_N(net537),
    .A2_N(net370),
    .B1(_04910_),
    .B2(_04911_),
    .X(_04912_));
 sky130_fd_sc_hd__and4bb_1 _13420_ (.A_N(_04910_),
    .B_N(_04911_),
    .C(net537),
    .D(net370),
    .X(_04913_));
 sky130_fd_sc_hd__a211o_1 _13421_ (.A1(_04783_),
    .A2(_04784_),
    .B1(_04912_),
    .C1(_04913_),
    .X(_04914_));
 sky130_fd_sc_hd__o211ai_1 _13422_ (.A1(_04912_),
    .A2(_04913_),
    .B1(_04783_),
    .C1(_04784_),
    .Y(_04915_));
 sky130_fd_sc_hd__and2_1 _13423_ (.A(_04914_),
    .B(_04915_),
    .X(_04916_));
 sky130_fd_sc_hd__nand2_1 _13424_ (.A(_04909_),
    .B(_04916_),
    .Y(_04917_));
 sky130_fd_sc_hd__xnor2_2 _13425_ (.A(_04909_),
    .B(_04916_),
    .Y(_04918_));
 sky130_fd_sc_hd__a21oi_4 _13426_ (.A1(_04767_),
    .A2(_04769_),
    .B1(_04918_),
    .Y(_04919_));
 sky130_fd_sc_hd__and3_1 _13427_ (.A(_04767_),
    .B(_04769_),
    .C(_04918_),
    .X(_04920_));
 sky130_fd_sc_hd__nor3b_4 _13428_ (.A(_04919_),
    .B(_04920_),
    .C_N(_04908_),
    .Y(_04921_));
 sky130_fd_sc_hd__o21ba_1 _13429_ (.A1(_04919_),
    .A2(_04920_),
    .B1_N(_04908_),
    .X(_04922_));
 sky130_fd_sc_hd__a211o_2 _13430_ (.A1(_04797_),
    .A2(_04800_),
    .B1(_04921_),
    .C1(_04922_),
    .X(_04923_));
 sky130_fd_sc_hd__o211ai_4 _13431_ (.A1(_04921_),
    .A2(_04922_),
    .B1(_04797_),
    .C1(_04800_),
    .Y(_04924_));
 sky130_fd_sc_hd__o211a_1 _13432_ (.A1(_04772_),
    .A2(_04774_),
    .B1(_04923_),
    .C1(_04924_),
    .X(_04925_));
 sky130_fd_sc_hd__o211ai_4 _13433_ (.A1(_04772_),
    .A2(_04774_),
    .B1(_04923_),
    .C1(_04924_),
    .Y(_04926_));
 sky130_fd_sc_hd__a211oi_2 _13434_ (.A1(_04923_),
    .A2(_04924_),
    .B1(_04772_),
    .C1(_04774_),
    .Y(_04927_));
 sky130_fd_sc_hd__a22o_1 _13435_ (.A1(net512),
    .A2(net397),
    .B1(net392),
    .B2(net517),
    .X(_04928_));
 sky130_fd_sc_hd__nand4_2 _13436_ (.A(net512),
    .B(net517),
    .C(net397),
    .D(net392),
    .Y(_04929_));
 sky130_fd_sc_hd__nand4_1 _13437_ (.A(net521),
    .B(net387),
    .C(_04928_),
    .D(_04929_),
    .Y(_04930_));
 sky130_fd_sc_hd__a22o_1 _13438_ (.A1(net521),
    .A2(net387),
    .B1(_04928_),
    .B2(_04929_),
    .X(_04931_));
 sky130_fd_sc_hd__and2_1 _13439_ (.A(_04930_),
    .B(_04931_),
    .X(_04932_));
 sky130_fd_sc_hd__nand2_1 _13440_ (.A(net508),
    .B(net403),
    .Y(_04933_));
 sky130_fd_sc_hd__a22o_1 _13441_ (.A1(net504),
    .A2(net407),
    .B1(net499),
    .B2(net411),
    .X(_04934_));
 sky130_fd_sc_hd__nand4_1 _13442_ (.A(net504),
    .B(net411),
    .C(net407),
    .D(net499),
    .Y(_04935_));
 sky130_fd_sc_hd__nand2_1 _13443_ (.A(_04934_),
    .B(_04935_),
    .Y(_04936_));
 sky130_fd_sc_hd__xor2_2 _13444_ (.A(_04933_),
    .B(_04936_),
    .X(_04937_));
 sky130_fd_sc_hd__or2_1 _13445_ (.A(_04788_),
    .B(_04789_),
    .X(_04938_));
 sky130_fd_sc_hd__and2_1 _13446_ (.A(_04937_),
    .B(_04938_),
    .X(_04939_));
 sky130_fd_sc_hd__xor2_2 _13447_ (.A(_04937_),
    .B(_04938_),
    .X(_04940_));
 sky130_fd_sc_hd__and2_1 _13448_ (.A(_04932_),
    .B(_04940_),
    .X(_04941_));
 sky130_fd_sc_hd__xnor2_2 _13449_ (.A(_04932_),
    .B(_04940_),
    .Y(_04942_));
 sky130_fd_sc_hd__a21o_4 _13450_ (.A1(_04809_),
    .A2(_04811_),
    .B1(_04942_),
    .X(_04943_));
 sky130_fd_sc_hd__nand3_4 _13451_ (.A(_04809_),
    .B(_04811_),
    .C(_04942_),
    .Y(_04944_));
 sky130_fd_sc_hd__o211a_1 _13452_ (.A1(_04793_),
    .A2(_04795_),
    .B1(_04943_),
    .C1(_04944_),
    .X(_04945_));
 sky130_fd_sc_hd__o211ai_4 _13453_ (.A1(_04793_),
    .A2(_04795_),
    .B1(_04943_),
    .C1(_04944_),
    .Y(_04946_));
 sky130_fd_sc_hd__a211oi_4 _13454_ (.A1(_04943_),
    .A2(_04944_),
    .B1(_04793_),
    .C1(_04795_),
    .Y(_04947_));
 sky130_fd_sc_hd__or2_1 _13455_ (.A(_04805_),
    .B(_04806_),
    .X(_04948_));
 sky130_fd_sc_hd__a31o_1 _13456_ (.A1(net429),
    .A2(net486),
    .A3(_04815_),
    .B1(_04814_),
    .X(_04949_));
 sky130_fd_sc_hd__a22o_1 _13457_ (.A1(net420),
    .A2(net491),
    .B1(net486),
    .B2(net424),
    .X(_04950_));
 sky130_fd_sc_hd__and4_1 _13458_ (.A(net424),
    .B(net420),
    .C(net491),
    .D(net487),
    .X(_04951_));
 sky130_fd_sc_hd__nand4_1 _13459_ (.A(net424),
    .B(net420),
    .C(net491),
    .D(net486),
    .Y(_04952_));
 sky130_fd_sc_hd__a22oi_1 _13460_ (.A1(net416),
    .A2(net495),
    .B1(_04950_),
    .B2(_04952_),
    .Y(_04953_));
 sky130_fd_sc_hd__and4_1 _13461_ (.A(net416),
    .B(net495),
    .C(_04950_),
    .D(_04952_),
    .X(_04954_));
 sky130_fd_sc_hd__or2_1 _13462_ (.A(_04953_),
    .B(_04954_),
    .X(_04955_));
 sky130_fd_sc_hd__and2b_1 _13463_ (.A_N(_04955_),
    .B(_04949_),
    .X(_04956_));
 sky130_fd_sc_hd__xnor2_2 _13464_ (.A(_04949_),
    .B(_04955_),
    .Y(_04957_));
 sky130_fd_sc_hd__and2_1 _13465_ (.A(_04948_),
    .B(_04957_),
    .X(_04958_));
 sky130_fd_sc_hd__xor2_2 _13466_ (.A(_04948_),
    .B(_04957_),
    .X(_04959_));
 sky130_fd_sc_hd__nand2_1 _13467_ (.A(net428),
    .B(net482),
    .Y(_04960_));
 sky130_fd_sc_hd__and4_1 _13468_ (.A(net438),
    .B(net433),
    .C(net478),
    .D(net474),
    .X(_04961_));
 sky130_fd_sc_hd__a22o_1 _13469_ (.A1(net433),
    .A2(net478),
    .B1(net474),
    .B2(net438),
    .X(_04962_));
 sky130_fd_sc_hd__and2b_1 _13470_ (.A_N(_04961_),
    .B(_04962_),
    .X(_04963_));
 sky130_fd_sc_hd__xnor2_2 _13471_ (.A(_04960_),
    .B(_04963_),
    .Y(_04964_));
 sky130_fd_sc_hd__and2_1 _13472_ (.A(net442),
    .B(net470),
    .X(_04965_));
 sky130_fd_sc_hd__nand4_1 _13473_ (.A(net451),
    .B(net447),
    .C(net466),
    .D(net463),
    .Y(_04966_));
 sky130_fd_sc_hd__a22o_1 _13474_ (.A1(net447),
    .A2(net466),
    .B1(net463),
    .B2(net451),
    .X(_04967_));
 sky130_fd_sc_hd__nand3_1 _13475_ (.A(_04965_),
    .B(_04966_),
    .C(_04967_),
    .Y(_04968_));
 sky130_fd_sc_hd__a21o_1 _13476_ (.A1(_04966_),
    .A2(_04967_),
    .B1(_04965_),
    .X(_04969_));
 sky130_fd_sc_hd__a21bo_1 _13477_ (.A1(_04818_),
    .A2(_04820_),
    .B1_N(_04819_),
    .X(_04970_));
 sky130_fd_sc_hd__nand3_1 _13478_ (.A(_04968_),
    .B(_04969_),
    .C(_04970_),
    .Y(_04971_));
 sky130_fd_sc_hd__a21o_1 _13479_ (.A1(_04968_),
    .A2(_04969_),
    .B1(_04970_),
    .X(_04972_));
 sky130_fd_sc_hd__nand3_2 _13480_ (.A(_04964_),
    .B(_04971_),
    .C(_04972_),
    .Y(_04973_));
 sky130_fd_sc_hd__a21o_1 _13481_ (.A1(_04971_),
    .A2(_04972_),
    .B1(_04964_),
    .X(_04974_));
 sky130_fd_sc_hd__a21bo_1 _13482_ (.A1(_04817_),
    .A2(_04825_),
    .B1_N(_04824_),
    .X(_04975_));
 sky130_fd_sc_hd__nand3_4 _13483_ (.A(_04973_),
    .B(_04974_),
    .C(_04975_),
    .Y(_04976_));
 sky130_fd_sc_hd__a21o_1 _13484_ (.A1(_04973_),
    .A2(_04974_),
    .B1(_04975_),
    .X(_04977_));
 sky130_fd_sc_hd__and3_1 _13485_ (.A(_04959_),
    .B(_04976_),
    .C(_04977_),
    .X(_04978_));
 sky130_fd_sc_hd__nand3_2 _13486_ (.A(_04959_),
    .B(_04976_),
    .C(_04977_),
    .Y(_04979_));
 sky130_fd_sc_hd__a21oi_2 _13487_ (.A1(_04976_),
    .A2(_04977_),
    .B1(_04959_),
    .Y(_04980_));
 sky130_fd_sc_hd__a211oi_4 _13488_ (.A1(_04829_),
    .A2(_04832_),
    .B1(_04978_),
    .C1(_04980_),
    .Y(_04981_));
 sky130_fd_sc_hd__o211a_1 _13489_ (.A1(_04978_),
    .A2(_04980_),
    .B1(_04829_),
    .C1(_04832_),
    .X(_04982_));
 sky130_fd_sc_hd__nor4_2 _13490_ (.A(_04945_),
    .B(_04947_),
    .C(_04981_),
    .D(_04982_),
    .Y(_04983_));
 sky130_fd_sc_hd__or4_2 _13491_ (.A(_04945_),
    .B(_04947_),
    .C(_04981_),
    .D(_04982_),
    .X(_04984_));
 sky130_fd_sc_hd__o22ai_4 _13492_ (.A1(_04945_),
    .A2(_04947_),
    .B1(_04981_),
    .B2(_04982_),
    .Y(_04985_));
 sky130_fd_sc_hd__o211a_2 _13493_ (.A1(_04834_),
    .A2(_04836_),
    .B1(_04984_),
    .C1(_04985_),
    .X(_04986_));
 sky130_fd_sc_hd__a211oi_4 _13494_ (.A1(_04984_),
    .A2(_04985_),
    .B1(_04834_),
    .C1(_04836_),
    .Y(_04987_));
 sky130_fd_sc_hd__nor4_1 _13495_ (.A(_04925_),
    .B(_04927_),
    .C(_04986_),
    .D(_04987_),
    .Y(_04988_));
 sky130_fd_sc_hd__or4_2 _13496_ (.A(_04925_),
    .B(_04927_),
    .C(_04986_),
    .D(_04987_),
    .X(_04989_));
 sky130_fd_sc_hd__o22ai_4 _13497_ (.A1(_04925_),
    .A2(_04927_),
    .B1(_04986_),
    .B2(_04987_),
    .Y(_04990_));
 sky130_fd_sc_hd__o211ai_4 _13498_ (.A1(_04839_),
    .A2(_04841_),
    .B1(_04989_),
    .C1(_04990_),
    .Y(_04991_));
 sky130_fd_sc_hd__a211o_1 _13499_ (.A1(_04989_),
    .A2(_04990_),
    .B1(_04839_),
    .C1(_04841_),
    .X(_04992_));
 sky130_fd_sc_hd__and4bb_1 _13500_ (.A_N(_04892_),
    .B_N(_04893_),
    .C(_04991_),
    .D(_04992_),
    .X(_04993_));
 sky130_fd_sc_hd__or4bb_2 _13501_ (.A(_04892_),
    .B(_04893_),
    .C_N(_04991_),
    .D_N(_04992_),
    .X(_04994_));
 sky130_fd_sc_hd__a2bb2oi_1 _13502_ (.A1_N(_04892_),
    .A2_N(_04893_),
    .B1(_04991_),
    .B2(_04992_),
    .Y(_04995_));
 sky130_fd_sc_hd__a211oi_1 _13503_ (.A1(_04844_),
    .A2(_04847_),
    .B1(_04993_),
    .C1(_04995_),
    .Y(_04996_));
 sky130_fd_sc_hd__a211o_1 _13504_ (.A1(_04844_),
    .A2(_04847_),
    .B1(_04993_),
    .C1(_04995_),
    .X(_04997_));
 sky130_fd_sc_hd__o211a_1 _13505_ (.A1(_04993_),
    .A2(_04995_),
    .B1(_04844_),
    .C1(_04847_),
    .X(_04998_));
 sky130_fd_sc_hd__a211o_1 _13506_ (.A1(_04742_),
    .A2(_04745_),
    .B1(_04996_),
    .C1(_04998_),
    .X(_04999_));
 sky130_fd_sc_hd__o211ai_1 _13507_ (.A1(_04996_),
    .A2(_04998_),
    .B1(_04742_),
    .C1(_04745_),
    .Y(_05000_));
 sky130_fd_sc_hd__nand2_2 _13508_ (.A(_04999_),
    .B(_05000_),
    .Y(_05001_));
 sky130_fd_sc_hd__nor2_2 _13509_ (.A(_04849_),
    .B(_04851_),
    .Y(_05002_));
 sky130_fd_sc_hd__or2_2 _13510_ (.A(_05001_),
    .B(_05002_),
    .X(_05003_));
 sky130_fd_sc_hd__xor2_4 _13511_ (.A(_05001_),
    .B(_05002_),
    .X(_05004_));
 sky130_fd_sc_hd__xnor2_4 _13512_ (.A(_04853_),
    .B(_05004_),
    .Y(_05005_));
 sky130_fd_sc_hd__xnor2_4 _13513_ (.A(_04865_),
    .B(_05005_),
    .Y(_05006_));
 sky130_fd_sc_hd__nor2_1 _13514_ (.A(net9),
    .B(_05006_),
    .Y(_05007_));
 sky130_fd_sc_hd__a221o_1 _13515_ (.A1(net600),
    .A2(net782),
    .B1(_02751_),
    .B2(net6),
    .C1(_05007_),
    .X(_05008_));
 sky130_fd_sc_hd__mux2_1 _13516_ (.A0(net734),
    .A1(_05008_),
    .S(net2),
    .X(_00277_));
 sky130_fd_sc_hd__nor2_1 _13517_ (.A(_04857_),
    .B(_05005_),
    .Y(_05009_));
 sky130_fd_sc_hd__or4_1 _13518_ (.A(_04587_),
    .B(_04718_),
    .C(_04857_),
    .D(_05005_),
    .X(_05010_));
 sky130_fd_sc_hd__o21bai_1 _13519_ (.A1(_04715_),
    .A2(_04854_),
    .B1_N(_04853_),
    .Y(_05011_));
 sky130_fd_sc_hd__nand2_1 _13520_ (.A(_05004_),
    .B(_05011_),
    .Y(_05012_));
 sky130_fd_sc_hd__o31ai_4 _13521_ (.A1(_04857_),
    .A2(_04859_),
    .A3(_05005_),
    .B1(_05012_),
    .Y(_05013_));
 sky130_fd_sc_hd__a31oi_4 _13522_ (.A1(_04456_),
    .A2(_04860_),
    .A3(_05009_),
    .B1(_05013_),
    .Y(_05014_));
 sky130_fd_sc_hd__nor2_1 _13523_ (.A(_04890_),
    .B(_04892_),
    .Y(_05015_));
 sky130_fd_sc_hd__a22oi_2 _13524_ (.A1(net580),
    .A2(net336),
    .B1(net333),
    .B2(net583),
    .Y(_05016_));
 sky130_fd_sc_hd__and4_1 _13525_ (.A(net580),
    .B(net584),
    .C(net336),
    .D(net333),
    .X(_05017_));
 sky130_fd_sc_hd__inv_2 _13526_ (.A(_05017_),
    .Y(_05018_));
 sky130_fd_sc_hd__or2_1 _13527_ (.A(_04872_),
    .B(_04874_),
    .X(_05019_));
 sky130_fd_sc_hd__a22oi_1 _13528_ (.A1(net562),
    .A2(net344),
    .B1(net340),
    .B2(net568),
    .Y(_05020_));
 sky130_fd_sc_hd__and4_1 _13529_ (.A(net562),
    .B(net568),
    .C(net344),
    .D(net340),
    .X(_05021_));
 sky130_fd_sc_hd__o2bb2a_1 _13530_ (.A1_N(net573),
    .A2_N(net337),
    .B1(_05020_),
    .B2(_05021_),
    .X(_05022_));
 sky130_fd_sc_hd__and4bb_1 _13531_ (.A_N(_05020_),
    .B_N(_05021_),
    .C(net573),
    .D(net337),
    .X(_05023_));
 sky130_fd_sc_hd__a211o_1 _13532_ (.A1(_04895_),
    .A2(_04897_),
    .B1(_05022_),
    .C1(_05023_),
    .X(_05024_));
 sky130_fd_sc_hd__o211ai_1 _13533_ (.A1(_05022_),
    .A2(_05023_),
    .B1(_04895_),
    .C1(_04897_),
    .Y(_05025_));
 sky130_fd_sc_hd__and2_1 _13534_ (.A(_05024_),
    .B(_05025_),
    .X(_05026_));
 sky130_fd_sc_hd__nand2_1 _13535_ (.A(_05019_),
    .B(_05026_),
    .Y(_05027_));
 sky130_fd_sc_hd__xnor2_1 _13536_ (.A(_05019_),
    .B(_05026_),
    .Y(_05028_));
 sky130_fd_sc_hd__a21oi_2 _13537_ (.A1(_04905_),
    .A2(_04907_),
    .B1(_05028_),
    .Y(_05029_));
 sky130_fd_sc_hd__inv_2 _13538_ (.A(_05029_),
    .Y(_05030_));
 sky130_fd_sc_hd__and3_1 _13539_ (.A(_04905_),
    .B(_04907_),
    .C(_05028_),
    .X(_05031_));
 sky130_fd_sc_hd__a211oi_2 _13540_ (.A1(_04876_),
    .A2(_04878_),
    .B1(_05029_),
    .C1(_05031_),
    .Y(_05032_));
 sky130_fd_sc_hd__a211o_1 _13541_ (.A1(_04876_),
    .A2(_04878_),
    .B1(_05029_),
    .C1(_05031_),
    .X(_05033_));
 sky130_fd_sc_hd__o211a_1 _13542_ (.A1(_05029_),
    .A2(_05031_),
    .B1(_04876_),
    .C1(_04878_),
    .X(_05034_));
 sky130_fd_sc_hd__a211oi_2 _13543_ (.A1(_04880_),
    .A2(_04882_),
    .B1(_05032_),
    .C1(_05034_),
    .Y(_05035_));
 sky130_fd_sc_hd__o211a_1 _13544_ (.A1(_05032_),
    .A2(_05034_),
    .B1(_04880_),
    .C1(_04882_),
    .X(_05036_));
 sky130_fd_sc_hd__nor4_2 _13545_ (.A(_05016_),
    .B(_05017_),
    .C(_05035_),
    .D(_05036_),
    .Y(_05037_));
 sky130_fd_sc_hd__o22a_1 _13546_ (.A1(_05016_),
    .A2(_05017_),
    .B1(_05035_),
    .B2(_05036_),
    .X(_05038_));
 sky130_fd_sc_hd__a211oi_4 _13547_ (.A1(_04923_),
    .A2(_04926_),
    .B1(_05037_),
    .C1(_05038_),
    .Y(_05039_));
 sky130_fd_sc_hd__inv_2 _13548_ (.A(_05039_),
    .Y(_05040_));
 sky130_fd_sc_hd__o211a_1 _13549_ (.A1(_05037_),
    .A2(_05038_),
    .B1(_04923_),
    .C1(_04926_),
    .X(_05041_));
 sky130_fd_sc_hd__a211oi_2 _13550_ (.A1(_04885_),
    .A2(_04888_),
    .B1(_05039_),
    .C1(_05041_),
    .Y(_05042_));
 sky130_fd_sc_hd__a211o_1 _13551_ (.A1(_04885_),
    .A2(_04888_),
    .B1(_05039_),
    .C1(_05041_),
    .X(_05043_));
 sky130_fd_sc_hd__o211a_1 _13552_ (.A1(_05039_),
    .A2(_05041_),
    .B1(_04885_),
    .C1(_04888_),
    .X(_05044_));
 sky130_fd_sc_hd__a22o_1 _13553_ (.A1(net550),
    .A2(net356),
    .B1(net355),
    .B2(net554),
    .X(_05045_));
 sky130_fd_sc_hd__nand4_2 _13554_ (.A(net550),
    .B(net554),
    .C(net356),
    .D(net354),
    .Y(_05046_));
 sky130_fd_sc_hd__a22o_1 _13555_ (.A1(net558),
    .A2(net348),
    .B1(_05045_),
    .B2(_05046_),
    .X(_05047_));
 sky130_fd_sc_hd__nand4_2 _13556_ (.A(net558),
    .B(net348),
    .C(_05045_),
    .D(_05046_),
    .Y(_05048_));
 sky130_fd_sc_hd__nand2_1 _13557_ (.A(_05047_),
    .B(_05048_),
    .Y(_05049_));
 sky130_fd_sc_hd__a22oi_1 _13558_ (.A1(net537),
    .A2(net632),
    .B1(net367),
    .B2(net542),
    .Y(_05050_));
 sky130_fd_sc_hd__and4_1 _13559_ (.A(net537),
    .B(net542),
    .C(net632),
    .D(net367),
    .X(_05051_));
 sky130_fd_sc_hd__o2bb2a_1 _13560_ (.A1_N(net546),
    .A2_N(net363),
    .B1(_05050_),
    .B2(_05051_),
    .X(_05052_));
 sky130_fd_sc_hd__and4bb_1 _13561_ (.A_N(_05050_),
    .B_N(_05051_),
    .C(\mul0.a[8] ),
    .D(net363),
    .X(_05053_));
 sky130_fd_sc_hd__or2_1 _13562_ (.A(_05052_),
    .B(_05053_),
    .X(_05054_));
 sky130_fd_sc_hd__o21ai_1 _13563_ (.A1(_04899_),
    .A2(_04902_),
    .B1(_04901_),
    .Y(_05055_));
 sky130_fd_sc_hd__nand2b_1 _13564_ (.A_N(_05054_),
    .B(_05055_),
    .Y(_05056_));
 sky130_fd_sc_hd__xor2_1 _13565_ (.A(_05054_),
    .B(_05055_),
    .X(_05057_));
 sky130_fd_sc_hd__or2_1 _13566_ (.A(_05049_),
    .B(_05057_),
    .X(_05058_));
 sky130_fd_sc_hd__nand2_1 _13567_ (.A(_05049_),
    .B(_05057_),
    .Y(_05059_));
 sky130_fd_sc_hd__and2_1 _13568_ (.A(_05058_),
    .B(_05059_),
    .X(_05060_));
 sky130_fd_sc_hd__or2_1 _13569_ (.A(_04911_),
    .B(_04913_),
    .X(_05061_));
 sky130_fd_sc_hd__a22oi_1 _13570_ (.A1(net521),
    .A2(net383),
    .B1(net377),
    .B2(net527),
    .Y(_05062_));
 sky130_fd_sc_hd__and4_1 _13571_ (.A(net524),
    .B(net527),
    .C(net383),
    .D(net377),
    .X(_05063_));
 sky130_fd_sc_hd__o2bb2a_1 _13572_ (.A1_N(net532),
    .A2_N(net374),
    .B1(_05062_),
    .B2(_05063_),
    .X(_05064_));
 sky130_fd_sc_hd__and4bb_1 _13573_ (.A_N(_05062_),
    .B_N(_05063_),
    .C(net532),
    .D(net370),
    .X(_05065_));
 sky130_fd_sc_hd__a211o_1 _13574_ (.A1(_04929_),
    .A2(_04930_),
    .B1(_05064_),
    .C1(_05065_),
    .X(_05066_));
 sky130_fd_sc_hd__o211ai_1 _13575_ (.A1(_05064_),
    .A2(_05065_),
    .B1(_04929_),
    .C1(_04930_),
    .Y(_05067_));
 sky130_fd_sc_hd__and2_1 _13576_ (.A(_05066_),
    .B(_05067_),
    .X(_05068_));
 sky130_fd_sc_hd__nand2_1 _13577_ (.A(_05061_),
    .B(_05068_),
    .Y(_05069_));
 sky130_fd_sc_hd__xnor2_2 _13578_ (.A(_05061_),
    .B(_05068_),
    .Y(_05070_));
 sky130_fd_sc_hd__a21oi_4 _13579_ (.A1(_04914_),
    .A2(_04917_),
    .B1(_05070_),
    .Y(_05071_));
 sky130_fd_sc_hd__and3_1 _13580_ (.A(_04914_),
    .B(_04917_),
    .C(_05070_),
    .X(_05072_));
 sky130_fd_sc_hd__nor3b_4 _13581_ (.A(_05071_),
    .B(_05072_),
    .C_N(_05060_),
    .Y(_05073_));
 sky130_fd_sc_hd__o21ba_1 _13582_ (.A1(_05071_),
    .A2(_05072_),
    .B1_N(_05060_),
    .X(_05074_));
 sky130_fd_sc_hd__a211o_2 _13583_ (.A1(_04943_),
    .A2(_04946_),
    .B1(_05073_),
    .C1(_05074_),
    .X(_05075_));
 sky130_fd_sc_hd__o211ai_4 _13584_ (.A1(_05073_),
    .A2(_05074_),
    .B1(_04943_),
    .C1(_04946_),
    .Y(_05076_));
 sky130_fd_sc_hd__o211a_1 _13585_ (.A1(_04919_),
    .A2(_04921_),
    .B1(_05075_),
    .C1(_05076_),
    .X(_05077_));
 sky130_fd_sc_hd__o211ai_2 _13586_ (.A1(_04919_),
    .A2(_04921_),
    .B1(_05075_),
    .C1(_05076_),
    .Y(_05078_));
 sky130_fd_sc_hd__a211oi_2 _13587_ (.A1(_05075_),
    .A2(_05076_),
    .B1(_04919_),
    .C1(_04921_),
    .Y(_05079_));
 sky130_fd_sc_hd__a22o_1 _13588_ (.A1(net508),
    .A2(net397),
    .B1(net392),
    .B2(net512),
    .X(_05080_));
 sky130_fd_sc_hd__nand4_2 _13589_ (.A(\mul0.a[16] ),
    .B(net512),
    .C(net397),
    .D(net392),
    .Y(_05081_));
 sky130_fd_sc_hd__a22o_1 _13590_ (.A1(net517),
    .A2(net387),
    .B1(_05080_),
    .B2(_05081_),
    .X(_05082_));
 sky130_fd_sc_hd__nand4_2 _13591_ (.A(net517),
    .B(net387),
    .C(_05080_),
    .D(_05081_),
    .Y(_05083_));
 sky130_fd_sc_hd__nand2_1 _13592_ (.A(_05082_),
    .B(_05083_),
    .Y(_05084_));
 sky130_fd_sc_hd__a22oi_1 _13593_ (.A1(net407),
    .A2(net499),
    .B1(net495),
    .B2(net411),
    .Y(_05085_));
 sky130_fd_sc_hd__and4_1 _13594_ (.A(net411),
    .B(net407),
    .C(net499),
    .D(net495),
    .X(_05086_));
 sky130_fd_sc_hd__o2bb2a_1 _13595_ (.A1_N(net504),
    .A2_N(net403),
    .B1(_05085_),
    .B2(_05086_),
    .X(_05087_));
 sky130_fd_sc_hd__and4bb_1 _13596_ (.A_N(_05085_),
    .B_N(_05086_),
    .C(net504),
    .D(net403),
    .X(_05088_));
 sky130_fd_sc_hd__or2_1 _13597_ (.A(_05087_),
    .B(_05088_),
    .X(_05089_));
 sky130_fd_sc_hd__o21ai_1 _13598_ (.A1(_04933_),
    .A2(_04936_),
    .B1(_04935_),
    .Y(_05090_));
 sky130_fd_sc_hd__nand2b_1 _13599_ (.A_N(_05089_),
    .B(_05090_),
    .Y(_05091_));
 sky130_fd_sc_hd__xor2_1 _13600_ (.A(_05089_),
    .B(_05090_),
    .X(_05092_));
 sky130_fd_sc_hd__or2_1 _13601_ (.A(_05084_),
    .B(_05092_),
    .X(_05093_));
 sky130_fd_sc_hd__xor2_1 _13602_ (.A(_05084_),
    .B(_05092_),
    .X(_05094_));
 sky130_fd_sc_hd__o21a_1 _13603_ (.A1(_04956_),
    .A2(_04958_),
    .B1(_05094_),
    .X(_05095_));
 sky130_fd_sc_hd__o21ai_2 _13604_ (.A1(_04956_),
    .A2(_04958_),
    .B1(_05094_),
    .Y(_05096_));
 sky130_fd_sc_hd__or3_2 _13605_ (.A(_04956_),
    .B(_04958_),
    .C(_05094_),
    .X(_05097_));
 sky130_fd_sc_hd__o211a_2 _13606_ (.A1(_04939_),
    .A2(_04941_),
    .B1(_05096_),
    .C1(_05097_),
    .X(_05098_));
 sky130_fd_sc_hd__a211oi_4 _13607_ (.A1(_05096_),
    .A2(_05097_),
    .B1(_04939_),
    .C1(_04941_),
    .Y(_05099_));
 sky130_fd_sc_hd__nor2_1 _13608_ (.A(_04951_),
    .B(_04954_),
    .Y(_05100_));
 sky130_fd_sc_hd__a31o_1 _13609_ (.A1(net428),
    .A2(net483),
    .A3(_04962_),
    .B1(_04961_),
    .X(_05101_));
 sky130_fd_sc_hd__a22o_1 _13610_ (.A1(net419),
    .A2(net487),
    .B1(net483),
    .B2(net423),
    .X(_05102_));
 sky130_fd_sc_hd__nand4_1 _13611_ (.A(net423),
    .B(net419),
    .C(net487),
    .D(net483),
    .Y(_05103_));
 sky130_fd_sc_hd__a22oi_1 _13612_ (.A1(net416),
    .A2(net491),
    .B1(_05102_),
    .B2(_05103_),
    .Y(_05104_));
 sky130_fd_sc_hd__and4_1 _13613_ (.A(net416),
    .B(net491),
    .C(_05102_),
    .D(_05103_),
    .X(_05105_));
 sky130_fd_sc_hd__or2_1 _13614_ (.A(_05104_),
    .B(_05105_),
    .X(_05106_));
 sky130_fd_sc_hd__and2b_1 _13615_ (.A_N(_05106_),
    .B(_05101_),
    .X(_05107_));
 sky130_fd_sc_hd__xnor2_2 _13616_ (.A(_05101_),
    .B(_05106_),
    .Y(_05108_));
 sky130_fd_sc_hd__and2b_1 _13617_ (.A_N(_05100_),
    .B(_05108_),
    .X(_05109_));
 sky130_fd_sc_hd__xnor2_2 _13618_ (.A(_05100_),
    .B(_05108_),
    .Y(_05110_));
 sky130_fd_sc_hd__nand2_1 _13619_ (.A(net428),
    .B(net478),
    .Y(_05111_));
 sky130_fd_sc_hd__and4_1 _13620_ (.A(net438),
    .B(net433),
    .C(net474),
    .D(net470),
    .X(_05112_));
 sky130_fd_sc_hd__a22o_1 _13621_ (.A1(net433),
    .A2(net474),
    .B1(net470),
    .B2(net438),
    .X(_05113_));
 sky130_fd_sc_hd__and2b_1 _13622_ (.A_N(_05112_),
    .B(_05113_),
    .X(_05114_));
 sky130_fd_sc_hd__xnor2_2 _13623_ (.A(_05111_),
    .B(_05114_),
    .Y(_05115_));
 sky130_fd_sc_hd__and2_1 _13624_ (.A(net442),
    .B(net466),
    .X(_05116_));
 sky130_fd_sc_hd__nand4_1 _13625_ (.A(net451),
    .B(net447),
    .C(net463),
    .D(net460),
    .Y(_05117_));
 sky130_fd_sc_hd__a22o_1 _13626_ (.A1(net447),
    .A2(net463),
    .B1(net460),
    .B2(net451),
    .X(_05118_));
 sky130_fd_sc_hd__nand3_1 _13627_ (.A(_05116_),
    .B(_05117_),
    .C(_05118_),
    .Y(_05119_));
 sky130_fd_sc_hd__a21o_1 _13628_ (.A1(_05117_),
    .A2(_05118_),
    .B1(_05116_),
    .X(_05120_));
 sky130_fd_sc_hd__a21bo_1 _13629_ (.A1(_04965_),
    .A2(_04967_),
    .B1_N(_04966_),
    .X(_05121_));
 sky130_fd_sc_hd__nand3_1 _13630_ (.A(_05119_),
    .B(_05120_),
    .C(_05121_),
    .Y(_05122_));
 sky130_fd_sc_hd__a21o_1 _13631_ (.A1(_05119_),
    .A2(_05120_),
    .B1(_05121_),
    .X(_05123_));
 sky130_fd_sc_hd__nand3_2 _13632_ (.A(_05115_),
    .B(_05122_),
    .C(_05123_),
    .Y(_05124_));
 sky130_fd_sc_hd__a21o_1 _13633_ (.A1(_05122_),
    .A2(_05123_),
    .B1(_05115_),
    .X(_05125_));
 sky130_fd_sc_hd__a21bo_1 _13634_ (.A1(_04964_),
    .A2(_04972_),
    .B1_N(_04971_),
    .X(_05126_));
 sky130_fd_sc_hd__nand3_4 _13635_ (.A(_05124_),
    .B(_05125_),
    .C(_05126_),
    .Y(_05127_));
 sky130_fd_sc_hd__a21o_1 _13636_ (.A1(_05124_),
    .A2(_05125_),
    .B1(_05126_),
    .X(_05128_));
 sky130_fd_sc_hd__and3_1 _13637_ (.A(_05110_),
    .B(_05127_),
    .C(_05128_),
    .X(_05129_));
 sky130_fd_sc_hd__nand3_2 _13638_ (.A(_05110_),
    .B(_05127_),
    .C(_05128_),
    .Y(_05130_));
 sky130_fd_sc_hd__a21oi_2 _13639_ (.A1(_05127_),
    .A2(_05128_),
    .B1(_05110_),
    .Y(_05131_));
 sky130_fd_sc_hd__a211oi_4 _13640_ (.A1(_04976_),
    .A2(_04979_),
    .B1(_05129_),
    .C1(_05131_),
    .Y(_05132_));
 sky130_fd_sc_hd__o211a_1 _13641_ (.A1(_05129_),
    .A2(_05131_),
    .B1(_04976_),
    .C1(_04979_),
    .X(_05133_));
 sky130_fd_sc_hd__nor4_2 _13642_ (.A(_05098_),
    .B(_05099_),
    .C(_05132_),
    .D(_05133_),
    .Y(_05134_));
 sky130_fd_sc_hd__or4_2 _13643_ (.A(_05098_),
    .B(_05099_),
    .C(_05132_),
    .D(_05133_),
    .X(_05135_));
 sky130_fd_sc_hd__o22ai_4 _13644_ (.A1(_05098_),
    .A2(_05099_),
    .B1(_05132_),
    .B2(_05133_),
    .Y(_05136_));
 sky130_fd_sc_hd__o211a_2 _13645_ (.A1(_04981_),
    .A2(_04983_),
    .B1(_05135_),
    .C1(_05136_),
    .X(_05137_));
 sky130_fd_sc_hd__a211oi_4 _13646_ (.A1(_05135_),
    .A2(_05136_),
    .B1(_04981_),
    .C1(_04983_),
    .Y(_05138_));
 sky130_fd_sc_hd__nor4_2 _13647_ (.A(_05077_),
    .B(_05079_),
    .C(_05137_),
    .D(_05138_),
    .Y(_05139_));
 sky130_fd_sc_hd__or4_1 _13648_ (.A(_05077_),
    .B(_05079_),
    .C(_05137_),
    .D(_05138_),
    .X(_05140_));
 sky130_fd_sc_hd__o22ai_2 _13649_ (.A1(_05077_),
    .A2(_05079_),
    .B1(_05137_),
    .B2(_05138_),
    .Y(_05141_));
 sky130_fd_sc_hd__o211a_2 _13650_ (.A1(_04986_),
    .A2(_04988_),
    .B1(_05140_),
    .C1(_05141_),
    .X(_05142_));
 sky130_fd_sc_hd__a211oi_2 _13651_ (.A1(_05140_),
    .A2(_05141_),
    .B1(_04986_),
    .C1(_04988_),
    .Y(_05143_));
 sky130_fd_sc_hd__nor4_4 _13652_ (.A(_05042_),
    .B(_05044_),
    .C(_05142_),
    .D(_05143_),
    .Y(_05144_));
 sky130_fd_sc_hd__o22a_1 _13653_ (.A1(_05042_),
    .A2(_05044_),
    .B1(_05142_),
    .B2(_05143_),
    .X(_05145_));
 sky130_fd_sc_hd__a211oi_4 _13654_ (.A1(_04991_),
    .A2(_04994_),
    .B1(_05144_),
    .C1(_05145_),
    .Y(_05146_));
 sky130_fd_sc_hd__o211a_1 _13655_ (.A1(_05144_),
    .A2(_05145_),
    .B1(_04991_),
    .C1(_04994_),
    .X(_05147_));
 sky130_fd_sc_hd__nor3_2 _13656_ (.A(_05015_),
    .B(_05146_),
    .C(_05147_),
    .Y(_05148_));
 sky130_fd_sc_hd__o21a_1 _13657_ (.A1(_05146_),
    .A2(_05147_),
    .B1(_05015_),
    .X(_05149_));
 sky130_fd_sc_hd__a211o_2 _13658_ (.A1(_04997_),
    .A2(_04999_),
    .B1(_05148_),
    .C1(_05149_),
    .X(_05150_));
 sky130_fd_sc_hd__o211ai_2 _13659_ (.A1(_05148_),
    .A2(_05149_),
    .B1(_04997_),
    .C1(_04999_),
    .Y(_05151_));
 sky130_fd_sc_hd__and2_2 _13660_ (.A(_05150_),
    .B(_05151_),
    .X(_05152_));
 sky130_fd_sc_hd__nand2b_1 _13661_ (.A_N(_05003_),
    .B(_05152_),
    .Y(_05153_));
 sky130_fd_sc_hd__xnor2_4 _13662_ (.A(_05003_),
    .B(_05152_),
    .Y(_05154_));
 sky130_fd_sc_hd__nand2b_1 _13663_ (.A_N(_05014_),
    .B(_05154_),
    .Y(_05155_));
 sky130_fd_sc_hd__xor2_4 _13664_ (.A(_05014_),
    .B(_05154_),
    .X(_05156_));
 sky130_fd_sc_hd__nor2_1 _13665_ (.A(_03057_),
    .B(_05156_),
    .Y(_05157_));
 sky130_fd_sc_hd__a221o_1 _13666_ (.A1(net600),
    .A2(net740),
    .B1(_02619_),
    .B2(net5),
    .C1(_05157_),
    .X(_05158_));
 sky130_fd_sc_hd__mux2_1 _13667_ (.A0(net697),
    .A1(_05158_),
    .S(net1),
    .X(_00278_));
 sky130_fd_sc_hd__nand2_2 _13668_ (.A(_05153_),
    .B(_05155_),
    .Y(_05159_));
 sky130_fd_sc_hd__nor2_1 _13669_ (.A(_05035_),
    .B(_05037_),
    .Y(_05160_));
 sky130_fd_sc_hd__a22o_1 _13670_ (.A1(net574),
    .A2(net336),
    .B1(net333),
    .B2(net578),
    .X(_05161_));
 sky130_fd_sc_hd__and3_1 _13671_ (.A(net574),
    .B(net578),
    .C(net333),
    .X(_05162_));
 sky130_fd_sc_hd__a21bo_1 _13672_ (.A1(net336),
    .A2(_05162_),
    .B1_N(_05161_),
    .X(_05163_));
 sky130_fd_sc_hd__nand2_1 _13673_ (.A(net584),
    .B(net330),
    .Y(_05164_));
 sky130_fd_sc_hd__xnor2_1 _13674_ (.A(_05163_),
    .B(_05164_),
    .Y(_05165_));
 sky130_fd_sc_hd__nor2_1 _13675_ (.A(_05018_),
    .B(_05165_),
    .Y(_05166_));
 sky130_fd_sc_hd__and2_1 _13676_ (.A(_05018_),
    .B(_05165_),
    .X(_05167_));
 sky130_fd_sc_hd__or2_1 _13677_ (.A(_05166_),
    .B(_05167_),
    .X(_05168_));
 sky130_fd_sc_hd__or2_1 _13678_ (.A(_05021_),
    .B(_05023_),
    .X(_05169_));
 sky130_fd_sc_hd__a22oi_1 _13679_ (.A1(net559),
    .A2(net344),
    .B1(net340),
    .B2(net562),
    .Y(_05170_));
 sky130_fd_sc_hd__and4_1 _13680_ (.A(net559),
    .B(net562),
    .C(net345),
    .D(net341),
    .X(_05171_));
 sky130_fd_sc_hd__o2bb2a_1 _13681_ (.A1_N(net568),
    .A2_N(net337),
    .B1(_05170_),
    .B2(_05171_),
    .X(_05172_));
 sky130_fd_sc_hd__and4bb_1 _13682_ (.A_N(_05170_),
    .B_N(_05171_),
    .C(net568),
    .D(net337),
    .X(_05173_));
 sky130_fd_sc_hd__a211o_1 _13683_ (.A1(_05046_),
    .A2(_05048_),
    .B1(_05172_),
    .C1(_05173_),
    .X(_05174_));
 sky130_fd_sc_hd__o211ai_1 _13684_ (.A1(_05172_),
    .A2(_05173_),
    .B1(_05046_),
    .C1(_05048_),
    .Y(_05175_));
 sky130_fd_sc_hd__and2_1 _13685_ (.A(_05174_),
    .B(_05175_),
    .X(_05176_));
 sky130_fd_sc_hd__nand2_1 _13686_ (.A(_05169_),
    .B(_05176_),
    .Y(_05177_));
 sky130_fd_sc_hd__xnor2_1 _13687_ (.A(_05169_),
    .B(_05176_),
    .Y(_05178_));
 sky130_fd_sc_hd__a21oi_2 _13688_ (.A1(_05056_),
    .A2(_05058_),
    .B1(_05178_),
    .Y(_05179_));
 sky130_fd_sc_hd__inv_2 _13689_ (.A(_05179_),
    .Y(_05180_));
 sky130_fd_sc_hd__and3_1 _13690_ (.A(_05056_),
    .B(_05058_),
    .C(_05178_),
    .X(_05181_));
 sky130_fd_sc_hd__a211oi_2 _13691_ (.A1(_05024_),
    .A2(_05027_),
    .B1(_05179_),
    .C1(_05181_),
    .Y(_05182_));
 sky130_fd_sc_hd__a211o_1 _13692_ (.A1(_05024_),
    .A2(_05027_),
    .B1(_05179_),
    .C1(_05181_),
    .X(_05183_));
 sky130_fd_sc_hd__o211a_1 _13693_ (.A1(_05179_),
    .A2(_05181_),
    .B1(_05024_),
    .C1(_05027_),
    .X(_05184_));
 sky130_fd_sc_hd__a211oi_2 _13694_ (.A1(_05030_),
    .A2(_05033_),
    .B1(_05182_),
    .C1(_05184_),
    .Y(_05185_));
 sky130_fd_sc_hd__inv_2 _13695_ (.A(_05185_),
    .Y(_05186_));
 sky130_fd_sc_hd__o211a_1 _13696_ (.A1(_05182_),
    .A2(_05184_),
    .B1(_05030_),
    .C1(_05033_),
    .X(_05187_));
 sky130_fd_sc_hd__nor3_1 _13697_ (.A(_05168_),
    .B(_05185_),
    .C(_05187_),
    .Y(_05188_));
 sky130_fd_sc_hd__or3_2 _13698_ (.A(_05168_),
    .B(_05185_),
    .C(_05187_),
    .X(_05189_));
 sky130_fd_sc_hd__o21a_1 _13699_ (.A1(_05185_),
    .A2(_05187_),
    .B1(_05168_),
    .X(_05190_));
 sky130_fd_sc_hd__a211oi_2 _13700_ (.A1(_05075_),
    .A2(_05078_),
    .B1(_05188_),
    .C1(_05190_),
    .Y(_05191_));
 sky130_fd_sc_hd__o211a_1 _13701_ (.A1(_05188_),
    .A2(_05190_),
    .B1(_05075_),
    .C1(_05078_),
    .X(_05192_));
 sky130_fd_sc_hd__nor3_1 _13702_ (.A(_05160_),
    .B(_05191_),
    .C(_05192_),
    .Y(_05193_));
 sky130_fd_sc_hd__o21a_1 _13703_ (.A1(_05191_),
    .A2(_05192_),
    .B1(_05160_),
    .X(_05194_));
 sky130_fd_sc_hd__a22o_1 _13704_ (.A1(net546),
    .A2(net356),
    .B1(net355),
    .B2(net551),
    .X(_05195_));
 sky130_fd_sc_hd__nand4_2 _13705_ (.A(net546),
    .B(net550),
    .C(net356),
    .D(net354),
    .Y(_05196_));
 sky130_fd_sc_hd__a22o_1 _13706_ (.A1(net555),
    .A2(net348),
    .B1(_05195_),
    .B2(_05196_),
    .X(_05197_));
 sky130_fd_sc_hd__nand4_1 _13707_ (.A(net555),
    .B(net348),
    .C(_05195_),
    .D(_05196_),
    .Y(_05198_));
 sky130_fd_sc_hd__nand2_1 _13708_ (.A(_05197_),
    .B(_05198_),
    .Y(_05199_));
 sky130_fd_sc_hd__a22oi_1 _13709_ (.A1(net532),
    .A2(net632),
    .B1(net367),
    .B2(net537),
    .Y(_05200_));
 sky130_fd_sc_hd__and4_1 _13710_ (.A(net532),
    .B(net537),
    .C(net632),
    .D(net367),
    .X(_05201_));
 sky130_fd_sc_hd__o2bb2a_1 _13711_ (.A1_N(net542),
    .A2_N(net363),
    .B1(_05200_),
    .B2(_05201_),
    .X(_05202_));
 sky130_fd_sc_hd__and4bb_1 _13712_ (.A_N(_05200_),
    .B_N(_05201_),
    .C(net542),
    .D(net363),
    .X(_05203_));
 sky130_fd_sc_hd__nor2_1 _13713_ (.A(_05202_),
    .B(_05203_),
    .Y(_05204_));
 sky130_fd_sc_hd__or2_1 _13714_ (.A(_05051_),
    .B(_05053_),
    .X(_05205_));
 sky130_fd_sc_hd__nand2_1 _13715_ (.A(_05204_),
    .B(_05205_),
    .Y(_05206_));
 sky130_fd_sc_hd__xnor2_1 _13716_ (.A(_05204_),
    .B(_05205_),
    .Y(_05207_));
 sky130_fd_sc_hd__or2_1 _13717_ (.A(_05199_),
    .B(_05207_),
    .X(_05208_));
 sky130_fd_sc_hd__nand2_1 _13718_ (.A(_05199_),
    .B(_05207_),
    .Y(_05209_));
 sky130_fd_sc_hd__and2_1 _13719_ (.A(_05208_),
    .B(_05209_),
    .X(_05210_));
 sky130_fd_sc_hd__or2_1 _13720_ (.A(_05063_),
    .B(_05065_),
    .X(_05211_));
 sky130_fd_sc_hd__a22o_1 _13721_ (.A1(net517),
    .A2(net383),
    .B1(net377),
    .B2(net524),
    .X(_05212_));
 sky130_fd_sc_hd__nand4_1 _13722_ (.A(net517),
    .B(net524),
    .C(net383),
    .D(net377),
    .Y(_05213_));
 sky130_fd_sc_hd__a22oi_2 _13723_ (.A1(net527),
    .A2(net374),
    .B1(_05212_),
    .B2(_05213_),
    .Y(_05214_));
 sky130_fd_sc_hd__and4_1 _13724_ (.A(net527),
    .B(net374),
    .C(_05212_),
    .D(_05213_),
    .X(_05215_));
 sky130_fd_sc_hd__a211o_1 _13725_ (.A1(_05081_),
    .A2(_05083_),
    .B1(_05214_),
    .C1(_05215_),
    .X(_05216_));
 sky130_fd_sc_hd__o211ai_1 _13726_ (.A1(_05214_),
    .A2(_05215_),
    .B1(_05081_),
    .C1(_05083_),
    .Y(_05217_));
 sky130_fd_sc_hd__and2_1 _13727_ (.A(_05216_),
    .B(_05217_),
    .X(_05218_));
 sky130_fd_sc_hd__nand2_1 _13728_ (.A(_05211_),
    .B(_05218_),
    .Y(_05219_));
 sky130_fd_sc_hd__xnor2_2 _13729_ (.A(_05211_),
    .B(_05218_),
    .Y(_05220_));
 sky130_fd_sc_hd__a21oi_2 _13730_ (.A1(_05066_),
    .A2(_05069_),
    .B1(_05220_),
    .Y(_05221_));
 sky130_fd_sc_hd__a21o_1 _13731_ (.A1(_05066_),
    .A2(_05069_),
    .B1(_05220_),
    .X(_05222_));
 sky130_fd_sc_hd__nand3_1 _13732_ (.A(_05066_),
    .B(_05069_),
    .C(_05220_),
    .Y(_05223_));
 sky130_fd_sc_hd__and3_1 _13733_ (.A(_05210_),
    .B(_05222_),
    .C(_05223_),
    .X(_05224_));
 sky130_fd_sc_hd__nand3_2 _13734_ (.A(_05210_),
    .B(_05222_),
    .C(_05223_),
    .Y(_05225_));
 sky130_fd_sc_hd__a21o_1 _13735_ (.A1(_05222_),
    .A2(_05223_),
    .B1(_05210_),
    .X(_05226_));
 sky130_fd_sc_hd__o211ai_4 _13736_ (.A1(_05095_),
    .A2(_05098_),
    .B1(_05225_),
    .C1(_05226_),
    .Y(_05227_));
 sky130_fd_sc_hd__a211o_2 _13737_ (.A1(_05225_),
    .A2(_05226_),
    .B1(_05095_),
    .C1(_05098_),
    .X(_05228_));
 sky130_fd_sc_hd__o211a_1 _13738_ (.A1(_05071_),
    .A2(_05073_),
    .B1(_05227_),
    .C1(_05228_),
    .X(_05229_));
 sky130_fd_sc_hd__o211ai_4 _13739_ (.A1(_05071_),
    .A2(_05073_),
    .B1(_05227_),
    .C1(_05228_),
    .Y(_05230_));
 sky130_fd_sc_hd__a211oi_2 _13740_ (.A1(_05227_),
    .A2(_05228_),
    .B1(_05071_),
    .C1(_05073_),
    .Y(_05231_));
 sky130_fd_sc_hd__a22o_1 _13741_ (.A1(net504),
    .A2(net397),
    .B1(net392),
    .B2(net508),
    .X(_05232_));
 sky130_fd_sc_hd__and4_1 _13742_ (.A(net504),
    .B(net508),
    .C(net397),
    .D(net392),
    .X(_05233_));
 sky130_fd_sc_hd__inv_2 _13743_ (.A(_05233_),
    .Y(_05234_));
 sky130_fd_sc_hd__nand2_1 _13744_ (.A(_05232_),
    .B(_05234_),
    .Y(_05235_));
 sky130_fd_sc_hd__nand2_1 _13745_ (.A(net512),
    .B(net387),
    .Y(_05236_));
 sky130_fd_sc_hd__xnor2_1 _13746_ (.A(_05235_),
    .B(_05236_),
    .Y(_05237_));
 sky130_fd_sc_hd__a22o_1 _13747_ (.A1(net407),
    .A2(net495),
    .B1(net491),
    .B2(net411),
    .X(_05238_));
 sky130_fd_sc_hd__nand4_4 _13748_ (.A(net411),
    .B(net407),
    .C(net495),
    .D(net491),
    .Y(_05239_));
 sky130_fd_sc_hd__a22o_1 _13749_ (.A1(net403),
    .A2(net499),
    .B1(_05238_),
    .B2(_05239_),
    .X(_05240_));
 sky130_fd_sc_hd__nand4_2 _13750_ (.A(net403),
    .B(net499),
    .C(_05238_),
    .D(_05239_),
    .Y(_05241_));
 sky130_fd_sc_hd__nand2_1 _13751_ (.A(_05240_),
    .B(_05241_),
    .Y(_05242_));
 sky130_fd_sc_hd__or2_1 _13752_ (.A(_05086_),
    .B(_05088_),
    .X(_05243_));
 sky130_fd_sc_hd__nand2b_1 _13753_ (.A_N(_05242_),
    .B(_05243_),
    .Y(_05244_));
 sky130_fd_sc_hd__xor2_1 _13754_ (.A(_05242_),
    .B(_05243_),
    .X(_05245_));
 sky130_fd_sc_hd__or2_1 _13755_ (.A(_05237_),
    .B(_05245_),
    .X(_05246_));
 sky130_fd_sc_hd__xor2_1 _13756_ (.A(_05237_),
    .B(_05245_),
    .X(_05247_));
 sky130_fd_sc_hd__o21a_2 _13757_ (.A1(_05107_),
    .A2(_05109_),
    .B1(_05247_),
    .X(_05248_));
 sky130_fd_sc_hd__nor3_2 _13758_ (.A(_05107_),
    .B(_05109_),
    .C(_05247_),
    .Y(_05249_));
 sky130_fd_sc_hd__a211oi_4 _13759_ (.A1(_05091_),
    .A2(_05093_),
    .B1(_05248_),
    .C1(_05249_),
    .Y(_05250_));
 sky130_fd_sc_hd__o211a_1 _13760_ (.A1(_05248_),
    .A2(_05249_),
    .B1(_05091_),
    .C1(_05093_),
    .X(_05251_));
 sky130_fd_sc_hd__a41o_1 _13761_ (.A1(net423),
    .A2(net419),
    .A3(net487),
    .A4(net482),
    .B1(_05105_),
    .X(_05252_));
 sky130_fd_sc_hd__a31o_1 _13762_ (.A1(net428),
    .A2(net478),
    .A3(_05113_),
    .B1(_05112_),
    .X(_05253_));
 sky130_fd_sc_hd__a22o_1 _13763_ (.A1(net419),
    .A2(net483),
    .B1(net478),
    .B2(net423),
    .X(_05254_));
 sky130_fd_sc_hd__nand4_2 _13764_ (.A(net423),
    .B(net419),
    .C(net483),
    .D(net478),
    .Y(_05255_));
 sky130_fd_sc_hd__a22o_1 _13765_ (.A1(net415),
    .A2(net487),
    .B1(_05254_),
    .B2(_05255_),
    .X(_05256_));
 sky130_fd_sc_hd__nand4_1 _13766_ (.A(net415),
    .B(net487),
    .C(_05254_),
    .D(_05255_),
    .Y(_05257_));
 sky130_fd_sc_hd__and3_1 _13767_ (.A(_05253_),
    .B(_05256_),
    .C(_05257_),
    .X(_05258_));
 sky130_fd_sc_hd__a21o_1 _13768_ (.A1(_05256_),
    .A2(_05257_),
    .B1(_05253_),
    .X(_05259_));
 sky130_fd_sc_hd__and2b_1 _13769_ (.A_N(_05258_),
    .B(_05259_),
    .X(_05260_));
 sky130_fd_sc_hd__xor2_2 _13770_ (.A(_05252_),
    .B(_05260_),
    .X(_05261_));
 sky130_fd_sc_hd__nand2_1 _13771_ (.A(net428),
    .B(net474),
    .Y(_05262_));
 sky130_fd_sc_hd__a22o_1 _13772_ (.A1(net433),
    .A2(net470),
    .B1(net466),
    .B2(net438),
    .X(_05263_));
 sky130_fd_sc_hd__and3_1 _13773_ (.A(net438),
    .B(net433),
    .C(net470),
    .X(_05264_));
 sky130_fd_sc_hd__a21bo_1 _13774_ (.A1(net466),
    .A2(_05264_),
    .B1_N(_05263_),
    .X(_05265_));
 sky130_fd_sc_hd__xor2_1 _13775_ (.A(_05262_),
    .B(_05265_),
    .X(_05266_));
 sky130_fd_sc_hd__and2_1 _13776_ (.A(net442),
    .B(net463),
    .X(_05267_));
 sky130_fd_sc_hd__a22o_1 _13777_ (.A1(net447),
    .A2(net460),
    .B1(net459),
    .B2(net451),
    .X(_05268_));
 sky130_fd_sc_hd__nand4_1 _13778_ (.A(net451),
    .B(net447),
    .C(net460),
    .D(net459),
    .Y(_05269_));
 sky130_fd_sc_hd__nand3_1 _13779_ (.A(_05267_),
    .B(_05268_),
    .C(_05269_),
    .Y(_05270_));
 sky130_fd_sc_hd__a21o_1 _13780_ (.A1(_05268_),
    .A2(_05269_),
    .B1(_05267_),
    .X(_05271_));
 sky130_fd_sc_hd__a21bo_1 _13781_ (.A1(_05116_),
    .A2(_05118_),
    .B1_N(_05117_),
    .X(_05272_));
 sky130_fd_sc_hd__nand3_1 _13782_ (.A(_05270_),
    .B(_05271_),
    .C(_05272_),
    .Y(_05273_));
 sky130_fd_sc_hd__a21o_1 _13783_ (.A1(_05270_),
    .A2(_05271_),
    .B1(_05272_),
    .X(_05274_));
 sky130_fd_sc_hd__nand3_1 _13784_ (.A(_05266_),
    .B(_05273_),
    .C(_05274_),
    .Y(_05275_));
 sky130_fd_sc_hd__a21o_1 _13785_ (.A1(_05273_),
    .A2(_05274_),
    .B1(_05266_),
    .X(_05276_));
 sky130_fd_sc_hd__a21bo_1 _13786_ (.A1(_05115_),
    .A2(_05123_),
    .B1_N(_05122_),
    .X(_05277_));
 sky130_fd_sc_hd__nand3_2 _13787_ (.A(_05275_),
    .B(_05276_),
    .C(_05277_),
    .Y(_05278_));
 sky130_fd_sc_hd__a21o_1 _13788_ (.A1(_05275_),
    .A2(_05276_),
    .B1(_05277_),
    .X(_05279_));
 sky130_fd_sc_hd__and3_1 _13789_ (.A(_05261_),
    .B(_05278_),
    .C(_05279_),
    .X(_05280_));
 sky130_fd_sc_hd__nand3_1 _13790_ (.A(_05261_),
    .B(_05278_),
    .C(_05279_),
    .Y(_05281_));
 sky130_fd_sc_hd__a21oi_2 _13791_ (.A1(_05278_),
    .A2(_05279_),
    .B1(_05261_),
    .Y(_05282_));
 sky130_fd_sc_hd__a211oi_4 _13792_ (.A1(_05127_),
    .A2(_05130_),
    .B1(_05280_),
    .C1(_05282_),
    .Y(_05283_));
 sky130_fd_sc_hd__o211a_2 _13793_ (.A1(_05280_),
    .A2(_05282_),
    .B1(_05127_),
    .C1(_05130_),
    .X(_05284_));
 sky130_fd_sc_hd__nor4_2 _13794_ (.A(_05250_),
    .B(_05251_),
    .C(_05283_),
    .D(_05284_),
    .Y(_05285_));
 sky130_fd_sc_hd__or4_2 _13795_ (.A(_05250_),
    .B(_05251_),
    .C(_05283_),
    .D(_05284_),
    .X(_05286_));
 sky130_fd_sc_hd__o22ai_4 _13796_ (.A1(_05250_),
    .A2(_05251_),
    .B1(_05283_),
    .B2(_05284_),
    .Y(_05287_));
 sky130_fd_sc_hd__o211a_2 _13797_ (.A1(_05132_),
    .A2(_05134_),
    .B1(_05286_),
    .C1(_05287_),
    .X(_05288_));
 sky130_fd_sc_hd__a211oi_4 _13798_ (.A1(_05286_),
    .A2(_05287_),
    .B1(_05132_),
    .C1(_05134_),
    .Y(_05289_));
 sky130_fd_sc_hd__nor4_1 _13799_ (.A(_05229_),
    .B(_05231_),
    .C(_05288_),
    .D(_05289_),
    .Y(_05290_));
 sky130_fd_sc_hd__or4_2 _13800_ (.A(_05229_),
    .B(_05231_),
    .C(_05288_),
    .D(_05289_),
    .X(_05291_));
 sky130_fd_sc_hd__o22ai_4 _13801_ (.A1(_05229_),
    .A2(_05231_),
    .B1(_05288_),
    .B2(_05289_),
    .Y(_05292_));
 sky130_fd_sc_hd__o211ai_4 _13802_ (.A1(_05137_),
    .A2(_05139_),
    .B1(_05291_),
    .C1(_05292_),
    .Y(_05293_));
 sky130_fd_sc_hd__a211o_1 _13803_ (.A1(_05291_),
    .A2(_05292_),
    .B1(_05137_),
    .C1(_05139_),
    .X(_05294_));
 sky130_fd_sc_hd__or4bb_4 _13804_ (.A(_05193_),
    .B(_05194_),
    .C_N(_05293_),
    .D_N(_05294_),
    .X(_05295_));
 sky130_fd_sc_hd__a2bb2o_1 _13805_ (.A1_N(_05193_),
    .A2_N(_05194_),
    .B1(_05293_),
    .B2(_05294_),
    .X(_05296_));
 sky130_fd_sc_hd__o211a_1 _13806_ (.A1(_05142_),
    .A2(_05144_),
    .B1(_05295_),
    .C1(_05296_),
    .X(_05297_));
 sky130_fd_sc_hd__a211oi_2 _13807_ (.A1(_05295_),
    .A2(_05296_),
    .B1(_05142_),
    .C1(_05144_),
    .Y(_05298_));
 sky130_fd_sc_hd__a211o_1 _13808_ (.A1(_05040_),
    .A2(_05043_),
    .B1(_05297_),
    .C1(_05298_),
    .X(_05299_));
 sky130_fd_sc_hd__o211ai_4 _13809_ (.A1(_05297_),
    .A2(_05298_),
    .B1(_05040_),
    .C1(_05043_),
    .Y(_05300_));
 sky130_fd_sc_hd__o211ai_4 _13810_ (.A1(_05146_),
    .A2(_05148_),
    .B1(_05299_),
    .C1(_05300_),
    .Y(_05301_));
 sky130_fd_sc_hd__a211o_1 _13811_ (.A1(_05299_),
    .A2(_05300_),
    .B1(_05146_),
    .C1(_05148_),
    .X(_05302_));
 sky130_fd_sc_hd__nand2_2 _13812_ (.A(_05301_),
    .B(_05302_),
    .Y(_05303_));
 sky130_fd_sc_hd__xnor2_2 _13813_ (.A(_05150_),
    .B(_05303_),
    .Y(_05304_));
 sky130_fd_sc_hd__xor2_4 _13814_ (.A(_05159_),
    .B(_05304_),
    .X(_05305_));
 sky130_fd_sc_hd__nor2_1 _13815_ (.A(_03057_),
    .B(_05305_),
    .Y(_05306_));
 sky130_fd_sc_hd__a221o_1 _13816_ (.A1(net600),
    .A2(\temp[12] ),
    .B1(_02626_),
    .B2(net5),
    .C1(_05306_),
    .X(_05307_));
 sky130_fd_sc_hd__mux2_1 _13817_ (.A0(net675),
    .A1(_05307_),
    .S(net1),
    .X(_00279_));
 sky130_fd_sc_hd__and2b_1 _13818_ (.A_N(_05297_),
    .B(_05299_),
    .X(_05308_));
 sky130_fd_sc_hd__nor2_1 _13819_ (.A(_05191_),
    .B(_05193_),
    .Y(_05309_));
 sky130_fd_sc_hd__a22o_1 _13820_ (.A1(net569),
    .A2(net336),
    .B1(net333),
    .B2(net574),
    .X(_05310_));
 sky130_fd_sc_hd__inv_2 _13821_ (.A(_05310_),
    .Y(_05311_));
 sky130_fd_sc_hd__and4_1 _13822_ (.A(net569),
    .B(net573),
    .C(net336),
    .D(net333),
    .X(_05312_));
 sky130_fd_sc_hd__o2bb2a_1 _13823_ (.A1_N(net578),
    .A2_N(net330),
    .B1(_05311_),
    .B2(_05312_),
    .X(_05313_));
 sky130_fd_sc_hd__and4b_1 _13824_ (.A_N(_05312_),
    .B(net330),
    .C(net578),
    .D(_05310_),
    .X(_05314_));
 sky130_fd_sc_hd__or2_1 _13825_ (.A(_05313_),
    .B(_05314_),
    .X(_05315_));
 sky130_fd_sc_hd__a32o_1 _13826_ (.A1(net584),
    .A2(net330),
    .A3(_05161_),
    .B1(_05162_),
    .B2(net336),
    .X(_05316_));
 sky130_fd_sc_hd__or3b_2 _13827_ (.A(_05313_),
    .B(_05314_),
    .C_N(_05316_),
    .X(_05317_));
 sky130_fd_sc_hd__xor2_1 _13828_ (.A(_05315_),
    .B(_05316_),
    .X(_05318_));
 sky130_fd_sc_hd__nand2_1 _13829_ (.A(net584),
    .B(net328),
    .Y(_05319_));
 sky130_fd_sc_hd__or2_1 _13830_ (.A(_05318_),
    .B(_05319_),
    .X(_05320_));
 sky130_fd_sc_hd__xor2_1 _13831_ (.A(_05318_),
    .B(_05319_),
    .X(_05321_));
 sky130_fd_sc_hd__and2_1 _13832_ (.A(_05166_),
    .B(_05321_),
    .X(_05322_));
 sky130_fd_sc_hd__nor2_1 _13833_ (.A(_05166_),
    .B(_05321_),
    .Y(_05323_));
 sky130_fd_sc_hd__or2_1 _13834_ (.A(_05322_),
    .B(_05323_),
    .X(_05324_));
 sky130_fd_sc_hd__or2_1 _13835_ (.A(_05171_),
    .B(_05173_),
    .X(_05325_));
 sky130_fd_sc_hd__a22o_1 _13836_ (.A1(net555),
    .A2(net345),
    .B1(net340),
    .B2(net559),
    .X(_05326_));
 sky130_fd_sc_hd__nand4_1 _13837_ (.A(net555),
    .B(net559),
    .C(net345),
    .D(net340),
    .Y(_05327_));
 sky130_fd_sc_hd__a22oi_2 _13838_ (.A1(net562),
    .A2(net337),
    .B1(_05326_),
    .B2(_05327_),
    .Y(_05328_));
 sky130_fd_sc_hd__and4_1 _13839_ (.A(net562),
    .B(net337),
    .C(_05326_),
    .D(_05327_),
    .X(_05329_));
 sky130_fd_sc_hd__a211o_1 _13840_ (.A1(_05196_),
    .A2(_05198_),
    .B1(_05328_),
    .C1(_05329_),
    .X(_05330_));
 sky130_fd_sc_hd__o211ai_1 _13841_ (.A1(_05328_),
    .A2(_05329_),
    .B1(_05196_),
    .C1(_05198_),
    .Y(_05331_));
 sky130_fd_sc_hd__and2_1 _13842_ (.A(_05330_),
    .B(_05331_),
    .X(_05332_));
 sky130_fd_sc_hd__nand2_1 _13843_ (.A(_05325_),
    .B(_05332_),
    .Y(_05333_));
 sky130_fd_sc_hd__xnor2_2 _13844_ (.A(_05325_),
    .B(_05332_),
    .Y(_05334_));
 sky130_fd_sc_hd__a21oi_4 _13845_ (.A1(_05206_),
    .A2(_05208_),
    .B1(_05334_),
    .Y(_05335_));
 sky130_fd_sc_hd__and3_1 _13846_ (.A(_05206_),
    .B(_05208_),
    .C(_05334_),
    .X(_05336_));
 sky130_fd_sc_hd__a211oi_4 _13847_ (.A1(_05174_),
    .A2(_05177_),
    .B1(_05335_),
    .C1(_05336_),
    .Y(_05337_));
 sky130_fd_sc_hd__o211a_1 _13848_ (.A1(_05335_),
    .A2(_05336_),
    .B1(_05174_),
    .C1(_05177_),
    .X(_05338_));
 sky130_fd_sc_hd__a211oi_2 _13849_ (.A1(_05180_),
    .A2(_05183_),
    .B1(_05337_),
    .C1(_05338_),
    .Y(_05339_));
 sky130_fd_sc_hd__o211a_1 _13850_ (.A1(_05337_),
    .A2(_05338_),
    .B1(_05180_),
    .C1(_05183_),
    .X(_05340_));
 sky130_fd_sc_hd__nor3_2 _13851_ (.A(_05324_),
    .B(_05339_),
    .C(_05340_),
    .Y(_05341_));
 sky130_fd_sc_hd__o21a_1 _13852_ (.A1(_05339_),
    .A2(_05340_),
    .B1(_05324_),
    .X(_05342_));
 sky130_fd_sc_hd__a211oi_4 _13853_ (.A1(_05227_),
    .A2(_05230_),
    .B1(_05341_),
    .C1(_05342_),
    .Y(_05343_));
 sky130_fd_sc_hd__o211a_1 _13854_ (.A1(_05341_),
    .A2(_05342_),
    .B1(_05227_),
    .C1(_05230_),
    .X(_05344_));
 sky130_fd_sc_hd__a211oi_4 _13855_ (.A1(_05186_),
    .A2(_05189_),
    .B1(_05343_),
    .C1(_05344_),
    .Y(_05345_));
 sky130_fd_sc_hd__o211a_1 _13856_ (.A1(_05343_),
    .A2(_05344_),
    .B1(_05186_),
    .C1(_05189_),
    .X(_05346_));
 sky130_fd_sc_hd__a22oi_2 _13857_ (.A1(net542),
    .A2(net356),
    .B1(net354),
    .B2(net546),
    .Y(_05347_));
 sky130_fd_sc_hd__and4_1 _13858_ (.A(net542),
    .B(net546),
    .C(net356),
    .D(net354),
    .X(_05348_));
 sky130_fd_sc_hd__nor2_1 _13859_ (.A(_05347_),
    .B(_05348_),
    .Y(_05349_));
 sky130_fd_sc_hd__nand2_1 _13860_ (.A(net550),
    .B(net348),
    .Y(_05350_));
 sky130_fd_sc_hd__xnor2_2 _13861_ (.A(_05349_),
    .B(_05350_),
    .Y(_05351_));
 sky130_fd_sc_hd__a22o_1 _13862_ (.A1(net527),
    .A2(net632),
    .B1(net367),
    .B2(net532),
    .X(_05352_));
 sky130_fd_sc_hd__and4_1 _13863_ (.A(net527),
    .B(net532),
    .C(net632),
    .D(net367),
    .X(_05353_));
 sky130_fd_sc_hd__nand4_1 _13864_ (.A(\mul0.a[12] ),
    .B(net532),
    .C(net632),
    .D(net367),
    .Y(_05354_));
 sky130_fd_sc_hd__a22o_1 _13865_ (.A1(net537),
    .A2(net363),
    .B1(_05352_),
    .B2(_05354_),
    .X(_05355_));
 sky130_fd_sc_hd__and4_1 _13866_ (.A(net537),
    .B(net363),
    .C(_05352_),
    .D(_05354_),
    .X(_05356_));
 sky130_fd_sc_hd__nand4_1 _13867_ (.A(net537),
    .B(net363),
    .C(_05352_),
    .D(_05354_),
    .Y(_05357_));
 sky130_fd_sc_hd__o211a_1 _13868_ (.A1(_05201_),
    .A2(_05203_),
    .B1(_05355_),
    .C1(_05357_),
    .X(_05358_));
 sky130_fd_sc_hd__a211o_1 _13869_ (.A1(_05355_),
    .A2(_05357_),
    .B1(_05201_),
    .C1(_05203_),
    .X(_05359_));
 sky130_fd_sc_hd__nand2b_1 _13870_ (.A_N(_05358_),
    .B(_05359_),
    .Y(_05360_));
 sky130_fd_sc_hd__xnor2_2 _13871_ (.A(_05351_),
    .B(_05360_),
    .Y(_05361_));
 sky130_fd_sc_hd__a41o_1 _13872_ (.A1(net517),
    .A2(net521),
    .A3(net383),
    .A4(net377),
    .B1(_05215_),
    .X(_05362_));
 sky130_fd_sc_hd__a31o_1 _13873_ (.A1(net512),
    .A2(net387),
    .A3(_05232_),
    .B1(_05233_),
    .X(_05363_));
 sky130_fd_sc_hd__a22o_1 _13874_ (.A1(\mul0.a[15] ),
    .A2(net383),
    .B1(net377),
    .B2(net517),
    .X(_05364_));
 sky130_fd_sc_hd__nand4_1 _13875_ (.A(\mul0.a[15] ),
    .B(net517),
    .C(net383),
    .D(net377),
    .Y(_05365_));
 sky130_fd_sc_hd__a22o_1 _13876_ (.A1(net524),
    .A2(net374),
    .B1(_05364_),
    .B2(_05365_),
    .X(_05366_));
 sky130_fd_sc_hd__nand4_1 _13877_ (.A(net524),
    .B(net374),
    .C(_05364_),
    .D(_05365_),
    .Y(_05367_));
 sky130_fd_sc_hd__and3_1 _13878_ (.A(_05363_),
    .B(_05366_),
    .C(_05367_),
    .X(_05368_));
 sky130_fd_sc_hd__a21o_1 _13879_ (.A1(_05366_),
    .A2(_05367_),
    .B1(_05363_),
    .X(_05369_));
 sky130_fd_sc_hd__and2b_1 _13880_ (.A_N(_05368_),
    .B(_05369_),
    .X(_05370_));
 sky130_fd_sc_hd__xnor2_1 _13881_ (.A(_05362_),
    .B(_05370_),
    .Y(_05371_));
 sky130_fd_sc_hd__a21o_2 _13882_ (.A1(_05216_),
    .A2(_05219_),
    .B1(_05371_),
    .X(_05372_));
 sky130_fd_sc_hd__nand3_2 _13883_ (.A(_05216_),
    .B(_05219_),
    .C(_05371_),
    .Y(_05373_));
 sky130_fd_sc_hd__nand3_4 _13884_ (.A(_05361_),
    .B(_05372_),
    .C(_05373_),
    .Y(_05374_));
 sky130_fd_sc_hd__a21o_1 _13885_ (.A1(_05372_),
    .A2(_05373_),
    .B1(_05361_),
    .X(_05375_));
 sky130_fd_sc_hd__o211ai_4 _13886_ (.A1(_05248_),
    .A2(_05250_),
    .B1(_05374_),
    .C1(_05375_),
    .Y(_05376_));
 sky130_fd_sc_hd__a211o_1 _13887_ (.A1(_05374_),
    .A2(_05375_),
    .B1(_05248_),
    .C1(_05250_),
    .X(_05377_));
 sky130_fd_sc_hd__o211a_1 _13888_ (.A1(_05221_),
    .A2(_05224_),
    .B1(_05376_),
    .C1(_05377_),
    .X(_05378_));
 sky130_fd_sc_hd__o211ai_2 _13889_ (.A1(_05221_),
    .A2(_05224_),
    .B1(_05376_),
    .C1(_05377_),
    .Y(_05379_));
 sky130_fd_sc_hd__a211oi_2 _13890_ (.A1(_05376_),
    .A2(_05377_),
    .B1(_05221_),
    .C1(_05224_),
    .Y(_05380_));
 sky130_fd_sc_hd__a21o_1 _13891_ (.A1(_05252_),
    .A2(_05259_),
    .B1(_05258_),
    .X(_05381_));
 sky130_fd_sc_hd__a22o_1 _13892_ (.A1(net504),
    .A2(net392),
    .B1(net499),
    .B2(net397),
    .X(_05382_));
 sky130_fd_sc_hd__and3_1 _13893_ (.A(net504),
    .B(net397),
    .C(net392),
    .X(_05383_));
 sky130_fd_sc_hd__a21bo_1 _13894_ (.A1(net499),
    .A2(_05383_),
    .B1_N(_05382_),
    .X(_05384_));
 sky130_fd_sc_hd__nand2_1 _13895_ (.A(net508),
    .B(net387),
    .Y(_05385_));
 sky130_fd_sc_hd__xor2_1 _13896_ (.A(_05384_),
    .B(_05385_),
    .X(_05386_));
 sky130_fd_sc_hd__a22o_1 _13897_ (.A1(net407),
    .A2(net491),
    .B1(net487),
    .B2(net411),
    .X(_05387_));
 sky130_fd_sc_hd__nand4_1 _13898_ (.A(net411),
    .B(net407),
    .C(net491),
    .D(net487),
    .Y(_05388_));
 sky130_fd_sc_hd__and2_1 _13899_ (.A(net403),
    .B(net495),
    .X(_05389_));
 sky130_fd_sc_hd__a21oi_1 _13900_ (.A1(_05387_),
    .A2(_05388_),
    .B1(_05389_),
    .Y(_05390_));
 sky130_fd_sc_hd__and3_1 _13901_ (.A(_05387_),
    .B(_05388_),
    .C(_05389_),
    .X(_05391_));
 sky130_fd_sc_hd__a211o_1 _13902_ (.A1(_05239_),
    .A2(_05241_),
    .B1(_05390_),
    .C1(_05391_),
    .X(_05392_));
 sky130_fd_sc_hd__o211ai_2 _13903_ (.A1(_05390_),
    .A2(_05391_),
    .B1(_05239_),
    .C1(_05241_),
    .Y(_05393_));
 sky130_fd_sc_hd__nand3_1 _13904_ (.A(_05386_),
    .B(_05392_),
    .C(_05393_),
    .Y(_05394_));
 sky130_fd_sc_hd__a21o_1 _13905_ (.A1(_05392_),
    .A2(_05393_),
    .B1(_05386_),
    .X(_05395_));
 sky130_fd_sc_hd__and3_2 _13906_ (.A(_05381_),
    .B(_05394_),
    .C(_05395_),
    .X(_05396_));
 sky130_fd_sc_hd__a21oi_1 _13907_ (.A1(_05394_),
    .A2(_05395_),
    .B1(_05381_),
    .Y(_05397_));
 sky130_fd_sc_hd__a211oi_2 _13908_ (.A1(_05244_),
    .A2(_05246_),
    .B1(_05396_),
    .C1(_05397_),
    .Y(_05398_));
 sky130_fd_sc_hd__o211a_1 _13909_ (.A1(_05396_),
    .A2(_05397_),
    .B1(_05244_),
    .C1(_05246_),
    .X(_05399_));
 sky130_fd_sc_hd__nand2_1 _13910_ (.A(_05255_),
    .B(_05257_),
    .Y(_05400_));
 sky130_fd_sc_hd__a32o_1 _13911_ (.A1(net428),
    .A2(net474),
    .A3(_05263_),
    .B1(_05264_),
    .B2(net466),
    .X(_05401_));
 sky130_fd_sc_hd__a22o_1 _13912_ (.A1(net419),
    .A2(net478),
    .B1(net474),
    .B2(net423),
    .X(_05402_));
 sky130_fd_sc_hd__nand4_1 _13913_ (.A(net423),
    .B(net419),
    .C(net478),
    .D(net474),
    .Y(_05403_));
 sky130_fd_sc_hd__a22o_1 _13914_ (.A1(net415),
    .A2(net482),
    .B1(_05402_),
    .B2(_05403_),
    .X(_05404_));
 sky130_fd_sc_hd__nand4_1 _13915_ (.A(net415),
    .B(net482),
    .C(_05402_),
    .D(_05403_),
    .Y(_05405_));
 sky130_fd_sc_hd__and3_1 _13916_ (.A(_05401_),
    .B(_05404_),
    .C(_05405_),
    .X(_05406_));
 sky130_fd_sc_hd__a21o_1 _13917_ (.A1(_05404_),
    .A2(_05405_),
    .B1(_05401_),
    .X(_05407_));
 sky130_fd_sc_hd__and2b_1 _13918_ (.A_N(_05406_),
    .B(_05407_),
    .X(_05408_));
 sky130_fd_sc_hd__xor2_1 _13919_ (.A(_05400_),
    .B(_05408_),
    .X(_05409_));
 sky130_fd_sc_hd__a22oi_1 _13920_ (.A1(net433),
    .A2(net466),
    .B1(net463),
    .B2(net438),
    .Y(_05410_));
 sky130_fd_sc_hd__and4_1 _13921_ (.A(net438),
    .B(net433),
    .C(net466),
    .D(net463),
    .X(_05411_));
 sky130_fd_sc_hd__and4bb_1 _13922_ (.A_N(_05410_),
    .B_N(_05411_),
    .C(net428),
    .D(net470),
    .X(_05412_));
 sky130_fd_sc_hd__o2bb2a_1 _13923_ (.A1_N(net428),
    .A2_N(net470),
    .B1(_05410_),
    .B2(_05411_),
    .X(_05413_));
 sky130_fd_sc_hd__nor2_1 _13924_ (.A(_05412_),
    .B(_05413_),
    .Y(_05414_));
 sky130_fd_sc_hd__and2_1 _13925_ (.A(net442),
    .B(net460),
    .X(_05415_));
 sky130_fd_sc_hd__a22o_1 _13926_ (.A1(net447),
    .A2(net459),
    .B1(net457),
    .B2(net452),
    .X(_05416_));
 sky130_fd_sc_hd__nand4_2 _13927_ (.A(net452),
    .B(\mul0.b[1] ),
    .C(net459),
    .D(net457),
    .Y(_05417_));
 sky130_fd_sc_hd__nand3_1 _13928_ (.A(_05415_),
    .B(_05416_),
    .C(_05417_),
    .Y(_05418_));
 sky130_fd_sc_hd__a21o_1 _13929_ (.A1(_05416_),
    .A2(_05417_),
    .B1(_05415_),
    .X(_05419_));
 sky130_fd_sc_hd__a21bo_1 _13930_ (.A1(_05267_),
    .A2(_05268_),
    .B1_N(_05269_),
    .X(_05420_));
 sky130_fd_sc_hd__nand3_1 _13931_ (.A(_05418_),
    .B(_05419_),
    .C(_05420_),
    .Y(_05421_));
 sky130_fd_sc_hd__a21o_1 _13932_ (.A1(_05418_),
    .A2(_05419_),
    .B1(_05420_),
    .X(_05422_));
 sky130_fd_sc_hd__nand3_2 _13933_ (.A(_05414_),
    .B(_05421_),
    .C(_05422_),
    .Y(_05423_));
 sky130_fd_sc_hd__a21o_1 _13934_ (.A1(_05421_),
    .A2(_05422_),
    .B1(_05414_),
    .X(_05424_));
 sky130_fd_sc_hd__a21bo_1 _13935_ (.A1(_05266_),
    .A2(_05274_),
    .B1_N(_05273_),
    .X(_05425_));
 sky130_fd_sc_hd__nand3_4 _13936_ (.A(_05423_),
    .B(_05424_),
    .C(_05425_),
    .Y(_05426_));
 sky130_fd_sc_hd__a21o_1 _13937_ (.A1(_05423_),
    .A2(_05424_),
    .B1(_05425_),
    .X(_05427_));
 sky130_fd_sc_hd__and3_1 _13938_ (.A(_05409_),
    .B(_05426_),
    .C(_05427_),
    .X(_05428_));
 sky130_fd_sc_hd__nand3_2 _13939_ (.A(_05409_),
    .B(_05426_),
    .C(_05427_),
    .Y(_05429_));
 sky130_fd_sc_hd__a21oi_1 _13940_ (.A1(_05426_),
    .A2(_05427_),
    .B1(_05409_),
    .Y(_05430_));
 sky130_fd_sc_hd__a211o_1 _13941_ (.A1(_05278_),
    .A2(_05281_),
    .B1(_05428_),
    .C1(_05430_),
    .X(_05431_));
 sky130_fd_sc_hd__o211ai_1 _13942_ (.A1(_05428_),
    .A2(_05430_),
    .B1(_05278_),
    .C1(_05281_),
    .Y(_05432_));
 sky130_fd_sc_hd__or4bb_4 _13943_ (.A(_05398_),
    .B(_05399_),
    .C_N(_05431_),
    .D_N(_05432_),
    .X(_05433_));
 sky130_fd_sc_hd__a2bb2o_1 _13944_ (.A1_N(_05398_),
    .A2_N(_05399_),
    .B1(_05431_),
    .B2(_05432_),
    .X(_05434_));
 sky130_fd_sc_hd__o211a_2 _13945_ (.A1(_05283_),
    .A2(_05285_),
    .B1(_05433_),
    .C1(_05434_),
    .X(_05435_));
 sky130_fd_sc_hd__a211oi_4 _13946_ (.A1(_05433_),
    .A2(_05434_),
    .B1(_05283_),
    .C1(_05285_),
    .Y(_05436_));
 sky130_fd_sc_hd__nor4_2 _13947_ (.A(_05378_),
    .B(_05380_),
    .C(_05435_),
    .D(_05436_),
    .Y(_05437_));
 sky130_fd_sc_hd__or4_1 _13948_ (.A(_05378_),
    .B(_05380_),
    .C(_05435_),
    .D(_05436_),
    .X(_05438_));
 sky130_fd_sc_hd__o22ai_2 _13949_ (.A1(_05378_),
    .A2(_05380_),
    .B1(_05435_),
    .B2(_05436_),
    .Y(_05439_));
 sky130_fd_sc_hd__o211a_2 _13950_ (.A1(_05288_),
    .A2(_05290_),
    .B1(_05438_),
    .C1(_05439_),
    .X(_05440_));
 sky130_fd_sc_hd__a211oi_2 _13951_ (.A1(_05438_),
    .A2(_05439_),
    .B1(_05288_),
    .C1(_05290_),
    .Y(_05441_));
 sky130_fd_sc_hd__nor4_4 _13952_ (.A(_05345_),
    .B(_05346_),
    .C(_05440_),
    .D(_05441_),
    .Y(_05442_));
 sky130_fd_sc_hd__o22a_1 _13953_ (.A1(_05345_),
    .A2(_05346_),
    .B1(_05440_),
    .B2(_05441_),
    .X(_05443_));
 sky130_fd_sc_hd__a211oi_4 _13954_ (.A1(_05293_),
    .A2(_05295_),
    .B1(_05442_),
    .C1(_05443_),
    .Y(_05444_));
 sky130_fd_sc_hd__o211a_1 _13955_ (.A1(_05442_),
    .A2(_05443_),
    .B1(_05293_),
    .C1(_05295_),
    .X(_05445_));
 sky130_fd_sc_hd__nor3_2 _13956_ (.A(_05309_),
    .B(_05444_),
    .C(_05445_),
    .Y(_05446_));
 sky130_fd_sc_hd__o21a_1 _13957_ (.A1(_05444_),
    .A2(_05445_),
    .B1(_05309_),
    .X(_05447_));
 sky130_fd_sc_hd__nor2_2 _13958_ (.A(_05446_),
    .B(_05447_),
    .Y(_05448_));
 sky130_fd_sc_hd__and2b_1 _13959_ (.A_N(_05308_),
    .B(_05448_),
    .X(_05449_));
 sky130_fd_sc_hd__xnor2_2 _13960_ (.A(_05308_),
    .B(_05448_),
    .Y(_05450_));
 sky130_fd_sc_hd__and2b_1 _13961_ (.A_N(_05301_),
    .B(_05450_),
    .X(_05451_));
 sky130_fd_sc_hd__xor2_4 _13962_ (.A(_05301_),
    .B(_05450_),
    .X(_05452_));
 sky130_fd_sc_hd__a21oi_2 _13963_ (.A1(_05150_),
    .A2(_05153_),
    .B1(_05303_),
    .Y(_05453_));
 sky130_fd_sc_hd__and2b_1 _13964_ (.A_N(_05304_),
    .B(_05154_),
    .X(_05454_));
 sky130_fd_sc_hd__and2b_1 _13965_ (.A_N(_05014_),
    .B(_05454_),
    .X(_05455_));
 sky130_fd_sc_hd__nor2_2 _13966_ (.A(_05453_),
    .B(_05455_),
    .Y(_05456_));
 sky130_fd_sc_hd__xor2_4 _13967_ (.A(_05452_),
    .B(_05456_),
    .X(_05457_));
 sky130_fd_sc_hd__a22o_1 _13968_ (.A1(net600),
    .A2(net693),
    .B1(_02632_),
    .B2(net5),
    .X(_05458_));
 sky130_fd_sc_hd__a21o_1 _13969_ (.A1(_03058_),
    .A2(_05457_),
    .B1(_05458_),
    .X(_05459_));
 sky130_fd_sc_hd__mux2_1 _13970_ (.A0(net779),
    .A1(_05459_),
    .S(net2),
    .X(_00280_));
 sky130_fd_sc_hd__o21ba_2 _13971_ (.A1(_05452_),
    .A2(_05456_),
    .B1_N(_05451_),
    .X(_05460_));
 sky130_fd_sc_hd__nor2_1 _13972_ (.A(_05343_),
    .B(_05345_),
    .Y(_05461_));
 sky130_fd_sc_hd__or2_1 _13973_ (.A(_05339_),
    .B(_05341_),
    .X(_05462_));
 sky130_fd_sc_hd__a22oi_1 _13974_ (.A1(net559),
    .A2(net337),
    .B1(net336),
    .B2(net562),
    .Y(_05463_));
 sky130_fd_sc_hd__and4_1 _13975_ (.A(net559),
    .B(net562),
    .C(net337),
    .D(net336),
    .X(_05464_));
 sky130_fd_sc_hd__o2bb2a_1 _13976_ (.A1_N(net568),
    .A2_N(net333),
    .B1(_05463_),
    .B2(_05464_),
    .X(_05465_));
 sky130_fd_sc_hd__and4bb_1 _13977_ (.A_N(_05463_),
    .B_N(_05464_),
    .C(net569),
    .D(net333),
    .X(_05466_));
 sky130_fd_sc_hd__nor2_1 _13978_ (.A(_05465_),
    .B(_05466_),
    .Y(_05467_));
 sky130_fd_sc_hd__nor2_1 _13979_ (.A(_05312_),
    .B(_05314_),
    .Y(_05468_));
 sky130_fd_sc_hd__or3_1 _13980_ (.A(_05465_),
    .B(_05466_),
    .C(_05468_),
    .X(_05469_));
 sky130_fd_sc_hd__xnor2_1 _13981_ (.A(_05467_),
    .B(_05468_),
    .Y(_05470_));
 sky130_fd_sc_hd__a22oi_2 _13982_ (.A1(net574),
    .A2(net330),
    .B1(net328),
    .B2(net578),
    .Y(_05471_));
 sky130_fd_sc_hd__and4_2 _13983_ (.A(net574),
    .B(net578),
    .C(net330),
    .D(net328),
    .X(_05472_));
 sky130_fd_sc_hd__o22a_1 _13984_ (.A1(net584),
    .A2(net57),
    .B1(_05471_),
    .B2(_05472_),
    .X(_05473_));
 sky130_fd_sc_hd__nor4_2 _13985_ (.A(net584),
    .B(net57),
    .C(_05471_),
    .D(_05472_),
    .Y(_05474_));
 sky130_fd_sc_hd__or2_1 _13986_ (.A(_05473_),
    .B(_05474_),
    .X(_05475_));
 sky130_fd_sc_hd__inv_2 _13987_ (.A(_05475_),
    .Y(_05476_));
 sky130_fd_sc_hd__nand2_1 _13988_ (.A(_05470_),
    .B(_05476_),
    .Y(_05477_));
 sky130_fd_sc_hd__or2_1 _13989_ (.A(_05470_),
    .B(_05476_),
    .X(_05478_));
 sky130_fd_sc_hd__nand2_1 _13990_ (.A(_05477_),
    .B(_05478_),
    .Y(_05479_));
 sky130_fd_sc_hd__a21oi_4 _13991_ (.A1(_05317_),
    .A2(_05320_),
    .B1(_05479_),
    .Y(_05480_));
 sky130_fd_sc_hd__and3_1 _13992_ (.A(_05317_),
    .B(_05320_),
    .C(_05479_),
    .X(_05481_));
 sky130_fd_sc_hd__a21oi_1 _13993_ (.A1(_05351_),
    .A2(_05359_),
    .B1(_05358_),
    .Y(_05482_));
 sky130_fd_sc_hd__a41o_1 _13994_ (.A1(net555),
    .A2(net559),
    .A3(net345),
    .A4(net341),
    .B1(_05329_),
    .X(_05483_));
 sky130_fd_sc_hd__o21bai_2 _13995_ (.A1(_05347_),
    .A2(_05350_),
    .B1_N(_05348_),
    .Y(_05484_));
 sky130_fd_sc_hd__a22o_1 _13996_ (.A1(net546),
    .A2(net348),
    .B1(net344),
    .B2(net551),
    .X(_05485_));
 sky130_fd_sc_hd__nand4_2 _13997_ (.A(net547),
    .B(net551),
    .C(net348),
    .D(net344),
    .Y(_05486_));
 sky130_fd_sc_hd__a22o_1 _13998_ (.A1(net555),
    .A2(net340),
    .B1(_05485_),
    .B2(_05486_),
    .X(_05487_));
 sky130_fd_sc_hd__nand4_2 _13999_ (.A(net555),
    .B(net340),
    .C(_05485_),
    .D(_05486_),
    .Y(_05488_));
 sky130_fd_sc_hd__nand3_2 _14000_ (.A(_05484_),
    .B(_05487_),
    .C(_05488_),
    .Y(_05489_));
 sky130_fd_sc_hd__a21o_1 _14001_ (.A1(_05487_),
    .A2(_05488_),
    .B1(_05484_),
    .X(_05490_));
 sky130_fd_sc_hd__nand3_2 _14002_ (.A(_05483_),
    .B(_05489_),
    .C(_05490_),
    .Y(_05491_));
 sky130_fd_sc_hd__a21o_1 _14003_ (.A1(_05489_),
    .A2(_05490_),
    .B1(_05483_),
    .X(_05492_));
 sky130_fd_sc_hd__and3b_2 _14004_ (.A_N(_05482_),
    .B(_05491_),
    .C(_05492_),
    .X(_05493_));
 sky130_fd_sc_hd__a21boi_2 _14005_ (.A1(_05491_),
    .A2(_05492_),
    .B1_N(_05482_),
    .Y(_05494_));
 sky130_fd_sc_hd__a211oi_2 _14006_ (.A1(_05330_),
    .A2(_05333_),
    .B1(_05493_),
    .C1(_05494_),
    .Y(_05495_));
 sky130_fd_sc_hd__inv_2 _14007_ (.A(_05495_),
    .Y(_05496_));
 sky130_fd_sc_hd__o211ai_2 _14008_ (.A1(_05493_),
    .A2(_05494_),
    .B1(_05330_),
    .C1(_05333_),
    .Y(_05497_));
 sky130_fd_sc_hd__o211a_1 _14009_ (.A1(_05335_),
    .A2(_05337_),
    .B1(_05496_),
    .C1(_05497_),
    .X(_05498_));
 sky130_fd_sc_hd__a211oi_2 _14010_ (.A1(_05496_),
    .A2(_05497_),
    .B1(_05335_),
    .C1(_05337_),
    .Y(_05499_));
 sky130_fd_sc_hd__nor4_2 _14011_ (.A(_05480_),
    .B(_05481_),
    .C(_05498_),
    .D(_05499_),
    .Y(_05500_));
 sky130_fd_sc_hd__o22a_1 _14012_ (.A1(_05480_),
    .A2(_05481_),
    .B1(_05498_),
    .B2(_05499_),
    .X(_05501_));
 sky130_fd_sc_hd__a211o_1 _14013_ (.A1(_05376_),
    .A2(_05379_),
    .B1(_05500_),
    .C1(_05501_),
    .X(_05502_));
 sky130_fd_sc_hd__o211ai_2 _14014_ (.A1(_05500_),
    .A2(_05501_),
    .B1(_05376_),
    .C1(_05379_),
    .Y(_05503_));
 sky130_fd_sc_hd__and3_1 _14015_ (.A(_05462_),
    .B(_05502_),
    .C(_05503_),
    .X(_05504_));
 sky130_fd_sc_hd__a21oi_1 _14016_ (.A1(_05502_),
    .A2(_05503_),
    .B1(_05462_),
    .Y(_05505_));
 sky130_fd_sc_hd__a22o_1 _14017_ (.A1(net533),
    .A2(net364),
    .B1(net356),
    .B2(net538),
    .X(_05506_));
 sky130_fd_sc_hd__nand4_4 _14018_ (.A(net533),
    .B(net538),
    .C(net364),
    .D(net360),
    .Y(_05507_));
 sky130_fd_sc_hd__a22o_1 _14019_ (.A1(net543),
    .A2(net354),
    .B1(_05506_),
    .B2(_05507_),
    .X(_05508_));
 sky130_fd_sc_hd__nand4_2 _14020_ (.A(net543),
    .B(net352),
    .C(_05506_),
    .D(_05507_),
    .Y(_05509_));
 sky130_fd_sc_hd__and2_1 _14021_ (.A(_05508_),
    .B(_05509_),
    .X(_05510_));
 sky130_fd_sc_hd__a22o_1 _14022_ (.A1(net519),
    .A2(net372),
    .B1(net632),
    .B2(net521),
    .X(_05511_));
 sky130_fd_sc_hd__and4_1 _14023_ (.A(net519),
    .B(net523),
    .C(net372),
    .D(net633),
    .X(_05512_));
 sky130_fd_sc_hd__nand4_1 _14024_ (.A(net519),
    .B(net521),
    .C(net372),
    .D(net632),
    .Y(_05513_));
 sky130_fd_sc_hd__a22o_1 _14025_ (.A1(net529),
    .A2(net366),
    .B1(_05511_),
    .B2(_05513_),
    .X(_05514_));
 sky130_fd_sc_hd__and4_1 _14026_ (.A(net527),
    .B(net367),
    .C(_05511_),
    .D(_05513_),
    .X(_05515_));
 sky130_fd_sc_hd__nand4_1 _14027_ (.A(net527),
    .B(net366),
    .C(_05511_),
    .D(_05513_),
    .Y(_05516_));
 sky130_fd_sc_hd__o211a_1 _14028_ (.A1(_05353_),
    .A2(_05356_),
    .B1(_05514_),
    .C1(_05516_),
    .X(_05517_));
 sky130_fd_sc_hd__a211o_1 _14029_ (.A1(_05514_),
    .A2(_05516_),
    .B1(_05353_),
    .C1(_05356_),
    .X(_05518_));
 sky130_fd_sc_hd__and2b_1 _14030_ (.A_N(_05517_),
    .B(_05518_),
    .X(_05519_));
 sky130_fd_sc_hd__xnor2_2 _14031_ (.A(_05510_),
    .B(_05519_),
    .Y(_05520_));
 sky130_fd_sc_hd__nand2_1 _14032_ (.A(_05365_),
    .B(_05367_),
    .Y(_05521_));
 sky130_fd_sc_hd__a32o_1 _14033_ (.A1(\mul0.a[16] ),
    .A2(net387),
    .A3(_05382_),
    .B1(_05383_),
    .B2(net499),
    .X(_05522_));
 sky130_fd_sc_hd__a22o_1 _14034_ (.A1(net504),
    .A2(net387),
    .B1(net383),
    .B2(\mul0.a[16] ),
    .X(_05523_));
 sky130_fd_sc_hd__nand4_2 _14035_ (.A(net504),
    .B(\mul0.a[16] ),
    .C(net387),
    .D(net383),
    .Y(_05524_));
 sky130_fd_sc_hd__a22o_1 _14036_ (.A1(\mul0.a[15] ),
    .A2(net377),
    .B1(_05523_),
    .B2(_05524_),
    .X(_05525_));
 sky130_fd_sc_hd__nand4_2 _14037_ (.A(\mul0.a[15] ),
    .B(net377),
    .C(_05523_),
    .D(_05524_),
    .Y(_05526_));
 sky130_fd_sc_hd__nand3_1 _14038_ (.A(_05522_),
    .B(_05525_),
    .C(_05526_),
    .Y(_05527_));
 sky130_fd_sc_hd__a21o_1 _14039_ (.A1(_05525_),
    .A2(_05526_),
    .B1(_05522_),
    .X(_05528_));
 sky130_fd_sc_hd__nand3_1 _14040_ (.A(_05521_),
    .B(_05527_),
    .C(_05528_),
    .Y(_05529_));
 sky130_fd_sc_hd__a21o_1 _14041_ (.A1(_05527_),
    .A2(_05528_),
    .B1(_05521_),
    .X(_05530_));
 sky130_fd_sc_hd__a21o_1 _14042_ (.A1(_05362_),
    .A2(_05369_),
    .B1(_05368_),
    .X(_05531_));
 sky130_fd_sc_hd__and3_1 _14043_ (.A(_05529_),
    .B(_05530_),
    .C(_05531_),
    .X(_05532_));
 sky130_fd_sc_hd__a21oi_1 _14044_ (.A1(_05529_),
    .A2(_05530_),
    .B1(_05531_),
    .Y(_05533_));
 sky130_fd_sc_hd__or3_1 _14045_ (.A(_05520_),
    .B(_05532_),
    .C(_05533_),
    .X(_05534_));
 sky130_fd_sc_hd__o21ai_1 _14046_ (.A1(_05532_),
    .A2(_05533_),
    .B1(_05520_),
    .Y(_05535_));
 sky130_fd_sc_hd__o211a_1 _14047_ (.A1(_05396_),
    .A2(_05398_),
    .B1(_05534_),
    .C1(_05535_),
    .X(_05536_));
 sky130_fd_sc_hd__a211oi_2 _14048_ (.A1(_05534_),
    .A2(_05535_),
    .B1(_05396_),
    .C1(_05398_),
    .Y(_05537_));
 sky130_fd_sc_hd__a211oi_2 _14049_ (.A1(_05372_),
    .A2(_05374_),
    .B1(_05536_),
    .C1(_05537_),
    .Y(_05538_));
 sky130_fd_sc_hd__o211a_1 _14050_ (.A1(_05536_),
    .A2(_05537_),
    .B1(_05372_),
    .C1(_05374_),
    .X(_05539_));
 sky130_fd_sc_hd__nand2_1 _14051_ (.A(_05392_),
    .B(_05394_),
    .Y(_05540_));
 sky130_fd_sc_hd__a21o_1 _14052_ (.A1(_05400_),
    .A2(_05407_),
    .B1(_05406_),
    .X(_05541_));
 sky130_fd_sc_hd__nand2_1 _14053_ (.A(net392),
    .B(net499),
    .Y(_05542_));
 sky130_fd_sc_hd__a22o_1 _14054_ (.A1(net397),
    .A2(net495),
    .B1(net491),
    .B2(net403),
    .X(_05543_));
 sky130_fd_sc_hd__and3_1 _14055_ (.A(net403),
    .B(net397),
    .C(net491),
    .X(_05544_));
 sky130_fd_sc_hd__a21bo_1 _14056_ (.A1(net495),
    .A2(_05544_),
    .B1_N(_05543_),
    .X(_05545_));
 sky130_fd_sc_hd__xor2_1 _14057_ (.A(_05542_),
    .B(_05545_),
    .X(_05546_));
 sky130_fd_sc_hd__and2_1 _14058_ (.A(net406),
    .B(net487),
    .X(_05547_));
 sky130_fd_sc_hd__a22o_1 _14059_ (.A1(net410),
    .A2(net483),
    .B1(net481),
    .B2(net415),
    .X(_05548_));
 sky130_fd_sc_hd__nand4_1 _14060_ (.A(net415),
    .B(net410),
    .C(net483),
    .D(net481),
    .Y(_05549_));
 sky130_fd_sc_hd__a21o_1 _14061_ (.A1(_05548_),
    .A2(_05549_),
    .B1(_05547_),
    .X(_05550_));
 sky130_fd_sc_hd__nand3_1 _14062_ (.A(_05547_),
    .B(_05548_),
    .C(_05549_),
    .Y(_05551_));
 sky130_fd_sc_hd__a21bo_1 _14063_ (.A1(_05387_),
    .A2(_05389_),
    .B1_N(_05388_),
    .X(_05552_));
 sky130_fd_sc_hd__nand3_1 _14064_ (.A(_05550_),
    .B(_05551_),
    .C(_05552_),
    .Y(_05553_));
 sky130_fd_sc_hd__a21o_1 _14065_ (.A1(_05550_),
    .A2(_05551_),
    .B1(_05552_),
    .X(_05554_));
 sky130_fd_sc_hd__nand3_1 _14066_ (.A(_05546_),
    .B(_05553_),
    .C(_05554_),
    .Y(_05555_));
 sky130_fd_sc_hd__a21o_1 _14067_ (.A1(_05553_),
    .A2(_05554_),
    .B1(_05546_),
    .X(_05556_));
 sky130_fd_sc_hd__nand3_2 _14068_ (.A(_05541_),
    .B(_05555_),
    .C(_05556_),
    .Y(_05557_));
 sky130_fd_sc_hd__a21o_1 _14069_ (.A1(_05555_),
    .A2(_05556_),
    .B1(_05541_),
    .X(_05558_));
 sky130_fd_sc_hd__nand3_1 _14070_ (.A(_05540_),
    .B(_05557_),
    .C(_05558_),
    .Y(_05559_));
 sky130_fd_sc_hd__a21o_1 _14071_ (.A1(_05557_),
    .A2(_05558_),
    .B1(_05540_),
    .X(_05560_));
 sky130_fd_sc_hd__nand2_1 _14072_ (.A(_05559_),
    .B(_05560_),
    .Y(_05561_));
 sky130_fd_sc_hd__nand2_1 _14073_ (.A(_05403_),
    .B(_05405_),
    .Y(_05562_));
 sky130_fd_sc_hd__a22o_1 _14074_ (.A1(net423),
    .A2(net470),
    .B1(net467),
    .B2(net428),
    .X(_05563_));
 sky130_fd_sc_hd__nand4_2 _14075_ (.A(net428),
    .B(net423),
    .C(net470),
    .D(net467),
    .Y(_05564_));
 sky130_fd_sc_hd__a22o_1 _14076_ (.A1(net419),
    .A2(net474),
    .B1(_05563_),
    .B2(_05564_),
    .X(_05565_));
 sky130_fd_sc_hd__nand4_2 _14077_ (.A(net419),
    .B(net474),
    .C(_05563_),
    .D(_05564_),
    .Y(_05566_));
 sky130_fd_sc_hd__o211a_1 _14078_ (.A1(_05411_),
    .A2(_05412_),
    .B1(_05565_),
    .C1(_05566_),
    .X(_05567_));
 sky130_fd_sc_hd__a211o_1 _14079_ (.A1(_05565_),
    .A2(_05566_),
    .B1(_05411_),
    .C1(_05412_),
    .X(_05568_));
 sky130_fd_sc_hd__nand2b_1 _14080_ (.A_N(_05567_),
    .B(_05568_),
    .Y(_05569_));
 sky130_fd_sc_hd__xnor2_2 _14081_ (.A(_05562_),
    .B(_05569_),
    .Y(_05570_));
 sky130_fd_sc_hd__nand2_1 _14082_ (.A(net433),
    .B(net463),
    .Y(_05571_));
 sky130_fd_sc_hd__a22o_1 _14083_ (.A1(net438),
    .A2(net460),
    .B1(net459),
    .B2(net442),
    .X(_05572_));
 sky130_fd_sc_hd__and3_1 _14084_ (.A(net442),
    .B(net438),
    .C(net459),
    .X(_05573_));
 sky130_fd_sc_hd__a21bo_1 _14085_ (.A1(net460),
    .A2(_05573_),
    .B1_N(_05572_),
    .X(_05574_));
 sky130_fd_sc_hd__xor2_2 _14086_ (.A(_05571_),
    .B(_05574_),
    .X(_05575_));
 sky130_fd_sc_hd__nand2_1 _14087_ (.A(net447),
    .B(net457),
    .Y(_05576_));
 sky130_fd_sc_hd__a21oi_1 _14088_ (.A1(net451),
    .A2(\mul0.a[31] ),
    .B1(\mul0.b[31] ),
    .Y(_05577_));
 sky130_fd_sc_hd__and3_1 _14089_ (.A(net451),
    .B(\mul0.a[31] ),
    .C(\mul0.b[31] ),
    .X(_05578_));
 sky130_fd_sc_hd__or3_1 _14090_ (.A(_05576_),
    .B(_05577_),
    .C(_05578_),
    .X(_05579_));
 sky130_fd_sc_hd__o21ai_1 _14091_ (.A1(_05577_),
    .A2(_05578_),
    .B1(_05576_),
    .Y(_05580_));
 sky130_fd_sc_hd__a21bo_1 _14092_ (.A1(_05415_),
    .A2(_05416_),
    .B1_N(_05417_),
    .X(_05581_));
 sky130_fd_sc_hd__nand3_1 _14093_ (.A(_05579_),
    .B(_05580_),
    .C(_05581_),
    .Y(_05582_));
 sky130_fd_sc_hd__a21o_1 _14094_ (.A1(_05579_),
    .A2(_05580_),
    .B1(_05581_),
    .X(_05583_));
 sky130_fd_sc_hd__nand3_2 _14095_ (.A(_05575_),
    .B(_05582_),
    .C(_05583_),
    .Y(_05584_));
 sky130_fd_sc_hd__a21o_1 _14096_ (.A1(_05582_),
    .A2(_05583_),
    .B1(_05575_),
    .X(_05585_));
 sky130_fd_sc_hd__a21bo_1 _14097_ (.A1(_05414_),
    .A2(_05422_),
    .B1_N(_05421_),
    .X(_05586_));
 sky130_fd_sc_hd__nand3_4 _14098_ (.A(_05584_),
    .B(_05585_),
    .C(_05586_),
    .Y(_05587_));
 sky130_fd_sc_hd__a21o_1 _14099_ (.A1(_05584_),
    .A2(_05585_),
    .B1(_05586_),
    .X(_05588_));
 sky130_fd_sc_hd__and3_1 _14100_ (.A(_05570_),
    .B(_05587_),
    .C(_05588_),
    .X(_05589_));
 sky130_fd_sc_hd__nand3_2 _14101_ (.A(_05570_),
    .B(_05587_),
    .C(_05588_),
    .Y(_05590_));
 sky130_fd_sc_hd__a21oi_2 _14102_ (.A1(_05587_),
    .A2(_05588_),
    .B1(_05570_),
    .Y(_05591_));
 sky130_fd_sc_hd__a211oi_4 _14103_ (.A1(_05426_),
    .A2(_05429_),
    .B1(_05589_),
    .C1(_05591_),
    .Y(_05592_));
 sky130_fd_sc_hd__o211a_1 _14104_ (.A1(_05589_),
    .A2(_05591_),
    .B1(_05426_),
    .C1(_05429_),
    .X(_05593_));
 sky130_fd_sc_hd__nor3_2 _14105_ (.A(_05561_),
    .B(_05592_),
    .C(_05593_),
    .Y(_05594_));
 sky130_fd_sc_hd__o21a_1 _14106_ (.A1(_05592_),
    .A2(_05593_),
    .B1(_05561_),
    .X(_05595_));
 sky130_fd_sc_hd__a211o_2 _14107_ (.A1(_05431_),
    .A2(_05433_),
    .B1(_05594_),
    .C1(_05595_),
    .X(_05596_));
 sky130_fd_sc_hd__o211ai_1 _14108_ (.A1(_05594_),
    .A2(_05595_),
    .B1(_05431_),
    .C1(_05433_),
    .Y(_05597_));
 sky130_fd_sc_hd__or4bb_4 _14109_ (.A(_05538_),
    .B(_05539_),
    .C_N(_05596_),
    .D_N(_05597_),
    .X(_05598_));
 sky130_fd_sc_hd__a2bb2o_1 _14110_ (.A1_N(_05538_),
    .A2_N(_05539_),
    .B1(_05596_),
    .B2(_05597_),
    .X(_05599_));
 sky130_fd_sc_hd__o211ai_4 _14111_ (.A1(_05435_),
    .A2(_05437_),
    .B1(_05598_),
    .C1(_05599_),
    .Y(_05600_));
 sky130_fd_sc_hd__a211o_1 _14112_ (.A1(_05598_),
    .A2(_05599_),
    .B1(_05435_),
    .C1(_05437_),
    .X(_05601_));
 sky130_fd_sc_hd__or4bb_4 _14113_ (.A(_05504_),
    .B(_05505_),
    .C_N(_05600_),
    .D_N(_05601_),
    .X(_05602_));
 sky130_fd_sc_hd__a2bb2o_1 _14114_ (.A1_N(_05504_),
    .A2_N(_05505_),
    .B1(_05600_),
    .B2(_05601_),
    .X(_05603_));
 sky130_fd_sc_hd__o211a_1 _14115_ (.A1(_05440_),
    .A2(_05442_),
    .B1(_05602_),
    .C1(_05603_),
    .X(_05604_));
 sky130_fd_sc_hd__a211oi_1 _14116_ (.A1(_05602_),
    .A2(_05603_),
    .B1(_05440_),
    .C1(_05442_),
    .Y(_05605_));
 sky130_fd_sc_hd__or3_1 _14117_ (.A(_05461_),
    .B(_05604_),
    .C(_05605_),
    .X(_05606_));
 sky130_fd_sc_hd__o21ai_1 _14118_ (.A1(_05604_),
    .A2(_05605_),
    .B1(_05461_),
    .Y(_05607_));
 sky130_fd_sc_hd__o211a_1 _14119_ (.A1(_05444_),
    .A2(_05446_),
    .B1(_05606_),
    .C1(_05607_),
    .X(_05608_));
 sky130_fd_sc_hd__a211oi_2 _14120_ (.A1(_05606_),
    .A2(_05607_),
    .B1(_05444_),
    .C1(_05446_),
    .Y(_05609_));
 sky130_fd_sc_hd__or3b_2 _14121_ (.A(_05608_),
    .B(_05609_),
    .C_N(_05322_),
    .X(_05610_));
 sky130_fd_sc_hd__o21bai_2 _14122_ (.A1(_05608_),
    .A2(_05609_),
    .B1_N(_05322_),
    .Y(_05611_));
 sky130_fd_sc_hd__and3_1 _14123_ (.A(_05449_),
    .B(_05610_),
    .C(_05611_),
    .X(_05612_));
 sky130_fd_sc_hd__a21oi_1 _14124_ (.A1(_05610_),
    .A2(_05611_),
    .B1(_05449_),
    .Y(_05613_));
 sky130_fd_sc_hd__or2_2 _14125_ (.A(_05612_),
    .B(_05613_),
    .X(_05614_));
 sky130_fd_sc_hd__xor2_4 _14126_ (.A(_05460_),
    .B(_05614_),
    .X(_05615_));
 sky130_fd_sc_hd__a22o_1 _14127_ (.A1(net600),
    .A2(\temp[14] ),
    .B1(_02638_),
    .B2(net5),
    .X(_05616_));
 sky130_fd_sc_hd__a21o_1 _14128_ (.A1(_03058_),
    .A2(_05615_),
    .B1(_05616_),
    .X(_05617_));
 sky130_fd_sc_hd__mux2_1 _14129_ (.A0(net786),
    .A1(_05617_),
    .S(net4),
    .X(_00281_));
 sky130_fd_sc_hd__a21bo_1 _14130_ (.A1(_05462_),
    .A2(_05503_),
    .B1_N(_05502_),
    .X(_05618_));
 sky130_fd_sc_hd__nor2_1 _14131_ (.A(_05498_),
    .B(_05500_),
    .Y(_05619_));
 sky130_fd_sc_hd__nor2_2 _14132_ (.A(_05536_),
    .B(_05538_),
    .Y(_05620_));
 sky130_fd_sc_hd__and4b_2 _14133_ (.A_N(net579),
    .B(net328),
    .C(net326),
    .D(net574),
    .X(_05621_));
 sky130_fd_sc_hd__o2bb2a_1 _14134_ (.A1_N(net574),
    .A2_N(net328),
    .B1(net57),
    .B2(net578),
    .X(_05622_));
 sky130_fd_sc_hd__nor2_1 _14135_ (.A(_05621_),
    .B(_05622_),
    .Y(_05623_));
 sky130_fd_sc_hd__inv_2 _14136_ (.A(_05623_),
    .Y(_05624_));
 sky130_fd_sc_hd__a22o_1 _14137_ (.A1(net559),
    .A2(net335),
    .B1(net332),
    .B2(net563),
    .X(_05625_));
 sky130_fd_sc_hd__and3_1 _14138_ (.A(net559),
    .B(net563),
    .C(net335),
    .X(_05626_));
 sky130_fd_sc_hd__a21bo_1 _14139_ (.A1(net332),
    .A2(_05626_),
    .B1_N(_05625_),
    .X(_05627_));
 sky130_fd_sc_hd__nand2_1 _14140_ (.A(net569),
    .B(net330),
    .Y(_05628_));
 sky130_fd_sc_hd__xnor2_1 _14141_ (.A(_05627_),
    .B(_05628_),
    .Y(_05629_));
 sky130_fd_sc_hd__or2_1 _14142_ (.A(_05464_),
    .B(_05466_),
    .X(_05630_));
 sky130_fd_sc_hd__and2b_1 _14143_ (.A_N(_05629_),
    .B(_05630_),
    .X(_05631_));
 sky130_fd_sc_hd__xor2_1 _14144_ (.A(_05629_),
    .B(_05630_),
    .X(_05632_));
 sky130_fd_sc_hd__nor2_1 _14145_ (.A(_05624_),
    .B(_05632_),
    .Y(_05633_));
 sky130_fd_sc_hd__xnor2_1 _14146_ (.A(_05624_),
    .B(_05632_),
    .Y(_05634_));
 sky130_fd_sc_hd__a21oi_1 _14147_ (.A1(_05469_),
    .A2(_05477_),
    .B1(_05634_),
    .Y(_05635_));
 sky130_fd_sc_hd__a21o_1 _14148_ (.A1(_05469_),
    .A2(_05477_),
    .B1(_05634_),
    .X(_05636_));
 sky130_fd_sc_hd__nand3_1 _14149_ (.A(_05469_),
    .B(_05477_),
    .C(_05634_),
    .Y(_05637_));
 sky130_fd_sc_hd__o211a_1 _14150_ (.A1(_05472_),
    .A2(_05474_),
    .B1(_05636_),
    .C1(_05637_),
    .X(_05638_));
 sky130_fd_sc_hd__a211oi_2 _14151_ (.A1(_05636_),
    .A2(_05637_),
    .B1(_05472_),
    .C1(_05474_),
    .Y(_05639_));
 sky130_fd_sc_hd__a21o_1 _14152_ (.A1(_05510_),
    .A2(_05518_),
    .B1(_05517_),
    .X(_05640_));
 sky130_fd_sc_hd__nand2_1 _14153_ (.A(_05486_),
    .B(_05488_),
    .Y(_05641_));
 sky130_fd_sc_hd__a22o_1 _14154_ (.A1(net547),
    .A2(net344),
    .B1(net340),
    .B2(net551),
    .X(_05642_));
 sky130_fd_sc_hd__nand4_1 _14155_ (.A(net547),
    .B(net551),
    .C(net344),
    .D(net340),
    .Y(_05643_));
 sky130_fd_sc_hd__a22oi_2 _14156_ (.A1(net555),
    .A2(net337),
    .B1(_05642_),
    .B2(_05643_),
    .Y(_05644_));
 sky130_fd_sc_hd__and4_1 _14157_ (.A(net555),
    .B(net337),
    .C(_05642_),
    .D(_05643_),
    .X(_05645_));
 sky130_fd_sc_hd__a211o_1 _14158_ (.A1(_05507_),
    .A2(_05509_),
    .B1(_05644_),
    .C1(_05645_),
    .X(_05646_));
 sky130_fd_sc_hd__o211ai_2 _14159_ (.A1(_05644_),
    .A2(_05645_),
    .B1(_05507_),
    .C1(_05509_),
    .Y(_05647_));
 sky130_fd_sc_hd__nand3_2 _14160_ (.A(_05641_),
    .B(_05646_),
    .C(_05647_),
    .Y(_05648_));
 sky130_fd_sc_hd__a21o_1 _14161_ (.A1(_05646_),
    .A2(_05647_),
    .B1(_05641_),
    .X(_05649_));
 sky130_fd_sc_hd__and3_1 _14162_ (.A(_05640_),
    .B(_05648_),
    .C(_05649_),
    .X(_05650_));
 sky130_fd_sc_hd__a21oi_1 _14163_ (.A1(_05648_),
    .A2(_05649_),
    .B1(_05640_),
    .Y(_05651_));
 sky130_fd_sc_hd__a211o_1 _14164_ (.A1(_05489_),
    .A2(_05491_),
    .B1(_05650_),
    .C1(_05651_),
    .X(_05652_));
 sky130_fd_sc_hd__o211ai_2 _14165_ (.A1(_05650_),
    .A2(_05651_),
    .B1(_05489_),
    .C1(_05491_),
    .Y(_05653_));
 sky130_fd_sc_hd__o211a_1 _14166_ (.A1(_05493_),
    .A2(_05495_),
    .B1(_05652_),
    .C1(_05653_),
    .X(_05654_));
 sky130_fd_sc_hd__a211oi_2 _14167_ (.A1(_05652_),
    .A2(_05653_),
    .B1(_05493_),
    .C1(_05495_),
    .Y(_05655_));
 sky130_fd_sc_hd__nor4_2 _14168_ (.A(_05638_),
    .B(_05639_),
    .C(_05654_),
    .D(_05655_),
    .Y(_05656_));
 sky130_fd_sc_hd__o22a_1 _14169_ (.A1(_05638_),
    .A2(_05639_),
    .B1(_05654_),
    .B2(_05655_),
    .X(_05657_));
 sky130_fd_sc_hd__nor2_1 _14170_ (.A(_05656_),
    .B(_05657_),
    .Y(_05658_));
 sky130_fd_sc_hd__xnor2_2 _14171_ (.A(_05620_),
    .B(_05658_),
    .Y(_05659_));
 sky130_fd_sc_hd__nand2b_1 _14172_ (.A_N(_05619_),
    .B(_05659_),
    .Y(_05660_));
 sky130_fd_sc_hd__xnor2_2 _14173_ (.A(_05619_),
    .B(_05659_),
    .Y(_05661_));
 sky130_fd_sc_hd__and2b_1 _14174_ (.A_N(_05532_),
    .B(_05534_),
    .X(_05662_));
 sky130_fd_sc_hd__a22o_1 _14175_ (.A1(net533),
    .A2(net360),
    .B1(net352),
    .B2(net538),
    .X(_05663_));
 sky130_fd_sc_hd__and3_1 _14176_ (.A(net533),
    .B(net538),
    .C(net360),
    .X(_05664_));
 sky130_fd_sc_hd__a21bo_1 _14177_ (.A1(net352),
    .A2(_05664_),
    .B1_N(_05663_),
    .X(_05665_));
 sky130_fd_sc_hd__nand2_1 _14178_ (.A(net543),
    .B(net351),
    .Y(_05666_));
 sky130_fd_sc_hd__xor2_2 _14179_ (.A(_05665_),
    .B(_05666_),
    .X(_05667_));
 sky130_fd_sc_hd__a22o_1 _14180_ (.A1(net519),
    .A2(net633),
    .B1(net366),
    .B2(net523),
    .X(_05668_));
 sky130_fd_sc_hd__and4_1 _14181_ (.A(net519),
    .B(net523),
    .C(net632),
    .D(net366),
    .X(_05669_));
 sky130_fd_sc_hd__nand4_1 _14182_ (.A(net519),
    .B(net523),
    .C(net633),
    .D(net366),
    .Y(_05670_));
 sky130_fd_sc_hd__a22o_1 _14183_ (.A1(net529),
    .A2(net361),
    .B1(_05668_),
    .B2(_05670_),
    .X(_05671_));
 sky130_fd_sc_hd__and4_1 _14184_ (.A(net529),
    .B(net361),
    .C(_05668_),
    .D(_05670_),
    .X(_05672_));
 sky130_fd_sc_hd__nand4_1 _14185_ (.A(net529),
    .B(net361),
    .C(_05668_),
    .D(_05670_),
    .Y(_05673_));
 sky130_fd_sc_hd__o211a_1 _14186_ (.A1(_05512_),
    .A2(_05515_),
    .B1(_05671_),
    .C1(_05673_),
    .X(_05674_));
 sky130_fd_sc_hd__a211o_1 _14187_ (.A1(_05671_),
    .A2(_05673_),
    .B1(_05512_),
    .C1(_05515_),
    .X(_05675_));
 sky130_fd_sc_hd__nand2b_1 _14188_ (.A_N(_05674_),
    .B(_05675_),
    .Y(_05676_));
 sky130_fd_sc_hd__xnor2_2 _14189_ (.A(_05667_),
    .B(_05676_),
    .Y(_05677_));
 sky130_fd_sc_hd__nand2_1 _14190_ (.A(_05524_),
    .B(_05526_),
    .Y(_05678_));
 sky130_fd_sc_hd__a32o_1 _14191_ (.A1(net392),
    .A2(net499),
    .A3(_05543_),
    .B1(_05544_),
    .B2(net495),
    .X(_05679_));
 sky130_fd_sc_hd__a22o_1 _14192_ (.A1(\mul0.a[17] ),
    .A2(net383),
    .B1(net377),
    .B2(net508),
    .X(_05680_));
 sky130_fd_sc_hd__nand4_2 _14193_ (.A(net504),
    .B(net508),
    .C(net383),
    .D(net377),
    .Y(_05681_));
 sky130_fd_sc_hd__a22o_1 _14194_ (.A1(net512),
    .A2(net374),
    .B1(_05680_),
    .B2(_05681_),
    .X(_05682_));
 sky130_fd_sc_hd__nand4_2 _14195_ (.A(net512),
    .B(net374),
    .C(_05680_),
    .D(_05681_),
    .Y(_05683_));
 sky130_fd_sc_hd__nand3_1 _14196_ (.A(_05679_),
    .B(_05682_),
    .C(_05683_),
    .Y(_05684_));
 sky130_fd_sc_hd__a21o_1 _14197_ (.A1(_05682_),
    .A2(_05683_),
    .B1(_05679_),
    .X(_05685_));
 sky130_fd_sc_hd__nand3_1 _14198_ (.A(_05678_),
    .B(_05684_),
    .C(_05685_),
    .Y(_05686_));
 sky130_fd_sc_hd__a21o_1 _14199_ (.A1(_05684_),
    .A2(_05685_),
    .B1(_05678_),
    .X(_05687_));
 sky130_fd_sc_hd__a21bo_1 _14200_ (.A1(_05521_),
    .A2(_05528_),
    .B1_N(_05527_),
    .X(_05688_));
 sky130_fd_sc_hd__nand3_1 _14201_ (.A(_05686_),
    .B(_05687_),
    .C(_05688_),
    .Y(_05689_));
 sky130_fd_sc_hd__a21o_1 _14202_ (.A1(_05686_),
    .A2(_05687_),
    .B1(_05688_),
    .X(_05690_));
 sky130_fd_sc_hd__and3_1 _14203_ (.A(_05677_),
    .B(_05689_),
    .C(_05690_),
    .X(_05691_));
 sky130_fd_sc_hd__a21oi_1 _14204_ (.A1(_05689_),
    .A2(_05690_),
    .B1(_05677_),
    .Y(_05692_));
 sky130_fd_sc_hd__a211o_1 _14205_ (.A1(_05557_),
    .A2(_05559_),
    .B1(_05691_),
    .C1(_05692_),
    .X(_05693_));
 sky130_fd_sc_hd__o211ai_1 _14206_ (.A1(_05691_),
    .A2(_05692_),
    .B1(_05557_),
    .C1(_05559_),
    .Y(_05694_));
 sky130_fd_sc_hd__nand2_2 _14207_ (.A(_05693_),
    .B(_05694_),
    .Y(_05695_));
 sky130_fd_sc_hd__xor2_1 _14208_ (.A(_05662_),
    .B(_05695_),
    .X(_05696_));
 sky130_fd_sc_hd__nand2_1 _14209_ (.A(_05553_),
    .B(_05555_),
    .Y(_05697_));
 sky130_fd_sc_hd__a21o_1 _14210_ (.A1(_05562_),
    .A2(_05568_),
    .B1(_05567_),
    .X(_05698_));
 sky130_fd_sc_hd__a22o_1 _14211_ (.A1(net392),
    .A2(net495),
    .B1(net491),
    .B2(net397),
    .X(_05699_));
 sky130_fd_sc_hd__nand4_1 _14212_ (.A(net397),
    .B(net392),
    .C(net495),
    .D(net491),
    .Y(_05700_));
 sky130_fd_sc_hd__nand2_1 _14213_ (.A(_05699_),
    .B(_05700_),
    .Y(_05701_));
 sky130_fd_sc_hd__and2_1 _14214_ (.A(net387),
    .B(net499),
    .X(_05702_));
 sky130_fd_sc_hd__xnor2_1 _14215_ (.A(_05701_),
    .B(_05702_),
    .Y(_05703_));
 sky130_fd_sc_hd__a22o_1 _14216_ (.A1(net406),
    .A2(net483),
    .B1(net481),
    .B2(net410),
    .X(_05704_));
 sky130_fd_sc_hd__nand4_1 _14217_ (.A(net410),
    .B(net406),
    .C(net483),
    .D(net481),
    .Y(_05705_));
 sky130_fd_sc_hd__and2_1 _14218_ (.A(net402),
    .B(net487),
    .X(_05706_));
 sky130_fd_sc_hd__a21o_1 _14219_ (.A1(_05704_),
    .A2(_05705_),
    .B1(_05706_),
    .X(_05707_));
 sky130_fd_sc_hd__nand3_1 _14220_ (.A(_05704_),
    .B(_05705_),
    .C(_05706_),
    .Y(_05708_));
 sky130_fd_sc_hd__a21bo_1 _14221_ (.A1(_05547_),
    .A2(_05548_),
    .B1_N(_05549_),
    .X(_05709_));
 sky130_fd_sc_hd__nand3_2 _14222_ (.A(_05707_),
    .B(_05708_),
    .C(_05709_),
    .Y(_05710_));
 sky130_fd_sc_hd__a21o_1 _14223_ (.A1(_05707_),
    .A2(_05708_),
    .B1(_05709_),
    .X(_05711_));
 sky130_fd_sc_hd__nand3_2 _14224_ (.A(_05703_),
    .B(_05710_),
    .C(_05711_),
    .Y(_05712_));
 sky130_fd_sc_hd__a21o_1 _14225_ (.A1(_05710_),
    .A2(_05711_),
    .B1(_05703_),
    .X(_05713_));
 sky130_fd_sc_hd__nand3_2 _14226_ (.A(_05698_),
    .B(_05712_),
    .C(_05713_),
    .Y(_05714_));
 sky130_fd_sc_hd__a21o_1 _14227_ (.A1(_05712_),
    .A2(_05713_),
    .B1(_05698_),
    .X(_05715_));
 sky130_fd_sc_hd__nand3_1 _14228_ (.A(_05697_),
    .B(_05714_),
    .C(_05715_),
    .Y(_05716_));
 sky130_fd_sc_hd__a21o_1 _14229_ (.A1(_05714_),
    .A2(_05715_),
    .B1(_05697_),
    .X(_05717_));
 sky130_fd_sc_hd__and2_1 _14230_ (.A(_05716_),
    .B(_05717_),
    .X(_05718_));
 sky130_fd_sc_hd__nand2_1 _14231_ (.A(_05564_),
    .B(_05566_),
    .Y(_05719_));
 sky130_fd_sc_hd__a32o_1 _14232_ (.A1(net433),
    .A2(net463),
    .A3(_05572_),
    .B1(_05573_),
    .B2(net460),
    .X(_05720_));
 sky130_fd_sc_hd__a22o_1 _14233_ (.A1(net419),
    .A2(net473),
    .B1(net467),
    .B2(net423),
    .X(_05721_));
 sky130_fd_sc_hd__nand4_2 _14234_ (.A(net423),
    .B(net419),
    .C(net470),
    .D(net467),
    .Y(_05722_));
 sky130_fd_sc_hd__a22o_1 _14235_ (.A1(net415),
    .A2(net477),
    .B1(_05721_),
    .B2(_05722_),
    .X(_05723_));
 sky130_fd_sc_hd__nand4_2 _14236_ (.A(net415),
    .B(net477),
    .C(_05721_),
    .D(_05722_),
    .Y(_05724_));
 sky130_fd_sc_hd__and3_1 _14237_ (.A(_05720_),
    .B(_05723_),
    .C(_05724_),
    .X(_05725_));
 sky130_fd_sc_hd__a21o_1 _14238_ (.A1(_05723_),
    .A2(_05724_),
    .B1(_05720_),
    .X(_05726_));
 sky130_fd_sc_hd__and2b_1 _14239_ (.A_N(_05725_),
    .B(_05726_),
    .X(_05727_));
 sky130_fd_sc_hd__xor2_2 _14240_ (.A(_05719_),
    .B(_05727_),
    .X(_05728_));
 sky130_fd_sc_hd__a22o_1 _14241_ (.A1(net433),
    .A2(net460),
    .B1(net459),
    .B2(net438),
    .X(_05729_));
 sky130_fd_sc_hd__and3_1 _14242_ (.A(net438),
    .B(net433),
    .C(net459),
    .X(_05730_));
 sky130_fd_sc_hd__a21bo_1 _14243_ (.A1(net460),
    .A2(_05730_),
    .B1_N(_05729_),
    .X(_05731_));
 sky130_fd_sc_hd__nand2_1 _14244_ (.A(net428),
    .B(net463),
    .Y(_05732_));
 sky130_fd_sc_hd__xor2_1 _14245_ (.A(_05731_),
    .B(_05732_),
    .X(_05733_));
 sky130_fd_sc_hd__o21bai_1 _14246_ (.A1(_05576_),
    .A2(_05577_),
    .B1_N(_05578_),
    .Y(_05734_));
 sky130_fd_sc_hd__or2_1 _14247_ (.A(net452),
    .B(\mul0.b[1] ),
    .X(_05735_));
 sky130_fd_sc_hd__and3_1 _14248_ (.A(net452),
    .B(\mul0.b[1] ),
    .C(net453),
    .X(_05736_));
 sky130_fd_sc_hd__a21boi_2 _14249_ (.A1(net452),
    .A2(\mul0.b[1] ),
    .B1_N(\mul0.a[31] ),
    .Y(_05737_));
 sky130_fd_sc_hd__nand2_1 _14250_ (.A(net442),
    .B(net457),
    .Y(_05738_));
 sky130_fd_sc_hd__and3_4 _14251_ (.A(_05735_),
    .B(_05737_),
    .C(_05738_),
    .X(_05739_));
 sky130_fd_sc_hd__a21oi_1 _14252_ (.A1(_05735_),
    .A2(_05737_),
    .B1(_05738_),
    .Y(_05740_));
 sky130_fd_sc_hd__o21ai_1 _14253_ (.A1(_05739_),
    .A2(_05740_),
    .B1(_05734_),
    .Y(_05741_));
 sky130_fd_sc_hd__or3_1 _14254_ (.A(_05734_),
    .B(_05739_),
    .C(_05740_),
    .X(_05742_));
 sky130_fd_sc_hd__nand3_1 _14255_ (.A(_05733_),
    .B(_05741_),
    .C(_05742_),
    .Y(_05743_));
 sky130_fd_sc_hd__a21o_1 _14256_ (.A1(_05741_),
    .A2(_05742_),
    .B1(_05733_),
    .X(_05744_));
 sky130_fd_sc_hd__a21bo_1 _14257_ (.A1(_05575_),
    .A2(_05583_),
    .B1_N(_05582_),
    .X(_05745_));
 sky130_fd_sc_hd__nand3_1 _14258_ (.A(_05743_),
    .B(_05744_),
    .C(_05745_),
    .Y(_05746_));
 sky130_fd_sc_hd__a21o_1 _14259_ (.A1(_05743_),
    .A2(_05744_),
    .B1(_05745_),
    .X(_05747_));
 sky130_fd_sc_hd__and3_1 _14260_ (.A(_05728_),
    .B(_05746_),
    .C(_05747_),
    .X(_05748_));
 sky130_fd_sc_hd__a21oi_2 _14261_ (.A1(_05746_),
    .A2(_05747_),
    .B1(_05728_),
    .Y(_05749_));
 sky130_fd_sc_hd__a211o_1 _14262_ (.A1(_05587_),
    .A2(_05590_),
    .B1(_05748_),
    .C1(_05749_),
    .X(_05750_));
 sky130_fd_sc_hd__o211ai_4 _14263_ (.A1(_05748_),
    .A2(_05749_),
    .B1(_05587_),
    .C1(_05590_),
    .Y(_05751_));
 sky130_fd_sc_hd__nand3_2 _14264_ (.A(_05718_),
    .B(_05750_),
    .C(_05751_),
    .Y(_05752_));
 sky130_fd_sc_hd__a21o_1 _14265_ (.A1(_05750_),
    .A2(_05751_),
    .B1(_05718_),
    .X(_05753_));
 sky130_fd_sc_hd__o211ai_4 _14266_ (.A1(_05592_),
    .A2(_05594_),
    .B1(_05752_),
    .C1(_05753_),
    .Y(_05754_));
 sky130_fd_sc_hd__a211o_1 _14267_ (.A1(_05752_),
    .A2(_05753_),
    .B1(_05592_),
    .C1(_05594_),
    .X(_05755_));
 sky130_fd_sc_hd__and3_1 _14268_ (.A(_05696_),
    .B(_05754_),
    .C(_05755_),
    .X(_05756_));
 sky130_fd_sc_hd__a21oi_2 _14269_ (.A1(_05754_),
    .A2(_05755_),
    .B1(_05696_),
    .Y(_05757_));
 sky130_fd_sc_hd__a211oi_1 _14270_ (.A1(_05596_),
    .A2(_05598_),
    .B1(_05756_),
    .C1(_05757_),
    .Y(_05758_));
 sky130_fd_sc_hd__a211o_1 _14271_ (.A1(_05596_),
    .A2(_05598_),
    .B1(_05756_),
    .C1(_05757_),
    .X(_05759_));
 sky130_fd_sc_hd__o211ai_4 _14272_ (.A1(_05756_),
    .A2(_05757_),
    .B1(_05596_),
    .C1(_05598_),
    .Y(_05760_));
 sky130_fd_sc_hd__and3_1 _14273_ (.A(_05661_),
    .B(_05759_),
    .C(_05760_),
    .X(_05761_));
 sky130_fd_sc_hd__a21oi_2 _14274_ (.A1(_05759_),
    .A2(_05760_),
    .B1(_05661_),
    .Y(_05762_));
 sky130_fd_sc_hd__a211o_1 _14275_ (.A1(_05600_),
    .A2(_05602_),
    .B1(_05761_),
    .C1(_05762_),
    .X(_05763_));
 sky130_fd_sc_hd__o211ai_4 _14276_ (.A1(_05761_),
    .A2(_05762_),
    .B1(_05600_),
    .C1(_05602_),
    .Y(_05764_));
 sky130_fd_sc_hd__and3_1 _14277_ (.A(_05618_),
    .B(_05763_),
    .C(_05764_),
    .X(_05765_));
 sky130_fd_sc_hd__a21oi_1 _14278_ (.A1(_05763_),
    .A2(_05764_),
    .B1(_05618_),
    .Y(_05766_));
 sky130_fd_sc_hd__or2_2 _14279_ (.A(_05765_),
    .B(_05766_),
    .X(_05767_));
 sky130_fd_sc_hd__and2b_1 _14280_ (.A_N(_05604_),
    .B(_05606_),
    .X(_05768_));
 sky130_fd_sc_hd__nor2_2 _14281_ (.A(_05767_),
    .B(_05768_),
    .Y(_05769_));
 sky130_fd_sc_hd__xor2_2 _14282_ (.A(_05767_),
    .B(_05768_),
    .X(_05770_));
 sky130_fd_sc_hd__and2_1 _14283_ (.A(_05480_),
    .B(_05770_),
    .X(_05771_));
 sky130_fd_sc_hd__xnor2_2 _14284_ (.A(_05480_),
    .B(_05770_),
    .Y(_05772_));
 sky130_fd_sc_hd__and2b_1 _14285_ (.A_N(_05608_),
    .B(_05610_),
    .X(_05773_));
 sky130_fd_sc_hd__or2_2 _14286_ (.A(_05772_),
    .B(_05773_),
    .X(_05774_));
 sky130_fd_sc_hd__nand2_1 _14287_ (.A(_05772_),
    .B(_05773_),
    .Y(_05775_));
 sky130_fd_sc_hd__and2_2 _14288_ (.A(_05774_),
    .B(_05775_),
    .X(_05776_));
 sky130_fd_sc_hd__xnor2_2 _14289_ (.A(_05772_),
    .B(_05773_),
    .Y(_05777_));
 sky130_fd_sc_hd__or2_1 _14290_ (.A(_05449_),
    .B(_05451_),
    .X(_05778_));
 sky130_fd_sc_hd__nor3_1 _14291_ (.A(_05452_),
    .B(_05612_),
    .C(_05613_),
    .Y(_05779_));
 sky130_fd_sc_hd__a32oi_2 _14292_ (.A1(_05610_),
    .A2(_05611_),
    .A3(_05778_),
    .B1(_05779_),
    .B2(_05453_),
    .Y(_05780_));
 sky130_fd_sc_hd__nand3_1 _14293_ (.A(_05013_),
    .B(_05454_),
    .C(_05779_),
    .Y(_05781_));
 sky130_fd_sc_hd__nand4b_1 _14294_ (.A_N(_05010_),
    .B(_05454_),
    .C(_05779_),
    .D(_04456_),
    .Y(_05782_));
 sky130_fd_sc_hd__and3_2 _14295_ (.A(_05780_),
    .B(_05781_),
    .C(_05782_),
    .X(_05783_));
 sky130_fd_sc_hd__xnor2_4 _14296_ (.A(_05776_),
    .B(_05783_),
    .Y(_05784_));
 sky130_fd_sc_hd__a22o_1 _14297_ (.A1(net599),
    .A2(net764),
    .B1(_02644_),
    .B2(net6),
    .X(_05785_));
 sky130_fd_sc_hd__a21o_1 _14298_ (.A1(_03058_),
    .A2(_05784_),
    .B1(_05785_),
    .X(_05786_));
 sky130_fd_sc_hd__mux2_1 _14299_ (.A0(net803),
    .A1(_05786_),
    .S(net4),
    .X(_00282_));
 sky130_fd_sc_hd__o21ai_4 _14300_ (.A1(_05777_),
    .A2(_05783_),
    .B1(_05774_),
    .Y(_05787_));
 sky130_fd_sc_hd__or2_1 _14301_ (.A(_05635_),
    .B(_05638_),
    .X(_05788_));
 sky130_fd_sc_hd__o31ai_4 _14302_ (.A1(_05620_),
    .A2(_05656_),
    .A3(_05657_),
    .B1(_05660_),
    .Y(_05789_));
 sky130_fd_sc_hd__nor2_2 _14303_ (.A(_05654_),
    .B(_05656_),
    .Y(_05790_));
 sky130_fd_sc_hd__o21ai_4 _14304_ (.A1(_05662_),
    .A2(_05695_),
    .B1(_05693_),
    .Y(_05791_));
 sky130_fd_sc_hd__a22o_1 _14305_ (.A1(net555),
    .A2(net335),
    .B1(net332),
    .B2(net560),
    .X(_05792_));
 sky130_fd_sc_hd__and3_1 _14306_ (.A(net555),
    .B(net560),
    .C(net332),
    .X(_05793_));
 sky130_fd_sc_hd__a21bo_2 _14307_ (.A1(net335),
    .A2(_05793_),
    .B1_N(_05792_),
    .X(_05794_));
 sky130_fd_sc_hd__nand2_2 _14308_ (.A(net563),
    .B(net329),
    .Y(_05795_));
 sky130_fd_sc_hd__xnor2_4 _14309_ (.A(_05794_),
    .B(_05795_),
    .Y(_05796_));
 sky130_fd_sc_hd__o2bb2a_2 _14310_ (.A1_N(net332),
    .A2_N(_05626_),
    .B1(_05627_),
    .B2(_05628_),
    .X(_05797_));
 sky130_fd_sc_hd__xnor2_2 _14311_ (.A(_05796_),
    .B(_05797_),
    .Y(_05798_));
 sky130_fd_sc_hd__and4b_2 _14312_ (.A_N(net574),
    .B(net328),
    .C(net326),
    .D(net569),
    .X(_05799_));
 sky130_fd_sc_hd__inv_2 _14313_ (.A(_05799_),
    .Y(_05800_));
 sky130_fd_sc_hd__o2bb2a_1 _14314_ (.A1_N(net569),
    .A2_N(net328),
    .B1(net57),
    .B2(net574),
    .X(_05801_));
 sky130_fd_sc_hd__nor2_1 _14315_ (.A(_05799_),
    .B(_05801_),
    .Y(_05802_));
 sky130_fd_sc_hd__xnor2_1 _14316_ (.A(_05798_),
    .B(_05802_),
    .Y(_05803_));
 sky130_fd_sc_hd__nor3_1 _14317_ (.A(_05631_),
    .B(_05633_),
    .C(_05803_),
    .Y(_05804_));
 sky130_fd_sc_hd__o21a_1 _14318_ (.A1(_05631_),
    .A2(_05633_),
    .B1(_05803_),
    .X(_05805_));
 sky130_fd_sc_hd__or2_2 _14319_ (.A(_05804_),
    .B(_05805_),
    .X(_05806_));
 sky130_fd_sc_hd__inv_2 _14320_ (.A(_05806_),
    .Y(_05807_));
 sky130_fd_sc_hd__xor2_4 _14321_ (.A(_05621_),
    .B(_05806_),
    .X(_05808_));
 sky130_fd_sc_hd__a21oi_1 _14322_ (.A1(_05667_),
    .A2(_05675_),
    .B1(_05674_),
    .Y(_05809_));
 sky130_fd_sc_hd__a41o_1 _14323_ (.A1(net547),
    .A2(net551),
    .A3(net344),
    .A4(net340),
    .B1(_05645_),
    .X(_05810_));
 sky130_fd_sc_hd__a32o_1 _14324_ (.A1(net543),
    .A2(net349),
    .A3(_05663_),
    .B1(_05664_),
    .B2(net352),
    .X(_05811_));
 sky130_fd_sc_hd__a22o_1 _14325_ (.A1(net543),
    .A2(net345),
    .B1(net341),
    .B2(net547),
    .X(_05812_));
 sky130_fd_sc_hd__nand4_2 _14326_ (.A(net543),
    .B(net547),
    .C(net345),
    .D(net341),
    .Y(_05813_));
 sky130_fd_sc_hd__a22o_1 _14327_ (.A1(net551),
    .A2(net339),
    .B1(_05812_),
    .B2(_05813_),
    .X(_05814_));
 sky130_fd_sc_hd__nand4_2 _14328_ (.A(net551),
    .B(net339),
    .C(_05812_),
    .D(_05813_),
    .Y(_05815_));
 sky130_fd_sc_hd__nand3_2 _14329_ (.A(_05811_),
    .B(_05814_),
    .C(_05815_),
    .Y(_05816_));
 sky130_fd_sc_hd__a21o_1 _14330_ (.A1(_05814_),
    .A2(_05815_),
    .B1(_05811_),
    .X(_05817_));
 sky130_fd_sc_hd__nand3_2 _14331_ (.A(_05810_),
    .B(_05816_),
    .C(_05817_),
    .Y(_05818_));
 sky130_fd_sc_hd__a21o_1 _14332_ (.A1(_05816_),
    .A2(_05817_),
    .B1(_05810_),
    .X(_05819_));
 sky130_fd_sc_hd__and3b_1 _14333_ (.A_N(_05809_),
    .B(_05818_),
    .C(_05819_),
    .X(_05820_));
 sky130_fd_sc_hd__a21boi_1 _14334_ (.A1(_05818_),
    .A2(_05819_),
    .B1_N(_05809_),
    .Y(_05821_));
 sky130_fd_sc_hd__a211oi_1 _14335_ (.A1(_05646_),
    .A2(_05648_),
    .B1(_05820_),
    .C1(_05821_),
    .Y(_05822_));
 sky130_fd_sc_hd__o211ai_1 _14336_ (.A1(_05820_),
    .A2(_05821_),
    .B1(_05646_),
    .C1(_05648_),
    .Y(_05823_));
 sky130_fd_sc_hd__nand2b_2 _14337_ (.A_N(_05822_),
    .B(_05823_),
    .Y(_05824_));
 sky130_fd_sc_hd__and2b_2 _14338_ (.A_N(_05650_),
    .B(_05652_),
    .X(_05825_));
 sky130_fd_sc_hd__nor2_1 _14339_ (.A(_05824_),
    .B(_05825_),
    .Y(_05826_));
 sky130_fd_sc_hd__xnor2_4 _14340_ (.A(_05824_),
    .B(_05825_),
    .Y(_05827_));
 sky130_fd_sc_hd__xnor2_4 _14341_ (.A(_05808_),
    .B(_05827_),
    .Y(_05828_));
 sky130_fd_sc_hd__and2b_1 _14342_ (.A_N(_05828_),
    .B(_05791_),
    .X(_05829_));
 sky130_fd_sc_hd__xnor2_4 _14343_ (.A(_05791_),
    .B(_05828_),
    .Y(_05830_));
 sky130_fd_sc_hd__and2b_1 _14344_ (.A_N(_05790_),
    .B(_05830_),
    .X(_05831_));
 sky130_fd_sc_hd__xnor2_4 _14345_ (.A(_05790_),
    .B(_05830_),
    .Y(_05832_));
 sky130_fd_sc_hd__a31o_1 _14346_ (.A1(_05686_),
    .A2(_05687_),
    .A3(_05688_),
    .B1(_05691_),
    .X(_05833_));
 sky130_fd_sc_hd__a22o_1 _14347_ (.A1(net529),
    .A2(net360),
    .B1(net352),
    .B2(net533),
    .X(_05834_));
 sky130_fd_sc_hd__and3_1 _14348_ (.A(net529),
    .B(net533),
    .C(net352),
    .X(_05835_));
 sky130_fd_sc_hd__a21bo_1 _14349_ (.A1(net360),
    .A2(_05835_),
    .B1_N(_05834_),
    .X(_05836_));
 sky130_fd_sc_hd__nand2_1 _14350_ (.A(net538),
    .B(net349),
    .Y(_05837_));
 sky130_fd_sc_hd__xor2_2 _14351_ (.A(_05836_),
    .B(_05837_),
    .X(_05838_));
 sky130_fd_sc_hd__a22o_1 _14352_ (.A1(net514),
    .A2(net632),
    .B1(net366),
    .B2(net519),
    .X(_05839_));
 sky130_fd_sc_hd__and4_1 _14353_ (.A(net514),
    .B(net519),
    .C(net632),
    .D(net366),
    .X(_05840_));
 sky130_fd_sc_hd__nand4_1 _14354_ (.A(net514),
    .B(net519),
    .C(net632),
    .D(net366),
    .Y(_05841_));
 sky130_fd_sc_hd__a22o_1 _14355_ (.A1(net523),
    .A2(net361),
    .B1(_05839_),
    .B2(_05841_),
    .X(_05842_));
 sky130_fd_sc_hd__and4_1 _14356_ (.A(net523),
    .B(net361),
    .C(_05839_),
    .D(_05841_),
    .X(_05843_));
 sky130_fd_sc_hd__nand4_1 _14357_ (.A(net523),
    .B(net362),
    .C(_05839_),
    .D(_05841_),
    .Y(_05844_));
 sky130_fd_sc_hd__o211a_1 _14358_ (.A1(_05669_),
    .A2(_05672_),
    .B1(_05842_),
    .C1(_05844_),
    .X(_05845_));
 sky130_fd_sc_hd__a211o_1 _14359_ (.A1(_05842_),
    .A2(_05844_),
    .B1(_05669_),
    .C1(_05672_),
    .X(_05846_));
 sky130_fd_sc_hd__nand2b_1 _14360_ (.A_N(_05845_),
    .B(_05846_),
    .Y(_05847_));
 sky130_fd_sc_hd__xnor2_2 _14361_ (.A(_05838_),
    .B(_05847_),
    .Y(_05848_));
 sky130_fd_sc_hd__nand2_1 _14362_ (.A(_05681_),
    .B(_05683_),
    .Y(_05849_));
 sky130_fd_sc_hd__a21bo_1 _14363_ (.A1(_05699_),
    .A2(_05702_),
    .B1_N(_05700_),
    .X(_05850_));
 sky130_fd_sc_hd__a22o_1 _14364_ (.A1(net504),
    .A2(net377),
    .B1(\mul0.a[18] ),
    .B2(net383),
    .X(_05851_));
 sky130_fd_sc_hd__nand4_2 _14365_ (.A(net504),
    .B(net383),
    .C(net377),
    .D(net499),
    .Y(_05852_));
 sky130_fd_sc_hd__a22o_1 _14366_ (.A1(net508),
    .A2(net374),
    .B1(_05851_),
    .B2(_05852_),
    .X(_05853_));
 sky130_fd_sc_hd__nand4_1 _14367_ (.A(net508),
    .B(net374),
    .C(_05851_),
    .D(_05852_),
    .Y(_05854_));
 sky130_fd_sc_hd__nand3_1 _14368_ (.A(_05850_),
    .B(_05853_),
    .C(_05854_),
    .Y(_05855_));
 sky130_fd_sc_hd__a21o_1 _14369_ (.A1(_05853_),
    .A2(_05854_),
    .B1(_05850_),
    .X(_05856_));
 sky130_fd_sc_hd__nand3_1 _14370_ (.A(_05849_),
    .B(_05855_),
    .C(_05856_),
    .Y(_05857_));
 sky130_fd_sc_hd__a21o_1 _14371_ (.A1(_05855_),
    .A2(_05856_),
    .B1(_05849_),
    .X(_05858_));
 sky130_fd_sc_hd__a21bo_1 _14372_ (.A1(_05678_),
    .A2(_05685_),
    .B1_N(_05684_),
    .X(_05859_));
 sky130_fd_sc_hd__nand3_1 _14373_ (.A(_05857_),
    .B(_05858_),
    .C(_05859_),
    .Y(_05860_));
 sky130_fd_sc_hd__a21o_1 _14374_ (.A1(_05857_),
    .A2(_05858_),
    .B1(_05859_),
    .X(_05861_));
 sky130_fd_sc_hd__and3_1 _14375_ (.A(_05848_),
    .B(_05860_),
    .C(_05861_),
    .X(_05862_));
 sky130_fd_sc_hd__a21oi_1 _14376_ (.A1(_05860_),
    .A2(_05861_),
    .B1(_05848_),
    .Y(_05863_));
 sky130_fd_sc_hd__a211o_1 _14377_ (.A1(_05714_),
    .A2(_05716_),
    .B1(_05862_),
    .C1(_05863_),
    .X(_05864_));
 sky130_fd_sc_hd__o211ai_2 _14378_ (.A1(_05862_),
    .A2(_05863_),
    .B1(_05714_),
    .C1(_05716_),
    .Y(_05865_));
 sky130_fd_sc_hd__and3_1 _14379_ (.A(_05833_),
    .B(_05864_),
    .C(_05865_),
    .X(_05866_));
 sky130_fd_sc_hd__a21oi_1 _14380_ (.A1(_05864_),
    .A2(_05865_),
    .B1(_05833_),
    .Y(_05867_));
 sky130_fd_sc_hd__nor2_2 _14381_ (.A(_05866_),
    .B(_05867_),
    .Y(_05868_));
 sky130_fd_sc_hd__a21o_1 _14382_ (.A1(_05719_),
    .A2(_05726_),
    .B1(_05725_),
    .X(_05869_));
 sky130_fd_sc_hd__a22o_1 _14383_ (.A1(net392),
    .A2(net490),
    .B1(net486),
    .B2(net397),
    .X(_05870_));
 sky130_fd_sc_hd__nand4_1 _14384_ (.A(net397),
    .B(net394),
    .C(net490),
    .D(net486),
    .Y(_05871_));
 sky130_fd_sc_hd__nand2_1 _14385_ (.A(_05870_),
    .B(_05871_),
    .Y(_05872_));
 sky130_fd_sc_hd__and2_1 _14386_ (.A(net387),
    .B(net494),
    .X(_05873_));
 sky130_fd_sc_hd__xnor2_1 _14387_ (.A(_05872_),
    .B(_05873_),
    .Y(_05874_));
 sky130_fd_sc_hd__a22o_1 _14388_ (.A1(net406),
    .A2(net481),
    .B1(net477),
    .B2(net410),
    .X(_05875_));
 sky130_fd_sc_hd__nand4_4 _14389_ (.A(net410),
    .B(net406),
    .C(net479),
    .D(net475),
    .Y(_05876_));
 sky130_fd_sc_hd__a22o_1 _14390_ (.A1(net402),
    .A2(net482),
    .B1(_05875_),
    .B2(_05876_),
    .X(_05877_));
 sky130_fd_sc_hd__nand4_4 _14391_ (.A(net402),
    .B(net482),
    .C(_05875_),
    .D(_05876_),
    .Y(_05878_));
 sky130_fd_sc_hd__a21bo_1 _14392_ (.A1(_05704_),
    .A2(_05706_),
    .B1_N(_05705_),
    .X(_05879_));
 sky130_fd_sc_hd__nand3_2 _14393_ (.A(_05877_),
    .B(_05878_),
    .C(_05879_),
    .Y(_05880_));
 sky130_fd_sc_hd__a21o_1 _14394_ (.A1(_05877_),
    .A2(_05878_),
    .B1(_05879_),
    .X(_05881_));
 sky130_fd_sc_hd__nand3_2 _14395_ (.A(_05874_),
    .B(_05880_),
    .C(_05881_),
    .Y(_05882_));
 sky130_fd_sc_hd__a21o_1 _14396_ (.A1(_05880_),
    .A2(_05881_),
    .B1(_05874_),
    .X(_05883_));
 sky130_fd_sc_hd__and3_1 _14397_ (.A(_05869_),
    .B(_05882_),
    .C(_05883_),
    .X(_05884_));
 sky130_fd_sc_hd__nand3_1 _14398_ (.A(_05869_),
    .B(_05882_),
    .C(_05883_),
    .Y(_05885_));
 sky130_fd_sc_hd__a21oi_1 _14399_ (.A1(_05882_),
    .A2(_05883_),
    .B1(_05869_),
    .Y(_05886_));
 sky130_fd_sc_hd__a211o_1 _14400_ (.A1(_05710_),
    .A2(_05712_),
    .B1(_05884_),
    .C1(_05886_),
    .X(_05887_));
 sky130_fd_sc_hd__o211ai_1 _14401_ (.A1(_05884_),
    .A2(_05886_),
    .B1(_05710_),
    .C1(_05712_),
    .Y(_05888_));
 sky130_fd_sc_hd__and2_2 _14402_ (.A(_05887_),
    .B(_05888_),
    .X(_05889_));
 sky130_fd_sc_hd__nand2_2 _14403_ (.A(_05722_),
    .B(_05724_),
    .Y(_05890_));
 sky130_fd_sc_hd__a32o_1 _14404_ (.A1(net428),
    .A2(net463),
    .A3(_05729_),
    .B1(_05730_),
    .B2(net460),
    .X(_05891_));
 sky130_fd_sc_hd__a22o_1 _14405_ (.A1(net419),
    .A2(net467),
    .B1(net464),
    .B2(net423),
    .X(_05892_));
 sky130_fd_sc_hd__nand4_2 _14406_ (.A(net423),
    .B(net419),
    .C(net467),
    .D(net464),
    .Y(_05893_));
 sky130_fd_sc_hd__a22o_1 _14407_ (.A1(net415),
    .A2(net473),
    .B1(_05892_),
    .B2(_05893_),
    .X(_05894_));
 sky130_fd_sc_hd__nand4_2 _14408_ (.A(net415),
    .B(net473),
    .C(_05892_),
    .D(_05893_),
    .Y(_05895_));
 sky130_fd_sc_hd__and3_1 _14409_ (.A(_05891_),
    .B(_05894_),
    .C(_05895_),
    .X(_05896_));
 sky130_fd_sc_hd__a21o_1 _14410_ (.A1(_05894_),
    .A2(_05895_),
    .B1(_05891_),
    .X(_05897_));
 sky130_fd_sc_hd__and2b_1 _14411_ (.A_N(_05896_),
    .B(_05897_),
    .X(_05898_));
 sky130_fd_sc_hd__xnor2_4 _14412_ (.A(_05890_),
    .B(_05898_),
    .Y(_05899_));
 sky130_fd_sc_hd__a22o_1 _14413_ (.A1(net433),
    .A2(net459),
    .B1(net457),
    .B2(net438),
    .X(_05900_));
 sky130_fd_sc_hd__a21bo_1 _14414_ (.A1(net457),
    .A2(_05730_),
    .B1_N(_05900_),
    .X(_05901_));
 sky130_fd_sc_hd__nand2_2 _14415_ (.A(net428),
    .B(net460),
    .Y(_05902_));
 sky130_fd_sc_hd__xor2_4 _14416_ (.A(_05901_),
    .B(_05902_),
    .X(_05903_));
 sky130_fd_sc_hd__mux2_4 _14417_ (.A0(_05736_),
    .A1(_05737_),
    .S(net442),
    .X(_05904_));
 sky130_fd_sc_hd__xor2_4 _14418_ (.A(_05739_),
    .B(_05904_),
    .X(_05905_));
 sky130_fd_sc_hd__xnor2_4 _14419_ (.A(_05903_),
    .B(_05905_),
    .Y(_05906_));
 sky130_fd_sc_hd__a21bo_1 _14420_ (.A1(_05733_),
    .A2(_05742_),
    .B1_N(_05741_),
    .X(_05907_));
 sky130_fd_sc_hd__nand2b_1 _14421_ (.A_N(_05906_),
    .B(_05907_),
    .Y(_05908_));
 sky130_fd_sc_hd__xor2_4 _14422_ (.A(_05906_),
    .B(_05907_),
    .X(_05909_));
 sky130_fd_sc_hd__xnor2_4 _14423_ (.A(_05899_),
    .B(_05909_),
    .Y(_05910_));
 sky130_fd_sc_hd__a21bo_2 _14424_ (.A1(_05728_),
    .A2(_05747_),
    .B1_N(_05746_),
    .X(_05911_));
 sky130_fd_sc_hd__and2b_1 _14425_ (.A_N(_05910_),
    .B(_05911_),
    .X(_05912_));
 sky130_fd_sc_hd__xnor2_4 _14426_ (.A(_05910_),
    .B(_05911_),
    .Y(_05913_));
 sky130_fd_sc_hd__xnor2_4 _14427_ (.A(_05889_),
    .B(_05913_),
    .Y(_05914_));
 sky130_fd_sc_hd__a21bo_2 _14428_ (.A1(_05718_),
    .A2(_05751_),
    .B1_N(_05750_),
    .X(_05915_));
 sky130_fd_sc_hd__and2b_1 _14429_ (.A_N(_05914_),
    .B(_05915_),
    .X(_05916_));
 sky130_fd_sc_hd__xnor2_4 _14430_ (.A(_05914_),
    .B(_05915_),
    .Y(_05917_));
 sky130_fd_sc_hd__xnor2_4 _14431_ (.A(_05868_),
    .B(_05917_),
    .Y(_05918_));
 sky130_fd_sc_hd__a21bo_2 _14432_ (.A1(_05696_),
    .A2(_05755_),
    .B1_N(_05754_),
    .X(_05919_));
 sky130_fd_sc_hd__and2b_1 _14433_ (.A_N(_05918_),
    .B(_05919_),
    .X(_05920_));
 sky130_fd_sc_hd__xnor2_4 _14434_ (.A(_05918_),
    .B(_05919_),
    .Y(_05921_));
 sky130_fd_sc_hd__xor2_2 _14435_ (.A(_05832_),
    .B(_05921_),
    .X(_05922_));
 sky130_fd_sc_hd__a21oi_2 _14436_ (.A1(_05661_),
    .A2(_05760_),
    .B1(_05758_),
    .Y(_05923_));
 sky130_fd_sc_hd__and2b_1 _14437_ (.A_N(_05923_),
    .B(_05922_),
    .X(_05924_));
 sky130_fd_sc_hd__xnor2_2 _14438_ (.A(_05922_),
    .B(_05923_),
    .Y(_05925_));
 sky130_fd_sc_hd__xnor2_2 _14439_ (.A(_05789_),
    .B(_05925_),
    .Y(_05926_));
 sky130_fd_sc_hd__a21boi_4 _14440_ (.A1(_05618_),
    .A2(_05764_),
    .B1_N(_05763_),
    .Y(_05927_));
 sky130_fd_sc_hd__nor2_1 _14441_ (.A(_05926_),
    .B(_05927_),
    .Y(_05928_));
 sky130_fd_sc_hd__xor2_2 _14442_ (.A(_05926_),
    .B(_05927_),
    .X(_05929_));
 sky130_fd_sc_hd__xor2_2 _14443_ (.A(_05788_),
    .B(_05929_),
    .X(_05930_));
 sky130_fd_sc_hd__o21ai_2 _14444_ (.A1(_05769_),
    .A2(_05771_),
    .B1(_05930_),
    .Y(_05931_));
 sky130_fd_sc_hd__inv_2 _14445_ (.A(_05931_),
    .Y(_05932_));
 sky130_fd_sc_hd__nor3_2 _14446_ (.A(_05769_),
    .B(_05771_),
    .C(_05930_),
    .Y(_05933_));
 sky130_fd_sc_hd__nor2_2 _14447_ (.A(_05932_),
    .B(_05933_),
    .Y(_05934_));
 sky130_fd_sc_hd__xnor2_4 _14448_ (.A(_05787_),
    .B(_05934_),
    .Y(_05935_));
 sky130_fd_sc_hd__nor2_1 _14449_ (.A(net9),
    .B(_05935_),
    .Y(_05936_));
 sky130_fd_sc_hd__a221o_1 _14450_ (.A1(net599),
    .A2(net703),
    .B1(_02648_),
    .B2(net6),
    .C1(_05936_),
    .X(_05937_));
 sky130_fd_sc_hd__mux2_1 _14451_ (.A0(net889),
    .A1(_05937_),
    .S(net3),
    .X(_00283_));
 sky130_fd_sc_hd__a21o_1 _14452_ (.A1(_05621_),
    .A2(_05807_),
    .B1(_05805_),
    .X(_05938_));
 sky130_fd_sc_hd__or2_2 _14453_ (.A(_05829_),
    .B(_05831_),
    .X(_05939_));
 sky130_fd_sc_hd__o21ba_2 _14454_ (.A1(_05808_),
    .A2(_05827_),
    .B1_N(_05826_),
    .X(_05940_));
 sky130_fd_sc_hd__a21bo_2 _14455_ (.A1(_05833_),
    .A2(_05865_),
    .B1_N(_05864_),
    .X(_05941_));
 sky130_fd_sc_hd__a22o_1 _14456_ (.A1(net551),
    .A2(net335),
    .B1(net332),
    .B2(net555),
    .X(_05942_));
 sky130_fd_sc_hd__and3_1 _14457_ (.A(net551),
    .B(net556),
    .C(net332),
    .X(_05943_));
 sky130_fd_sc_hd__a21bo_2 _14458_ (.A1(net335),
    .A2(_05943_),
    .B1_N(_05942_),
    .X(_05944_));
 sky130_fd_sc_hd__nand2_2 _14459_ (.A(net560),
    .B(net329),
    .Y(_05945_));
 sky130_fd_sc_hd__xnor2_4 _14460_ (.A(_05944_),
    .B(_05945_),
    .Y(_05946_));
 sky130_fd_sc_hd__o2bb2a_2 _14461_ (.A1_N(net335),
    .A2_N(_05793_),
    .B1(_05794_),
    .B2(_05795_),
    .X(_05947_));
 sky130_fd_sc_hd__xnor2_2 _14462_ (.A(_05946_),
    .B(_05947_),
    .Y(_05948_));
 sky130_fd_sc_hd__and4b_2 _14463_ (.A_N(net569),
    .B(net328),
    .C(net326),
    .D(net563),
    .X(_05949_));
 sky130_fd_sc_hd__inv_2 _14464_ (.A(_05949_),
    .Y(_05950_));
 sky130_fd_sc_hd__o2bb2a_1 _14465_ (.A1_N(net563),
    .A2_N(net328),
    .B1(net57),
    .B2(net569),
    .X(_05951_));
 sky130_fd_sc_hd__nor2_1 _14466_ (.A(_05949_),
    .B(_05951_),
    .Y(_05952_));
 sky130_fd_sc_hd__xnor2_1 _14467_ (.A(_05948_),
    .B(_05952_),
    .Y(_05953_));
 sky130_fd_sc_hd__o32ai_4 _14468_ (.A1(_05798_),
    .A2(_05799_),
    .A3(_05801_),
    .B1(_05797_),
    .B2(_05796_),
    .Y(_05954_));
 sky130_fd_sc_hd__xnor2_1 _14469_ (.A(_05953_),
    .B(_05954_),
    .Y(_05955_));
 sky130_fd_sc_hd__nor2_1 _14470_ (.A(_05800_),
    .B(_05955_),
    .Y(_05956_));
 sky130_fd_sc_hd__and2_1 _14471_ (.A(_05800_),
    .B(_05955_),
    .X(_05957_));
 sky130_fd_sc_hd__or2_2 _14472_ (.A(_05956_),
    .B(_05957_),
    .X(_05958_));
 sky130_fd_sc_hd__a21oi_1 _14473_ (.A1(_05838_),
    .A2(_05846_),
    .B1(_05845_),
    .Y(_05959_));
 sky130_fd_sc_hd__nand2_1 _14474_ (.A(_05813_),
    .B(_05815_),
    .Y(_05960_));
 sky130_fd_sc_hd__a32o_1 _14475_ (.A1(net538),
    .A2(net349),
    .A3(_05834_),
    .B1(_05835_),
    .B2(net356),
    .X(_05961_));
 sky130_fd_sc_hd__a22o_1 _14476_ (.A1(net538),
    .A2(net345),
    .B1(net341),
    .B2(net543),
    .X(_05962_));
 sky130_fd_sc_hd__nand4_2 _14477_ (.A(net538),
    .B(net543),
    .C(net345),
    .D(net341),
    .Y(_05963_));
 sky130_fd_sc_hd__a22o_1 _14478_ (.A1(net547),
    .A2(net339),
    .B1(_05962_),
    .B2(_05963_),
    .X(_05964_));
 sky130_fd_sc_hd__nand4_2 _14479_ (.A(net547),
    .B(net339),
    .C(_05962_),
    .D(_05963_),
    .Y(_05965_));
 sky130_fd_sc_hd__nand3_2 _14480_ (.A(_05961_),
    .B(_05964_),
    .C(_05965_),
    .Y(_05966_));
 sky130_fd_sc_hd__a21o_1 _14481_ (.A1(_05964_),
    .A2(_05965_),
    .B1(_05961_),
    .X(_05967_));
 sky130_fd_sc_hd__nand3_2 _14482_ (.A(_05960_),
    .B(_05966_),
    .C(_05967_),
    .Y(_05968_));
 sky130_fd_sc_hd__a21o_1 _14483_ (.A1(_05966_),
    .A2(_05967_),
    .B1(_05960_),
    .X(_05969_));
 sky130_fd_sc_hd__and3b_1 _14484_ (.A_N(_05959_),
    .B(_05968_),
    .C(_05969_),
    .X(_05970_));
 sky130_fd_sc_hd__a21boi_1 _14485_ (.A1(_05968_),
    .A2(_05969_),
    .B1_N(_05959_),
    .Y(_05971_));
 sky130_fd_sc_hd__a211oi_1 _14486_ (.A1(_05816_),
    .A2(_05818_),
    .B1(_05970_),
    .C1(_05971_),
    .Y(_05972_));
 sky130_fd_sc_hd__o211ai_1 _14487_ (.A1(_05970_),
    .A2(_05971_),
    .B1(_05816_),
    .C1(_05818_),
    .Y(_05973_));
 sky130_fd_sc_hd__nand2b_2 _14488_ (.A_N(_05972_),
    .B(_05973_),
    .Y(_05974_));
 sky130_fd_sc_hd__nor2_2 _14489_ (.A(_05820_),
    .B(_05822_),
    .Y(_05975_));
 sky130_fd_sc_hd__nor2_1 _14490_ (.A(_05974_),
    .B(_05975_),
    .Y(_05976_));
 sky130_fd_sc_hd__xnor2_4 _14491_ (.A(_05974_),
    .B(_05975_),
    .Y(_05977_));
 sky130_fd_sc_hd__xnor2_4 _14492_ (.A(_05958_),
    .B(_05977_),
    .Y(_05978_));
 sky130_fd_sc_hd__and2b_1 _14493_ (.A_N(_05978_),
    .B(_05941_),
    .X(_05979_));
 sky130_fd_sc_hd__xnor2_4 _14494_ (.A(_05941_),
    .B(_05978_),
    .Y(_05980_));
 sky130_fd_sc_hd__and2b_1 _14495_ (.A_N(_05940_),
    .B(_05980_),
    .X(_05981_));
 sky130_fd_sc_hd__xnor2_4 _14496_ (.A(_05940_),
    .B(_05980_),
    .Y(_05982_));
 sky130_fd_sc_hd__a31o_2 _14497_ (.A1(_05857_),
    .A2(_05858_),
    .A3(_05859_),
    .B1(_05862_),
    .X(_05983_));
 sky130_fd_sc_hd__a22o_1 _14498_ (.A1(net523),
    .A2(net357),
    .B1(net352),
    .B2(net529),
    .X(_05984_));
 sky130_fd_sc_hd__and3_1 _14499_ (.A(net523),
    .B(net529),
    .C(net352),
    .X(_05985_));
 sky130_fd_sc_hd__a21bo_1 _14500_ (.A1(net356),
    .A2(_05985_),
    .B1_N(_05984_),
    .X(_05986_));
 sky130_fd_sc_hd__nand2_1 _14501_ (.A(net533),
    .B(net349),
    .Y(_05987_));
 sky130_fd_sc_hd__xor2_2 _14502_ (.A(_05986_),
    .B(_05987_),
    .X(_05988_));
 sky130_fd_sc_hd__a22o_1 _14503_ (.A1(net510),
    .A2(net632),
    .B1(net366),
    .B2(net514),
    .X(_05989_));
 sky130_fd_sc_hd__and4_1 _14504_ (.A(net509),
    .B(net514),
    .C(net633),
    .D(net366),
    .X(_05990_));
 sky130_fd_sc_hd__nand4_1 _14505_ (.A(net510),
    .B(net514),
    .C(net633),
    .D(net366),
    .Y(_05991_));
 sky130_fd_sc_hd__a22o_1 _14506_ (.A1(net519),
    .A2(net361),
    .B1(_05989_),
    .B2(_05991_),
    .X(_05992_));
 sky130_fd_sc_hd__and4_1 _14507_ (.A(net519),
    .B(net361),
    .C(_05989_),
    .D(_05991_),
    .X(_05993_));
 sky130_fd_sc_hd__nand4_1 _14508_ (.A(net519),
    .B(net361),
    .C(_05989_),
    .D(_05991_),
    .Y(_05994_));
 sky130_fd_sc_hd__o211a_1 _14509_ (.A1(_05840_),
    .A2(_05843_),
    .B1(_05992_),
    .C1(_05994_),
    .X(_05995_));
 sky130_fd_sc_hd__a211o_1 _14510_ (.A1(_05992_),
    .A2(_05994_),
    .B1(_05840_),
    .C1(_05843_),
    .X(_05996_));
 sky130_fd_sc_hd__nand2b_1 _14511_ (.A_N(_05995_),
    .B(_05996_),
    .Y(_05997_));
 sky130_fd_sc_hd__xnor2_2 _14512_ (.A(_05988_),
    .B(_05997_),
    .Y(_05998_));
 sky130_fd_sc_hd__nand2_1 _14513_ (.A(_05852_),
    .B(_05854_),
    .Y(_05999_));
 sky130_fd_sc_hd__a21bo_1 _14514_ (.A1(_05870_),
    .A2(_05873_),
    .B1_N(_05871_),
    .X(_06000_));
 sky130_fd_sc_hd__a22o_1 _14515_ (.A1(net377),
    .A2(net502),
    .B1(net497),
    .B2(net385),
    .X(_06001_));
 sky130_fd_sc_hd__nand4_2 _14516_ (.A(net383),
    .B(net380),
    .C(net502),
    .D(net497),
    .Y(_06002_));
 sky130_fd_sc_hd__a22o_1 _14517_ (.A1(net504),
    .A2(net372),
    .B1(_06001_),
    .B2(_06002_),
    .X(_06003_));
 sky130_fd_sc_hd__nand4_2 _14518_ (.A(\mul0.a[17] ),
    .B(net372),
    .C(_06001_),
    .D(_06002_),
    .Y(_06004_));
 sky130_fd_sc_hd__nand3_1 _14519_ (.A(_06000_),
    .B(_06003_),
    .C(_06004_),
    .Y(_06005_));
 sky130_fd_sc_hd__a21o_1 _14520_ (.A1(_06003_),
    .A2(_06004_),
    .B1(_06000_),
    .X(_06006_));
 sky130_fd_sc_hd__nand3_1 _14521_ (.A(_05999_),
    .B(_06005_),
    .C(_06006_),
    .Y(_06007_));
 sky130_fd_sc_hd__a21o_1 _14522_ (.A1(_06005_),
    .A2(_06006_),
    .B1(_05999_),
    .X(_06008_));
 sky130_fd_sc_hd__a21bo_1 _14523_ (.A1(_05849_),
    .A2(_05856_),
    .B1_N(_05855_),
    .X(_06009_));
 sky130_fd_sc_hd__nand3_1 _14524_ (.A(_06007_),
    .B(_06008_),
    .C(_06009_),
    .Y(_06010_));
 sky130_fd_sc_hd__a21o_1 _14525_ (.A1(_06007_),
    .A2(_06008_),
    .B1(_06009_),
    .X(_06011_));
 sky130_fd_sc_hd__and3_1 _14526_ (.A(_05998_),
    .B(_06010_),
    .C(_06011_),
    .X(_06012_));
 sky130_fd_sc_hd__a21oi_1 _14527_ (.A1(_06010_),
    .A2(_06011_),
    .B1(_05998_),
    .Y(_06013_));
 sky130_fd_sc_hd__a211oi_2 _14528_ (.A1(_05885_),
    .A2(_05887_),
    .B1(_06012_),
    .C1(_06013_),
    .Y(_06014_));
 sky130_fd_sc_hd__o211a_1 _14529_ (.A1(_06012_),
    .A2(_06013_),
    .B1(_05885_),
    .C1(_05887_),
    .X(_06015_));
 sky130_fd_sc_hd__nor2_2 _14530_ (.A(_06014_),
    .B(_06015_),
    .Y(_06016_));
 sky130_fd_sc_hd__xor2_4 _14531_ (.A(_05983_),
    .B(_06016_),
    .X(_06017_));
 sky130_fd_sc_hd__nand2_1 _14532_ (.A(_05880_),
    .B(_05882_),
    .Y(_06018_));
 sky130_fd_sc_hd__a21o_1 _14533_ (.A1(_05890_),
    .A2(_05897_),
    .B1(_05896_),
    .X(_06019_));
 sky130_fd_sc_hd__a22o_1 _14534_ (.A1(net392),
    .A2(net488),
    .B1(net484),
    .B2(net399),
    .X(_06020_));
 sky130_fd_sc_hd__and3_1 _14535_ (.A(net399),
    .B(net394),
    .C(net488),
    .X(_06021_));
 sky130_fd_sc_hd__a21bo_1 _14536_ (.A1(net484),
    .A2(_06021_),
    .B1_N(_06020_),
    .X(_06022_));
 sky130_fd_sc_hd__nand2_1 _14537_ (.A(net387),
    .B(net493),
    .Y(_06023_));
 sky130_fd_sc_hd__xor2_1 _14538_ (.A(_06022_),
    .B(_06023_),
    .X(_06024_));
 sky130_fd_sc_hd__a22o_1 _14539_ (.A1(net406),
    .A2(net475),
    .B1(net471),
    .B2(net412),
    .X(_06025_));
 sky130_fd_sc_hd__nand4_2 _14540_ (.A(net410),
    .B(net406),
    .C(net475),
    .D(net471),
    .Y(_06026_));
 sky130_fd_sc_hd__inv_2 _14541_ (.A(_06026_),
    .Y(_06027_));
 sky130_fd_sc_hd__a22oi_2 _14542_ (.A1(net402),
    .A2(net479),
    .B1(_06025_),
    .B2(_06026_),
    .Y(_06028_));
 sky130_fd_sc_hd__and4_2 _14543_ (.A(net402),
    .B(net479),
    .C(_06025_),
    .D(_06026_),
    .X(_06029_));
 sky130_fd_sc_hd__a211o_2 _14544_ (.A1(_05876_),
    .A2(_05878_),
    .B1(_06028_),
    .C1(_06029_),
    .X(_06030_));
 sky130_fd_sc_hd__o211ai_2 _14545_ (.A1(_06028_),
    .A2(_06029_),
    .B1(_05876_),
    .C1(_05878_),
    .Y(_06031_));
 sky130_fd_sc_hd__nand3_2 _14546_ (.A(_06024_),
    .B(_06030_),
    .C(_06031_),
    .Y(_06032_));
 sky130_fd_sc_hd__a21o_1 _14547_ (.A1(_06030_),
    .A2(_06031_),
    .B1(_06024_),
    .X(_06033_));
 sky130_fd_sc_hd__nand3_1 _14548_ (.A(_06019_),
    .B(_06032_),
    .C(_06033_),
    .Y(_06034_));
 sky130_fd_sc_hd__inv_2 _14549_ (.A(_06034_),
    .Y(_06035_));
 sky130_fd_sc_hd__a21o_1 _14550_ (.A1(_06032_),
    .A2(_06033_),
    .B1(_06019_),
    .X(_06036_));
 sky130_fd_sc_hd__and3_1 _14551_ (.A(_06018_),
    .B(_06034_),
    .C(_06036_),
    .X(_06037_));
 sky130_fd_sc_hd__a21oi_1 _14552_ (.A1(_06034_),
    .A2(_06036_),
    .B1(_06018_),
    .Y(_06038_));
 sky130_fd_sc_hd__nor2_2 _14553_ (.A(_06037_),
    .B(_06038_),
    .Y(_06039_));
 sky130_fd_sc_hd__nand2_2 _14554_ (.A(_05893_),
    .B(_05895_),
    .Y(_06040_));
 sky130_fd_sc_hd__a32o_1 _14555_ (.A1(net428),
    .A2(net460),
    .A3(_05900_),
    .B1(_05730_),
    .B2(net457),
    .X(_06041_));
 sky130_fd_sc_hd__a22o_1 _14556_ (.A1(net419),
    .A2(net464),
    .B1(net460),
    .B2(net423),
    .X(_06042_));
 sky130_fd_sc_hd__nand4_2 _14557_ (.A(net423),
    .B(net419),
    .C(net464),
    .D(net460),
    .Y(_06043_));
 sky130_fd_sc_hd__a22o_1 _14558_ (.A1(net415),
    .A2(net466),
    .B1(_06042_),
    .B2(_06043_),
    .X(_06044_));
 sky130_fd_sc_hd__nand4_2 _14559_ (.A(net415),
    .B(net467),
    .C(_06042_),
    .D(_06043_),
    .Y(_06045_));
 sky130_fd_sc_hd__and3_1 _14560_ (.A(_06041_),
    .B(_06044_),
    .C(_06045_),
    .X(_06046_));
 sky130_fd_sc_hd__a21o_1 _14561_ (.A1(_06044_),
    .A2(_06045_),
    .B1(_06041_),
    .X(_06047_));
 sky130_fd_sc_hd__and2b_1 _14562_ (.A_N(_06046_),
    .B(_06047_),
    .X(_06048_));
 sky130_fd_sc_hd__xor2_4 _14563_ (.A(_06040_),
    .B(_06048_),
    .X(_06049_));
 sky130_fd_sc_hd__a22o_1 _14564_ (.A1(net433),
    .A2(net456),
    .B1(net453),
    .B2(net438),
    .X(_06050_));
 sky130_fd_sc_hd__nand4_1 _14565_ (.A(net439),
    .B(net434),
    .C(net456),
    .D(net453),
    .Y(_06051_));
 sky130_fd_sc_hd__and2_1 _14566_ (.A(net429),
    .B(net459),
    .X(_06052_));
 sky130_fd_sc_hd__a21o_1 _14567_ (.A1(_06050_),
    .A2(_06051_),
    .B1(_06052_),
    .X(_06053_));
 sky130_fd_sc_hd__nand3_1 _14568_ (.A(_06050_),
    .B(_06051_),
    .C(_06052_),
    .Y(_06054_));
 sky130_fd_sc_hd__o211a_1 _14569_ (.A1(_05739_),
    .A2(_05904_),
    .B1(_06053_),
    .C1(_06054_),
    .X(_06055_));
 sky130_fd_sc_hd__a211oi_1 _14570_ (.A1(_06053_),
    .A2(_06054_),
    .B1(_05739_),
    .C1(_05904_),
    .Y(_06056_));
 sky130_fd_sc_hd__nor2_2 _14571_ (.A(_06055_),
    .B(_06056_),
    .Y(_06057_));
 sky130_fd_sc_hd__and2_2 _14572_ (.A(net442),
    .B(_05736_),
    .X(_06058_));
 sky130_fd_sc_hd__a21oi_2 _14573_ (.A1(_05903_),
    .A2(_05905_),
    .B1(_06058_),
    .Y(_06059_));
 sky130_fd_sc_hd__and2b_1 _14574_ (.A_N(_06059_),
    .B(_06057_),
    .X(_06060_));
 sky130_fd_sc_hd__xnor2_4 _14575_ (.A(_06057_),
    .B(_06059_),
    .Y(_06061_));
 sky130_fd_sc_hd__xor2_4 _14576_ (.A(_06049_),
    .B(_06061_),
    .X(_06062_));
 sky130_fd_sc_hd__o21a_2 _14577_ (.A1(_05899_),
    .A2(_05909_),
    .B1(_05908_),
    .X(_06063_));
 sky130_fd_sc_hd__and2b_1 _14578_ (.A_N(_06063_),
    .B(_06062_),
    .X(_06064_));
 sky130_fd_sc_hd__xnor2_4 _14579_ (.A(_06062_),
    .B(_06063_),
    .Y(_06065_));
 sky130_fd_sc_hd__xor2_4 _14580_ (.A(_06039_),
    .B(_06065_),
    .X(_06066_));
 sky130_fd_sc_hd__a21o_2 _14581_ (.A1(_05889_),
    .A2(_05913_),
    .B1(_05912_),
    .X(_06067_));
 sky130_fd_sc_hd__nand2_1 _14582_ (.A(_06066_),
    .B(_06067_),
    .Y(_06068_));
 sky130_fd_sc_hd__xor2_4 _14583_ (.A(_06066_),
    .B(_06067_),
    .X(_06069_));
 sky130_fd_sc_hd__xnor2_4 _14584_ (.A(_06017_),
    .B(_06069_),
    .Y(_06070_));
 sky130_fd_sc_hd__a21oi_4 _14585_ (.A1(_05868_),
    .A2(_05917_),
    .B1(_05916_),
    .Y(_06071_));
 sky130_fd_sc_hd__nor2_1 _14586_ (.A(_06070_),
    .B(_06071_),
    .Y(_06072_));
 sky130_fd_sc_hd__xor2_4 _14587_ (.A(_06070_),
    .B(_06071_),
    .X(_06073_));
 sky130_fd_sc_hd__xor2_4 _14588_ (.A(_05982_),
    .B(_06073_),
    .X(_06074_));
 sky130_fd_sc_hd__a21oi_4 _14589_ (.A1(_05832_),
    .A2(_05921_),
    .B1(_05920_),
    .Y(_06075_));
 sky130_fd_sc_hd__nand2b_1 _14590_ (.A_N(_06075_),
    .B(_06074_),
    .Y(_06076_));
 sky130_fd_sc_hd__xnor2_4 _14591_ (.A(_06074_),
    .B(_06075_),
    .Y(_06077_));
 sky130_fd_sc_hd__xnor2_2 _14592_ (.A(_05939_),
    .B(_06077_),
    .Y(_06078_));
 sky130_fd_sc_hd__a21oi_2 _14593_ (.A1(_05789_),
    .A2(_05925_),
    .B1(_05924_),
    .Y(_06079_));
 sky130_fd_sc_hd__nor2_1 _14594_ (.A(_06078_),
    .B(_06079_),
    .Y(_06080_));
 sky130_fd_sc_hd__xor2_2 _14595_ (.A(_06078_),
    .B(_06079_),
    .X(_06081_));
 sky130_fd_sc_hd__xnor2_1 _14596_ (.A(_05938_),
    .B(_06081_),
    .Y(_06082_));
 sky130_fd_sc_hd__a21oi_1 _14597_ (.A1(_05788_),
    .A2(_05929_),
    .B1(_05928_),
    .Y(_06083_));
 sky130_fd_sc_hd__nor2_1 _14598_ (.A(_06082_),
    .B(_06083_),
    .Y(_06084_));
 sky130_fd_sc_hd__xor2_1 _14599_ (.A(_06082_),
    .B(_06083_),
    .X(_06085_));
 sky130_fd_sc_hd__a21oi_2 _14600_ (.A1(_05774_),
    .A2(_05931_),
    .B1(_05933_),
    .Y(_06086_));
 sky130_fd_sc_hd__and3b_1 _14601_ (.A_N(_05783_),
    .B(_05934_),
    .C(_05776_),
    .X(_06087_));
 sky130_fd_sc_hd__o21a_1 _14602_ (.A1(_06086_),
    .A2(_06087_),
    .B1(_06085_),
    .X(_06088_));
 sky130_fd_sc_hd__nor3_1 _14603_ (.A(_06085_),
    .B(_06086_),
    .C(_06087_),
    .Y(_06089_));
 sky130_fd_sc_hd__or2_4 _14604_ (.A(_06088_),
    .B(_06089_),
    .X(_06090_));
 sky130_fd_sc_hd__nor2_1 _14605_ (.A(net9),
    .B(_06090_),
    .Y(_06091_));
 sky130_fd_sc_hd__a221o_1 _14606_ (.A1(net599),
    .A2(net757),
    .B1(_02653_),
    .B2(net6),
    .C1(_06091_),
    .X(_06092_));
 sky130_fd_sc_hd__mux2_1 _14607_ (.A0(net862),
    .A1(_06092_),
    .S(net4),
    .X(_00284_));
 sky130_fd_sc_hd__or2_2 _14608_ (.A(_06084_),
    .B(_06088_),
    .X(_06093_));
 sky130_fd_sc_hd__a21oi_4 _14609_ (.A1(_05938_),
    .A2(_06081_),
    .B1(_06080_),
    .Y(_06094_));
 sky130_fd_sc_hd__a21o_2 _14610_ (.A1(_05953_),
    .A2(_05954_),
    .B1(_05956_),
    .X(_06095_));
 sky130_fd_sc_hd__or2_2 _14611_ (.A(_05979_),
    .B(_05981_),
    .X(_06096_));
 sky130_fd_sc_hd__o21ba_2 _14612_ (.A1(_05958_),
    .A2(_05977_),
    .B1_N(_05976_),
    .X(_06097_));
 sky130_fd_sc_hd__a21o_2 _14613_ (.A1(_05983_),
    .A2(_06016_),
    .B1(_06014_),
    .X(_06098_));
 sky130_fd_sc_hd__a22o_1 _14614_ (.A1(net547),
    .A2(net334),
    .B1(net331),
    .B2(net551),
    .X(_06099_));
 sky130_fd_sc_hd__and3_1 _14615_ (.A(net547),
    .B(net551),
    .C(net331),
    .X(_06100_));
 sky130_fd_sc_hd__a21bo_2 _14616_ (.A1(net334),
    .A2(_06100_),
    .B1_N(_06099_),
    .X(_06101_));
 sky130_fd_sc_hd__nand2_2 _14617_ (.A(net556),
    .B(net329),
    .Y(_06102_));
 sky130_fd_sc_hd__xnor2_4 _14618_ (.A(_06101_),
    .B(_06102_),
    .Y(_06103_));
 sky130_fd_sc_hd__o2bb2a_2 _14619_ (.A1_N(net335),
    .A2_N(_05943_),
    .B1(_05944_),
    .B2(_05945_),
    .X(_06104_));
 sky130_fd_sc_hd__xnor2_2 _14620_ (.A(_06103_),
    .B(_06104_),
    .Y(_06105_));
 sky130_fd_sc_hd__and4b_2 _14621_ (.A_N(net563),
    .B(net327),
    .C(net326),
    .D(net560),
    .X(_06106_));
 sky130_fd_sc_hd__inv_2 _14622_ (.A(_06106_),
    .Y(_06107_));
 sky130_fd_sc_hd__o2bb2a_1 _14623_ (.A1_N(net560),
    .A2_N(net327),
    .B1(net57),
    .B2(net563),
    .X(_06108_));
 sky130_fd_sc_hd__nor2_1 _14624_ (.A(_06106_),
    .B(_06108_),
    .Y(_06109_));
 sky130_fd_sc_hd__xnor2_1 _14625_ (.A(_06105_),
    .B(_06109_),
    .Y(_06110_));
 sky130_fd_sc_hd__o32ai_4 _14626_ (.A1(_05948_),
    .A2(_05949_),
    .A3(_05951_),
    .B1(_05947_),
    .B2(_05946_),
    .Y(_06111_));
 sky130_fd_sc_hd__xnor2_1 _14627_ (.A(_06110_),
    .B(_06111_),
    .Y(_06112_));
 sky130_fd_sc_hd__nor2_1 _14628_ (.A(_05950_),
    .B(_06112_),
    .Y(_06113_));
 sky130_fd_sc_hd__and2_1 _14629_ (.A(_05950_),
    .B(_06112_),
    .X(_06114_));
 sky130_fd_sc_hd__or2_2 _14630_ (.A(_06113_),
    .B(_06114_),
    .X(_06115_));
 sky130_fd_sc_hd__a21oi_1 _14631_ (.A1(_05988_),
    .A2(_05996_),
    .B1(_05995_),
    .Y(_06116_));
 sky130_fd_sc_hd__nand2_1 _14632_ (.A(_05963_),
    .B(_05965_),
    .Y(_06117_));
 sky130_fd_sc_hd__a32o_1 _14633_ (.A1(net533),
    .A2(net349),
    .A3(_05984_),
    .B1(_05985_),
    .B2(net357),
    .X(_06118_));
 sky130_fd_sc_hd__a22o_1 _14634_ (.A1(net534),
    .A2(net346),
    .B1(net342),
    .B2(net538),
    .X(_06119_));
 sky130_fd_sc_hd__nand4_2 _14635_ (.A(net534),
    .B(net538),
    .C(net346),
    .D(net341),
    .Y(_06120_));
 sky130_fd_sc_hd__a22o_1 _14636_ (.A1(net543),
    .A2(net338),
    .B1(_06119_),
    .B2(_06120_),
    .X(_06121_));
 sky130_fd_sc_hd__nand4_2 _14637_ (.A(net543),
    .B(net338),
    .C(_06119_),
    .D(_06120_),
    .Y(_06122_));
 sky130_fd_sc_hd__nand3_2 _14638_ (.A(_06118_),
    .B(_06121_),
    .C(_06122_),
    .Y(_06123_));
 sky130_fd_sc_hd__a21o_1 _14639_ (.A1(_06121_),
    .A2(_06122_),
    .B1(_06118_),
    .X(_06124_));
 sky130_fd_sc_hd__nand3_2 _14640_ (.A(_06117_),
    .B(_06123_),
    .C(_06124_),
    .Y(_06125_));
 sky130_fd_sc_hd__a21o_1 _14641_ (.A1(_06123_),
    .A2(_06124_),
    .B1(_06117_),
    .X(_06126_));
 sky130_fd_sc_hd__and3b_1 _14642_ (.A_N(_06116_),
    .B(_06125_),
    .C(_06126_),
    .X(_06127_));
 sky130_fd_sc_hd__a21boi_1 _14643_ (.A1(_06125_),
    .A2(_06126_),
    .B1_N(_06116_),
    .Y(_06128_));
 sky130_fd_sc_hd__a211oi_1 _14644_ (.A1(_05966_),
    .A2(_05968_),
    .B1(_06127_),
    .C1(_06128_),
    .Y(_06129_));
 sky130_fd_sc_hd__o211ai_1 _14645_ (.A1(_06127_),
    .A2(_06128_),
    .B1(_05966_),
    .C1(_05968_),
    .Y(_06130_));
 sky130_fd_sc_hd__nand2b_2 _14646_ (.A_N(_06129_),
    .B(_06130_),
    .Y(_06131_));
 sky130_fd_sc_hd__nor2_2 _14647_ (.A(_05970_),
    .B(_05972_),
    .Y(_06132_));
 sky130_fd_sc_hd__nor2_1 _14648_ (.A(_06131_),
    .B(_06132_),
    .Y(_06133_));
 sky130_fd_sc_hd__xnor2_4 _14649_ (.A(_06131_),
    .B(_06132_),
    .Y(_06134_));
 sky130_fd_sc_hd__xnor2_4 _14650_ (.A(_06115_),
    .B(_06134_),
    .Y(_06135_));
 sky130_fd_sc_hd__and2b_1 _14651_ (.A_N(_06135_),
    .B(_06098_),
    .X(_06136_));
 sky130_fd_sc_hd__xnor2_4 _14652_ (.A(_06098_),
    .B(_06135_),
    .Y(_06137_));
 sky130_fd_sc_hd__and2b_1 _14653_ (.A_N(_06097_),
    .B(_06137_),
    .X(_06138_));
 sky130_fd_sc_hd__xnor2_4 _14654_ (.A(_06097_),
    .B(_06137_),
    .Y(_06139_));
 sky130_fd_sc_hd__a31o_2 _14655_ (.A1(_06007_),
    .A2(_06008_),
    .A3(_06009_),
    .B1(_06012_),
    .X(_06140_));
 sky130_fd_sc_hd__a22o_1 _14656_ (.A1(net518),
    .A2(net357),
    .B1(net352),
    .B2(net522),
    .X(_06141_));
 sky130_fd_sc_hd__and3_1 _14657_ (.A(net518),
    .B(net522),
    .C(net352),
    .X(_06142_));
 sky130_fd_sc_hd__a21bo_1 _14658_ (.A1(net357),
    .A2(_06142_),
    .B1_N(_06141_),
    .X(_06143_));
 sky130_fd_sc_hd__nand2_1 _14659_ (.A(net529),
    .B(net349),
    .Y(_06144_));
 sky130_fd_sc_hd__xor2_2 _14660_ (.A(_06143_),
    .B(_06144_),
    .X(_06145_));
 sky130_fd_sc_hd__a22o_1 _14661_ (.A1(net506),
    .A2(net633),
    .B1(net366),
    .B2(net510),
    .X(_06146_));
 sky130_fd_sc_hd__and4_1 _14662_ (.A(net506),
    .B(net510),
    .C(net633),
    .D(net366),
    .X(_06147_));
 sky130_fd_sc_hd__nand4_1 _14663_ (.A(net505),
    .B(net510),
    .C(net633),
    .D(net367),
    .Y(_06148_));
 sky130_fd_sc_hd__a22o_1 _14664_ (.A1(net514),
    .A2(net361),
    .B1(_06146_),
    .B2(_06148_),
    .X(_06149_));
 sky130_fd_sc_hd__and4_1 _14665_ (.A(net514),
    .B(net361),
    .C(_06146_),
    .D(_06148_),
    .X(_06150_));
 sky130_fd_sc_hd__nand4_1 _14666_ (.A(net514),
    .B(net361),
    .C(_06146_),
    .D(_06148_),
    .Y(_06151_));
 sky130_fd_sc_hd__o211a_1 _14667_ (.A1(_05990_),
    .A2(_05993_),
    .B1(_06149_),
    .C1(_06151_),
    .X(_06152_));
 sky130_fd_sc_hd__a211o_1 _14668_ (.A1(_06149_),
    .A2(_06151_),
    .B1(_05990_),
    .C1(_05993_),
    .X(_06153_));
 sky130_fd_sc_hd__nand2b_1 _14669_ (.A_N(_06152_),
    .B(_06153_),
    .Y(_06154_));
 sky130_fd_sc_hd__xnor2_2 _14670_ (.A(_06145_),
    .B(_06154_),
    .Y(_06155_));
 sky130_fd_sc_hd__nand2_1 _14671_ (.A(_06002_),
    .B(_06004_),
    .Y(_06156_));
 sky130_fd_sc_hd__a32o_1 _14672_ (.A1(net389),
    .A2(net493),
    .A3(_06020_),
    .B1(_06021_),
    .B2(net484),
    .X(_06157_));
 sky130_fd_sc_hd__a22o_1 _14673_ (.A1(net380),
    .A2(net497),
    .B1(net493),
    .B2(net385),
    .X(_06158_));
 sky130_fd_sc_hd__nand4_2 _14674_ (.A(net385),
    .B(net380),
    .C(net497),
    .D(net493),
    .Y(_06159_));
 sky130_fd_sc_hd__a22o_1 _14675_ (.A1(net372),
    .A2(net502),
    .B1(_06158_),
    .B2(_06159_),
    .X(_06160_));
 sky130_fd_sc_hd__nand4_2 _14676_ (.A(net372),
    .B(net502),
    .C(_06158_),
    .D(_06159_),
    .Y(_06161_));
 sky130_fd_sc_hd__nand3_1 _14677_ (.A(_06157_),
    .B(_06160_),
    .C(_06161_),
    .Y(_06162_));
 sky130_fd_sc_hd__a21o_1 _14678_ (.A1(_06160_),
    .A2(_06161_),
    .B1(_06157_),
    .X(_06163_));
 sky130_fd_sc_hd__nand3_1 _14679_ (.A(_06156_),
    .B(_06162_),
    .C(_06163_),
    .Y(_06164_));
 sky130_fd_sc_hd__a21o_1 _14680_ (.A1(_06162_),
    .A2(_06163_),
    .B1(_06156_),
    .X(_06165_));
 sky130_fd_sc_hd__a21bo_1 _14681_ (.A1(_05999_),
    .A2(_06006_),
    .B1_N(_06005_),
    .X(_06166_));
 sky130_fd_sc_hd__nand3_1 _14682_ (.A(_06164_),
    .B(_06165_),
    .C(_06166_),
    .Y(_06167_));
 sky130_fd_sc_hd__a21o_1 _14683_ (.A1(_06164_),
    .A2(_06165_),
    .B1(_06166_),
    .X(_06168_));
 sky130_fd_sc_hd__nand3_1 _14684_ (.A(_06155_),
    .B(_06167_),
    .C(_06168_),
    .Y(_06169_));
 sky130_fd_sc_hd__a21o_1 _14685_ (.A1(_06167_),
    .A2(_06168_),
    .B1(_06155_),
    .X(_06170_));
 sky130_fd_sc_hd__o211a_1 _14686_ (.A1(_06035_),
    .A2(_06037_),
    .B1(_06169_),
    .C1(_06170_),
    .X(_06171_));
 sky130_fd_sc_hd__a211oi_1 _14687_ (.A1(_06169_),
    .A2(_06170_),
    .B1(_06035_),
    .C1(_06037_),
    .Y(_06172_));
 sky130_fd_sc_hd__nor2_2 _14688_ (.A(_06171_),
    .B(_06172_),
    .Y(_06173_));
 sky130_fd_sc_hd__xor2_4 _14689_ (.A(_06140_),
    .B(_06173_),
    .X(_06174_));
 sky130_fd_sc_hd__nand2_2 _14690_ (.A(_06030_),
    .B(_06032_),
    .Y(_06175_));
 sky130_fd_sc_hd__a21o_1 _14691_ (.A1(_06040_),
    .A2(_06047_),
    .B1(_06046_),
    .X(_06176_));
 sky130_fd_sc_hd__a22o_1 _14692_ (.A1(net393),
    .A2(net484),
    .B1(net479),
    .B2(net398),
    .X(_06177_));
 sky130_fd_sc_hd__and3_1 _14693_ (.A(net398),
    .B(net393),
    .C(net484),
    .X(_06178_));
 sky130_fd_sc_hd__a21bo_1 _14694_ (.A1(net479),
    .A2(_06178_),
    .B1_N(_06177_),
    .X(_06179_));
 sky130_fd_sc_hd__nand2_1 _14695_ (.A(net388),
    .B(net488),
    .Y(_06180_));
 sky130_fd_sc_hd__xor2_1 _14696_ (.A(_06179_),
    .B(_06180_),
    .X(_06181_));
 sky130_fd_sc_hd__a22o_1 _14697_ (.A1(\mul0.b[10] ),
    .A2(net471),
    .B1(net469),
    .B2(net411),
    .X(_06182_));
 sky130_fd_sc_hd__nand4_2 _14698_ (.A(net412),
    .B(net407),
    .C(net471),
    .D(net469),
    .Y(_06183_));
 sky130_fd_sc_hd__inv_2 _14699_ (.A(_06183_),
    .Y(_06184_));
 sky130_fd_sc_hd__a22o_1 _14700_ (.A1(net402),
    .A2(net475),
    .B1(_06182_),
    .B2(_06183_),
    .X(_06185_));
 sky130_fd_sc_hd__and4_1 _14701_ (.A(net402),
    .B(net475),
    .C(_06182_),
    .D(_06183_),
    .X(_06186_));
 sky130_fd_sc_hd__nand4_2 _14702_ (.A(net402),
    .B(net475),
    .C(_06182_),
    .D(_06183_),
    .Y(_06187_));
 sky130_fd_sc_hd__o211ai_4 _14703_ (.A1(_06027_),
    .A2(_06029_),
    .B1(_06185_),
    .C1(_06187_),
    .Y(_06188_));
 sky130_fd_sc_hd__a211o_1 _14704_ (.A1(_06185_),
    .A2(_06187_),
    .B1(_06027_),
    .C1(_06029_),
    .X(_06189_));
 sky130_fd_sc_hd__nand3_2 _14705_ (.A(_06181_),
    .B(_06188_),
    .C(_06189_),
    .Y(_06190_));
 sky130_fd_sc_hd__a21o_1 _14706_ (.A1(_06188_),
    .A2(_06189_),
    .B1(_06181_),
    .X(_06191_));
 sky130_fd_sc_hd__and3_2 _14707_ (.A(_06176_),
    .B(_06190_),
    .C(_06191_),
    .X(_06192_));
 sky130_fd_sc_hd__a21oi_1 _14708_ (.A1(_06190_),
    .A2(_06191_),
    .B1(_06176_),
    .Y(_06193_));
 sky130_fd_sc_hd__or2_2 _14709_ (.A(_06192_),
    .B(_06193_),
    .X(_06194_));
 sky130_fd_sc_hd__a211oi_2 _14710_ (.A1(_06030_),
    .A2(_06032_),
    .B1(_06192_),
    .C1(_06193_),
    .Y(_06195_));
 sky130_fd_sc_hd__xnor2_4 _14711_ (.A(_06175_),
    .B(_06194_),
    .Y(_06196_));
 sky130_fd_sc_hd__and3_1 _14712_ (.A(net439),
    .B(net434),
    .C(net453),
    .X(_06197_));
 sky130_fd_sc_hd__nand3_2 _14713_ (.A(net438),
    .B(net433),
    .C(net453),
    .Y(_06198_));
 sky130_fd_sc_hd__o21a_2 _14714_ (.A1(net438),
    .A2(net433),
    .B1(net453),
    .X(_06199_));
 sky130_fd_sc_hd__a22o_1 _14715_ (.A1(net429),
    .A2(net456),
    .B1(_06198_),
    .B2(_06199_),
    .X(_06200_));
 sky130_fd_sc_hd__nand4_2 _14716_ (.A(net429),
    .B(net456),
    .C(_06198_),
    .D(_06199_),
    .Y(_06201_));
 sky130_fd_sc_hd__a211o_1 _14717_ (.A1(_06200_),
    .A2(_06201_),
    .B1(_05739_),
    .C1(_05904_),
    .X(_06202_));
 sky130_fd_sc_hd__o211a_1 _14718_ (.A1(_05739_),
    .A2(_05904_),
    .B1(_06200_),
    .C1(_06201_),
    .X(_06203_));
 sky130_fd_sc_hd__o211ai_2 _14719_ (.A1(_05739_),
    .A2(_05904_),
    .B1(_06200_),
    .C1(_06201_),
    .Y(_06204_));
 sky130_fd_sc_hd__a211oi_1 _14720_ (.A1(_06202_),
    .A2(_06204_),
    .B1(_06055_),
    .C1(_06058_),
    .Y(_06205_));
 sky130_fd_sc_hd__a211o_1 _14721_ (.A1(_06202_),
    .A2(_06204_),
    .B1(_06055_),
    .C1(_06058_),
    .X(_06206_));
 sky130_fd_sc_hd__o211a_1 _14722_ (.A1(_06055_),
    .A2(_06058_),
    .B1(_06202_),
    .C1(_06204_),
    .X(_06207_));
 sky130_fd_sc_hd__nor2_2 _14723_ (.A(_06205_),
    .B(_06207_),
    .Y(_06208_));
 sky130_fd_sc_hd__nand2_1 _14724_ (.A(_06043_),
    .B(_06045_),
    .Y(_06209_));
 sky130_fd_sc_hd__a21bo_1 _14725_ (.A1(_06050_),
    .A2(_06052_),
    .B1_N(_06051_),
    .X(_06210_));
 sky130_fd_sc_hd__a22o_1 _14726_ (.A1(net420),
    .A2(net461),
    .B1(net459),
    .B2(net423),
    .X(_06211_));
 sky130_fd_sc_hd__nand4_2 _14727_ (.A(net424),
    .B(net420),
    .C(net461),
    .D(net459),
    .Y(_06212_));
 sky130_fd_sc_hd__a22o_1 _14728_ (.A1(net415),
    .A2(net464),
    .B1(_06211_),
    .B2(_06212_),
    .X(_06213_));
 sky130_fd_sc_hd__nand4_2 _14729_ (.A(net416),
    .B(net464),
    .C(_06211_),
    .D(_06212_),
    .Y(_06214_));
 sky130_fd_sc_hd__nand3_1 _14730_ (.A(_06210_),
    .B(_06213_),
    .C(_06214_),
    .Y(_06215_));
 sky130_fd_sc_hd__a21o_1 _14731_ (.A1(_06213_),
    .A2(_06214_),
    .B1(_06210_),
    .X(_06216_));
 sky130_fd_sc_hd__nand3_1 _14732_ (.A(_06209_),
    .B(_06215_),
    .C(_06216_),
    .Y(_06217_));
 sky130_fd_sc_hd__a21o_1 _14733_ (.A1(_06215_),
    .A2(_06216_),
    .B1(_06209_),
    .X(_06218_));
 sky130_fd_sc_hd__and2_2 _14734_ (.A(_06217_),
    .B(_06218_),
    .X(_06219_));
 sky130_fd_sc_hd__xnor2_4 _14735_ (.A(_06208_),
    .B(_06219_),
    .Y(_06220_));
 sky130_fd_sc_hd__a21oi_4 _14736_ (.A1(_06049_),
    .A2(_06061_),
    .B1(_06060_),
    .Y(_06221_));
 sky130_fd_sc_hd__nor2_1 _14737_ (.A(_06220_),
    .B(_06221_),
    .Y(_06222_));
 sky130_fd_sc_hd__xor2_4 _14738_ (.A(_06220_),
    .B(_06221_),
    .X(_06223_));
 sky130_fd_sc_hd__xor2_4 _14739_ (.A(_06196_),
    .B(_06223_),
    .X(_06224_));
 sky130_fd_sc_hd__a21oi_4 _14740_ (.A1(_06039_),
    .A2(_06065_),
    .B1(_06064_),
    .Y(_06225_));
 sky130_fd_sc_hd__and2b_1 _14741_ (.A_N(_06225_),
    .B(_06224_),
    .X(_06226_));
 sky130_fd_sc_hd__xnor2_4 _14742_ (.A(_06224_),
    .B(_06225_),
    .Y(_06227_));
 sky130_fd_sc_hd__xnor2_4 _14743_ (.A(_06174_),
    .B(_06227_),
    .Y(_06228_));
 sky130_fd_sc_hd__a21boi_4 _14744_ (.A1(_06017_),
    .A2(_06069_),
    .B1_N(_06068_),
    .Y(_06229_));
 sky130_fd_sc_hd__nor2_1 _14745_ (.A(_06228_),
    .B(_06229_),
    .Y(_06230_));
 sky130_fd_sc_hd__xor2_4 _14746_ (.A(_06228_),
    .B(_06229_),
    .X(_06231_));
 sky130_fd_sc_hd__xor2_4 _14747_ (.A(_06139_),
    .B(_06231_),
    .X(_06232_));
 sky130_fd_sc_hd__a21oi_4 _14748_ (.A1(_05982_),
    .A2(_06073_),
    .B1(_06072_),
    .Y(_06233_));
 sky130_fd_sc_hd__nand2b_1 _14749_ (.A_N(_06233_),
    .B(_06232_),
    .Y(_06234_));
 sky130_fd_sc_hd__xnor2_4 _14750_ (.A(_06232_),
    .B(_06233_),
    .Y(_06235_));
 sky130_fd_sc_hd__xnor2_4 _14751_ (.A(_06096_),
    .B(_06235_),
    .Y(_06236_));
 sky130_fd_sc_hd__a21boi_4 _14752_ (.A1(_05939_),
    .A2(_06077_),
    .B1_N(_06076_),
    .Y(_06237_));
 sky130_fd_sc_hd__nor2_1 _14753_ (.A(_06236_),
    .B(_06237_),
    .Y(_06238_));
 sky130_fd_sc_hd__xor2_4 _14754_ (.A(_06236_),
    .B(_06237_),
    .X(_06239_));
 sky130_fd_sc_hd__xnor2_4 _14755_ (.A(_06095_),
    .B(_06239_),
    .Y(_06240_));
 sky130_fd_sc_hd__nor2_1 _14756_ (.A(_06094_),
    .B(_06240_),
    .Y(_06241_));
 sky130_fd_sc_hd__nand2_1 _14757_ (.A(_06094_),
    .B(_06240_),
    .Y(_06242_));
 sky130_fd_sc_hd__xor2_4 _14758_ (.A(_06094_),
    .B(_06240_),
    .X(_06243_));
 sky130_fd_sc_hd__xnor2_4 _14759_ (.A(_06093_),
    .B(_06243_),
    .Y(_06244_));
 sky130_fd_sc_hd__nor2_1 _14760_ (.A(net9),
    .B(_06244_),
    .Y(_06245_));
 sky130_fd_sc_hd__a221o_1 _14761_ (.A1(\state[4] ),
    .A2(\temp[18] ),
    .B1(_02663_),
    .B2(net6),
    .C1(_06245_),
    .X(_06246_));
 sky130_fd_sc_hd__mux2_1 _14762_ (.A0(net729),
    .A1(_06246_),
    .S(_03055_),
    .X(_00285_));
 sky130_fd_sc_hd__a21o_1 _14763_ (.A1(_06110_),
    .A2(_06111_),
    .B1(_06113_),
    .X(_06247_));
 sky130_fd_sc_hd__or2_1 _14764_ (.A(_06136_),
    .B(_06138_),
    .X(_06248_));
 sky130_fd_sc_hd__o21ba_1 _14765_ (.A1(_06115_),
    .A2(_06134_),
    .B1_N(_06133_),
    .X(_06249_));
 sky130_fd_sc_hd__a21oi_2 _14766_ (.A1(_06140_),
    .A2(_06173_),
    .B1(_06171_),
    .Y(_06250_));
 sky130_fd_sc_hd__a22o_1 _14767_ (.A1(net543),
    .A2(net334),
    .B1(net331),
    .B2(net547),
    .X(_06251_));
 sky130_fd_sc_hd__nand4_2 _14768_ (.A(net543),
    .B(net547),
    .C(net334),
    .D(net331),
    .Y(_06252_));
 sky130_fd_sc_hd__nand2_1 _14769_ (.A(_06251_),
    .B(_06252_),
    .Y(_06253_));
 sky130_fd_sc_hd__nand2_1 _14770_ (.A(net551),
    .B(net329),
    .Y(_06254_));
 sky130_fd_sc_hd__xnor2_2 _14771_ (.A(_06253_),
    .B(_06254_),
    .Y(_06255_));
 sky130_fd_sc_hd__o2bb2a_2 _14772_ (.A1_N(net334),
    .A2_N(_06100_),
    .B1(_06101_),
    .B2(_06102_),
    .X(_06256_));
 sky130_fd_sc_hd__xnor2_2 _14773_ (.A(_06255_),
    .B(_06256_),
    .Y(_06257_));
 sky130_fd_sc_hd__and4b_2 _14774_ (.A_N(net560),
    .B(net327),
    .C(net326),
    .D(net556),
    .X(_06258_));
 sky130_fd_sc_hd__inv_2 _14775_ (.A(_06258_),
    .Y(_06259_));
 sky130_fd_sc_hd__o2bb2a_1 _14776_ (.A1_N(net556),
    .A2_N(net327),
    .B1(net57),
    .B2(net560),
    .X(_06260_));
 sky130_fd_sc_hd__nor2_1 _14777_ (.A(_06258_),
    .B(_06260_),
    .Y(_06261_));
 sky130_fd_sc_hd__xnor2_1 _14778_ (.A(_06257_),
    .B(_06261_),
    .Y(_06262_));
 sky130_fd_sc_hd__o32ai_4 _14779_ (.A1(_06105_),
    .A2(_06106_),
    .A3(_06108_),
    .B1(_06104_),
    .B2(_06103_),
    .Y(_06263_));
 sky130_fd_sc_hd__xnor2_1 _14780_ (.A(_06262_),
    .B(_06263_),
    .Y(_06264_));
 sky130_fd_sc_hd__nor2_1 _14781_ (.A(_06107_),
    .B(_06264_),
    .Y(_06265_));
 sky130_fd_sc_hd__and2_1 _14782_ (.A(_06107_),
    .B(_06264_),
    .X(_06266_));
 sky130_fd_sc_hd__or2_1 _14783_ (.A(_06265_),
    .B(_06266_),
    .X(_06267_));
 sky130_fd_sc_hd__a21oi_1 _14784_ (.A1(_06145_),
    .A2(_06153_),
    .B1(_06152_),
    .Y(_06268_));
 sky130_fd_sc_hd__nand2_1 _14785_ (.A(_06120_),
    .B(_06122_),
    .Y(_06269_));
 sky130_fd_sc_hd__a32o_1 _14786_ (.A1(net528),
    .A2(net349),
    .A3(_06141_),
    .B1(_06142_),
    .B2(net357),
    .X(_06270_));
 sky130_fd_sc_hd__a22o_1 _14787_ (.A1(net528),
    .A2(net346),
    .B1(net342),
    .B2(net534),
    .X(_06271_));
 sky130_fd_sc_hd__nand4_2 _14788_ (.A(net528),
    .B(net534),
    .C(net346),
    .D(net342),
    .Y(_06272_));
 sky130_fd_sc_hd__a22o_1 _14789_ (.A1(net538),
    .A2(net338),
    .B1(_06271_),
    .B2(_06272_),
    .X(_06273_));
 sky130_fd_sc_hd__nand4_2 _14790_ (.A(net538),
    .B(net338),
    .C(_06271_),
    .D(_06272_),
    .Y(_06274_));
 sky130_fd_sc_hd__nand3_2 _14791_ (.A(_06270_),
    .B(_06273_),
    .C(_06274_),
    .Y(_06275_));
 sky130_fd_sc_hd__a21o_1 _14792_ (.A1(_06273_),
    .A2(_06274_),
    .B1(_06270_),
    .X(_06276_));
 sky130_fd_sc_hd__nand3_2 _14793_ (.A(_06269_),
    .B(_06275_),
    .C(_06276_),
    .Y(_06277_));
 sky130_fd_sc_hd__a21o_1 _14794_ (.A1(_06275_),
    .A2(_06276_),
    .B1(_06269_),
    .X(_06278_));
 sky130_fd_sc_hd__and3b_1 _14795_ (.A_N(_06268_),
    .B(_06277_),
    .C(_06278_),
    .X(_06279_));
 sky130_fd_sc_hd__a21boi_1 _14796_ (.A1(_06277_),
    .A2(_06278_),
    .B1_N(_06268_),
    .Y(_06280_));
 sky130_fd_sc_hd__a211oi_2 _14797_ (.A1(_06123_),
    .A2(_06125_),
    .B1(_06279_),
    .C1(_06280_),
    .Y(_06281_));
 sky130_fd_sc_hd__o211ai_1 _14798_ (.A1(_06279_),
    .A2(_06280_),
    .B1(_06123_),
    .C1(_06125_),
    .Y(_06282_));
 sky130_fd_sc_hd__and2b_1 _14799_ (.A_N(_06281_),
    .B(_06282_),
    .X(_06283_));
 sky130_fd_sc_hd__nor2_1 _14800_ (.A(_06127_),
    .B(_06129_),
    .Y(_06284_));
 sky130_fd_sc_hd__and2b_1 _14801_ (.A_N(_06284_),
    .B(_06283_),
    .X(_06285_));
 sky130_fd_sc_hd__xnor2_1 _14802_ (.A(_06283_),
    .B(_06284_),
    .Y(_06286_));
 sky130_fd_sc_hd__and2b_1 _14803_ (.A_N(_06267_),
    .B(_06286_),
    .X(_06287_));
 sky130_fd_sc_hd__xnor2_1 _14804_ (.A(_06267_),
    .B(_06286_),
    .Y(_06288_));
 sky130_fd_sc_hd__and2b_1 _14805_ (.A_N(_06250_),
    .B(_06288_),
    .X(_06289_));
 sky130_fd_sc_hd__xnor2_1 _14806_ (.A(_06250_),
    .B(_06288_),
    .Y(_06290_));
 sky130_fd_sc_hd__and2b_1 _14807_ (.A_N(_06249_),
    .B(_06290_),
    .X(_06291_));
 sky130_fd_sc_hd__xnor2_1 _14808_ (.A(_06249_),
    .B(_06290_),
    .Y(_06292_));
 sky130_fd_sc_hd__nand2_1 _14809_ (.A(_06167_),
    .B(_06169_),
    .Y(_06293_));
 sky130_fd_sc_hd__a22o_1 _14810_ (.A1(net513),
    .A2(net357),
    .B1(net352),
    .B2(net518),
    .X(_06294_));
 sky130_fd_sc_hd__and3_1 _14811_ (.A(net513),
    .B(net518),
    .C(net352),
    .X(_06295_));
 sky130_fd_sc_hd__a21bo_1 _14812_ (.A1(net357),
    .A2(_06295_),
    .B1_N(_06294_),
    .X(_06296_));
 sky130_fd_sc_hd__nand2_1 _14813_ (.A(net523),
    .B(net349),
    .Y(_06297_));
 sky130_fd_sc_hd__xor2_2 _14814_ (.A(_06296_),
    .B(_06297_),
    .X(_06298_));
 sky130_fd_sc_hd__a22o_1 _14815_ (.A1(net500),
    .A2(net634),
    .B1(net366),
    .B2(net506),
    .X(_06299_));
 sky130_fd_sc_hd__and4_1 _14816_ (.A(net505),
    .B(net501),
    .C(net634),
    .D(net366),
    .X(_06300_));
 sky130_fd_sc_hd__nand4_1 _14817_ (.A(net506),
    .B(net500),
    .C(net633),
    .D(net366),
    .Y(_06301_));
 sky130_fd_sc_hd__a22o_1 _14818_ (.A1(net510),
    .A2(net361),
    .B1(_06299_),
    .B2(_06301_),
    .X(_06302_));
 sky130_fd_sc_hd__and4_1 _14819_ (.A(net510),
    .B(net361),
    .C(_06299_),
    .D(_06301_),
    .X(_06303_));
 sky130_fd_sc_hd__nand4_1 _14820_ (.A(net510),
    .B(net361),
    .C(_06299_),
    .D(_06301_),
    .Y(_06304_));
 sky130_fd_sc_hd__o211a_1 _14821_ (.A1(_06147_),
    .A2(_06150_),
    .B1(_06302_),
    .C1(_06304_),
    .X(_06305_));
 sky130_fd_sc_hd__a211o_1 _14822_ (.A1(_06302_),
    .A2(_06304_),
    .B1(_06147_),
    .C1(_06150_),
    .X(_06306_));
 sky130_fd_sc_hd__nand2b_1 _14823_ (.A_N(_06305_),
    .B(_06306_),
    .Y(_06307_));
 sky130_fd_sc_hd__xnor2_2 _14824_ (.A(_06298_),
    .B(_06307_),
    .Y(_06308_));
 sky130_fd_sc_hd__nand2_1 _14825_ (.A(_06159_),
    .B(_06161_),
    .Y(_06309_));
 sky130_fd_sc_hd__a32o_1 _14826_ (.A1(net388),
    .A2(net488),
    .A3(_06177_),
    .B1(_06178_),
    .B2(net479),
    .X(_06310_));
 sky130_fd_sc_hd__a22o_1 _14827_ (.A1(net378),
    .A2(net493),
    .B1(net488),
    .B2(net384),
    .X(_06311_));
 sky130_fd_sc_hd__nand4_2 _14828_ (.A(net385),
    .B(net380),
    .C(net493),
    .D(net488),
    .Y(_06312_));
 sky130_fd_sc_hd__a22o_1 _14829_ (.A1(net372),
    .A2(net497),
    .B1(_06311_),
    .B2(_06312_),
    .X(_06313_));
 sky130_fd_sc_hd__nand4_2 _14830_ (.A(net372),
    .B(net497),
    .C(_06311_),
    .D(_06312_),
    .Y(_06314_));
 sky130_fd_sc_hd__nand3_1 _14831_ (.A(_06310_),
    .B(_06313_),
    .C(_06314_),
    .Y(_06315_));
 sky130_fd_sc_hd__a21o_1 _14832_ (.A1(_06313_),
    .A2(_06314_),
    .B1(_06310_),
    .X(_06316_));
 sky130_fd_sc_hd__nand3_1 _14833_ (.A(_06309_),
    .B(_06315_),
    .C(_06316_),
    .Y(_06317_));
 sky130_fd_sc_hd__a21o_1 _14834_ (.A1(_06315_),
    .A2(_06316_),
    .B1(_06309_),
    .X(_06318_));
 sky130_fd_sc_hd__a21bo_1 _14835_ (.A1(_06156_),
    .A2(_06163_),
    .B1_N(_06162_),
    .X(_06319_));
 sky130_fd_sc_hd__nand3_2 _14836_ (.A(_06317_),
    .B(_06318_),
    .C(_06319_),
    .Y(_06320_));
 sky130_fd_sc_hd__inv_2 _14837_ (.A(_06320_),
    .Y(_06321_));
 sky130_fd_sc_hd__a21o_1 _14838_ (.A1(_06317_),
    .A2(_06318_),
    .B1(_06319_),
    .X(_06322_));
 sky130_fd_sc_hd__and3_1 _14839_ (.A(_06308_),
    .B(_06320_),
    .C(_06322_),
    .X(_06323_));
 sky130_fd_sc_hd__nand3_1 _14840_ (.A(_06308_),
    .B(_06320_),
    .C(_06322_),
    .Y(_06324_));
 sky130_fd_sc_hd__a21o_1 _14841_ (.A1(_06320_),
    .A2(_06322_),
    .B1(_06308_),
    .X(_06325_));
 sky130_fd_sc_hd__o211ai_2 _14842_ (.A1(_06192_),
    .A2(_06195_),
    .B1(_06324_),
    .C1(_06325_),
    .Y(_06326_));
 sky130_fd_sc_hd__a211o_1 _14843_ (.A1(_06324_),
    .A2(_06325_),
    .B1(_06192_),
    .C1(_06195_),
    .X(_06327_));
 sky130_fd_sc_hd__and3_1 _14844_ (.A(_06293_),
    .B(_06326_),
    .C(_06327_),
    .X(_06328_));
 sky130_fd_sc_hd__a21oi_1 _14845_ (.A1(_06326_),
    .A2(_06327_),
    .B1(_06293_),
    .Y(_06329_));
 sky130_fd_sc_hd__nor2_1 _14846_ (.A(_06328_),
    .B(_06329_),
    .Y(_06330_));
 sky130_fd_sc_hd__a22o_1 _14847_ (.A1(net428),
    .A2(net453),
    .B1(_06198_),
    .B2(_06199_),
    .X(_06331_));
 sky130_fd_sc_hd__nand3_1 _14848_ (.A(net428),
    .B(_06198_),
    .C(_06199_),
    .Y(_06332_));
 sky130_fd_sc_hd__a211o_2 _14849_ (.A1(_06331_),
    .A2(_06332_),
    .B1(_05739_),
    .C1(_05904_),
    .X(_06333_));
 sky130_fd_sc_hd__o211ai_2 _14850_ (.A1(_05739_),
    .A2(_05904_),
    .B1(_06331_),
    .C1(_06332_),
    .Y(_06334_));
 sky130_fd_sc_hd__o211a_1 _14851_ (.A1(_06058_),
    .A2(_06203_),
    .B1(_06333_),
    .C1(_06334_),
    .X(_06335_));
 sky130_fd_sc_hd__o211ai_1 _14852_ (.A1(_06058_),
    .A2(_06203_),
    .B1(_06333_),
    .C1(_06334_),
    .Y(_06336_));
 sky130_fd_sc_hd__a211o_1 _14853_ (.A1(_06333_),
    .A2(_06334_),
    .B1(_06058_),
    .C1(_06203_),
    .X(_06337_));
 sky130_fd_sc_hd__nand2_1 _14854_ (.A(_06212_),
    .B(_06214_),
    .Y(_06338_));
 sky130_fd_sc_hd__a31o_1 _14855_ (.A1(net429),
    .A2(net456),
    .A3(_06199_),
    .B1(_06197_),
    .X(_06339_));
 sky130_fd_sc_hd__a22o_1 _14856_ (.A1(net419),
    .A2(\mul0.a[29] ),
    .B1(net456),
    .B2(net425),
    .X(_06340_));
 sky130_fd_sc_hd__nand4_2 _14857_ (.A(net424),
    .B(\mul0.b[7] ),
    .C(\mul0.a[29] ),
    .D(net456),
    .Y(_06341_));
 sky130_fd_sc_hd__a22o_1 _14858_ (.A1(net415),
    .A2(net461),
    .B1(_06340_),
    .B2(_06341_),
    .X(_06342_));
 sky130_fd_sc_hd__nand4_1 _14859_ (.A(net415),
    .B(net461),
    .C(_06340_),
    .D(_06341_),
    .Y(_06343_));
 sky130_fd_sc_hd__nand3_1 _14860_ (.A(_06339_),
    .B(_06342_),
    .C(_06343_),
    .Y(_06344_));
 sky130_fd_sc_hd__a21o_1 _14861_ (.A1(_06342_),
    .A2(_06343_),
    .B1(_06339_),
    .X(_06345_));
 sky130_fd_sc_hd__nand3_1 _14862_ (.A(_06338_),
    .B(_06344_),
    .C(_06345_),
    .Y(_06346_));
 sky130_fd_sc_hd__a21o_1 _14863_ (.A1(_06344_),
    .A2(_06345_),
    .B1(_06338_),
    .X(_06347_));
 sky130_fd_sc_hd__a22o_1 _14864_ (.A1(_06336_),
    .A2(_06337_),
    .B1(_06346_),
    .B2(_06347_),
    .X(_06348_));
 sky130_fd_sc_hd__nand4_1 _14865_ (.A(_06336_),
    .B(_06337_),
    .C(_06346_),
    .D(_06347_),
    .Y(_06349_));
 sky130_fd_sc_hd__a31o_1 _14866_ (.A1(_06206_),
    .A2(_06217_),
    .A3(_06218_),
    .B1(_06207_),
    .X(_06350_));
 sky130_fd_sc_hd__a21oi_2 _14867_ (.A1(_06348_),
    .A2(_06349_),
    .B1(_06350_),
    .Y(_06351_));
 sky130_fd_sc_hd__and3_1 _14868_ (.A(_06348_),
    .B(_06349_),
    .C(_06350_),
    .X(_06352_));
 sky130_fd_sc_hd__a21bo_1 _14869_ (.A1(_06209_),
    .A2(_06216_),
    .B1_N(_06215_),
    .X(_06353_));
 sky130_fd_sc_hd__a22o_1 _14870_ (.A1(net393),
    .A2(net481),
    .B1(net475),
    .B2(net399),
    .X(_06354_));
 sky130_fd_sc_hd__and3_1 _14871_ (.A(net399),
    .B(net393),
    .C(net479),
    .X(_06355_));
 sky130_fd_sc_hd__a21bo_1 _14872_ (.A1(net477),
    .A2(_06355_),
    .B1_N(_06354_),
    .X(_06356_));
 sky130_fd_sc_hd__nand2_1 _14873_ (.A(net388),
    .B(net483),
    .Y(_06357_));
 sky130_fd_sc_hd__xor2_1 _14874_ (.A(_06356_),
    .B(_06357_),
    .X(_06358_));
 sky130_fd_sc_hd__a22o_1 _14875_ (.A1(net407),
    .A2(net468),
    .B1(net465),
    .B2(net411),
    .X(_06359_));
 sky130_fd_sc_hd__nand4_4 _14876_ (.A(net411),
    .B(net407),
    .C(net468),
    .D(net465),
    .Y(_06360_));
 sky130_fd_sc_hd__a22o_1 _14877_ (.A1(\mul0.b[11] ),
    .A2(net471),
    .B1(_06359_),
    .B2(_06360_),
    .X(_06361_));
 sky130_fd_sc_hd__nand4_4 _14878_ (.A(\mul0.b[11] ),
    .B(net471),
    .C(_06359_),
    .D(_06360_),
    .Y(_06362_));
 sky130_fd_sc_hd__o211ai_4 _14879_ (.A1(_06184_),
    .A2(_06186_),
    .B1(_06361_),
    .C1(_06362_),
    .Y(_06363_));
 sky130_fd_sc_hd__a211o_1 _14880_ (.A1(_06361_),
    .A2(_06362_),
    .B1(_06184_),
    .C1(_06186_),
    .X(_06364_));
 sky130_fd_sc_hd__nand3_2 _14881_ (.A(_06358_),
    .B(_06363_),
    .C(_06364_),
    .Y(_06365_));
 sky130_fd_sc_hd__a21o_1 _14882_ (.A1(_06363_),
    .A2(_06364_),
    .B1(_06358_),
    .X(_06366_));
 sky130_fd_sc_hd__and3_2 _14883_ (.A(_06353_),
    .B(_06365_),
    .C(_06366_),
    .X(_06367_));
 sky130_fd_sc_hd__a21oi_2 _14884_ (.A1(_06365_),
    .A2(_06366_),
    .B1(_06353_),
    .Y(_06368_));
 sky130_fd_sc_hd__a211oi_4 _14885_ (.A1(_06188_),
    .A2(_06190_),
    .B1(_06367_),
    .C1(_06368_),
    .Y(_06369_));
 sky130_fd_sc_hd__o211a_1 _14886_ (.A1(_06367_),
    .A2(_06368_),
    .B1(_06188_),
    .C1(_06190_),
    .X(_06370_));
 sky130_fd_sc_hd__nor4_2 _14887_ (.A(_06351_),
    .B(_06352_),
    .C(_06369_),
    .D(_06370_),
    .Y(_06371_));
 sky130_fd_sc_hd__o22a_1 _14888_ (.A1(_06351_),
    .A2(_06352_),
    .B1(_06369_),
    .B2(_06370_),
    .X(_06372_));
 sky130_fd_sc_hd__nor2_2 _14889_ (.A(_06371_),
    .B(_06372_),
    .Y(_06373_));
 sky130_fd_sc_hd__a21oi_2 _14890_ (.A1(_06196_),
    .A2(_06223_),
    .B1(_06222_),
    .Y(_06374_));
 sky130_fd_sc_hd__and2b_1 _14891_ (.A_N(_06374_),
    .B(_06373_),
    .X(_06375_));
 sky130_fd_sc_hd__xnor2_2 _14892_ (.A(_06373_),
    .B(_06374_),
    .Y(_06376_));
 sky130_fd_sc_hd__xnor2_2 _14893_ (.A(_06330_),
    .B(_06376_),
    .Y(_06377_));
 sky130_fd_sc_hd__a21oi_2 _14894_ (.A1(_06174_),
    .A2(_06227_),
    .B1(_06226_),
    .Y(_06378_));
 sky130_fd_sc_hd__nor2_1 _14895_ (.A(_06377_),
    .B(_06378_),
    .Y(_06379_));
 sky130_fd_sc_hd__xor2_2 _14896_ (.A(_06377_),
    .B(_06378_),
    .X(_06380_));
 sky130_fd_sc_hd__xor2_1 _14897_ (.A(_06292_),
    .B(_06380_),
    .X(_06381_));
 sky130_fd_sc_hd__a21oi_2 _14898_ (.A1(_06139_),
    .A2(_06231_),
    .B1(_06230_),
    .Y(_06382_));
 sky130_fd_sc_hd__nand2b_1 _14899_ (.A_N(_06382_),
    .B(_06381_),
    .Y(_06383_));
 sky130_fd_sc_hd__xnor2_1 _14900_ (.A(_06381_),
    .B(_06382_),
    .Y(_06384_));
 sky130_fd_sc_hd__xnor2_1 _14901_ (.A(_06248_),
    .B(_06384_),
    .Y(_06385_));
 sky130_fd_sc_hd__a21boi_2 _14902_ (.A1(_06096_),
    .A2(_06235_),
    .B1_N(_06234_),
    .Y(_06386_));
 sky130_fd_sc_hd__or2_1 _14903_ (.A(_06385_),
    .B(_06386_),
    .X(_06387_));
 sky130_fd_sc_hd__xor2_1 _14904_ (.A(_06385_),
    .B(_06386_),
    .X(_06388_));
 sky130_fd_sc_hd__nand2_1 _14905_ (.A(_06247_),
    .B(_06388_),
    .Y(_06389_));
 sky130_fd_sc_hd__xnor2_1 _14906_ (.A(_06247_),
    .B(_06388_),
    .Y(_06390_));
 sky130_fd_sc_hd__a21oi_1 _14907_ (.A1(_06095_),
    .A2(_06239_),
    .B1(_06238_),
    .Y(_06391_));
 sky130_fd_sc_hd__nor2_1 _14908_ (.A(_06390_),
    .B(_06391_),
    .Y(_06392_));
 sky130_fd_sc_hd__and2_1 _14909_ (.A(_06390_),
    .B(_06391_),
    .X(_06393_));
 sky130_fd_sc_hd__nor2_2 _14910_ (.A(_06392_),
    .B(_06393_),
    .Y(_06394_));
 sky130_fd_sc_hd__nand2_1 _14911_ (.A(_06085_),
    .B(_06243_),
    .Y(_06395_));
 sky130_fd_sc_hd__inv_2 _14912_ (.A(_06395_),
    .Y(_06396_));
 sky130_fd_sc_hd__or4b_1 _14913_ (.A(_05777_),
    .B(_06395_),
    .C(_05933_),
    .D_N(_05931_),
    .X(_06397_));
 sky130_fd_sc_hd__a31o_1 _14914_ (.A1(_05780_),
    .A2(_05781_),
    .A3(_05782_),
    .B1(_06397_),
    .X(_06398_));
 sky130_fd_sc_hd__a221oi_4 _14915_ (.A1(_06084_),
    .A2(_06242_),
    .B1(_06396_),
    .B2(_06086_),
    .C1(_06241_),
    .Y(_06399_));
 sky130_fd_sc_hd__and2_2 _14916_ (.A(_06398_),
    .B(_06399_),
    .X(_06400_));
 sky130_fd_sc_hd__nand2b_1 _14917_ (.A_N(_06400_),
    .B(_06394_),
    .Y(_06401_));
 sky130_fd_sc_hd__xnor2_4 _14918_ (.A(_06394_),
    .B(_06400_),
    .Y(_06402_));
 sky130_fd_sc_hd__a22o_1 _14919_ (.A1(\state[4] ),
    .A2(\temp[19] ),
    .B1(_02671_),
    .B2(net5),
    .X(_06403_));
 sky130_fd_sc_hd__a21o_1 _14920_ (.A1(_03058_),
    .A2(_06402_),
    .B1(_06403_),
    .X(_06404_));
 sky130_fd_sc_hd__mux2_1 _14921_ (.A0(net748),
    .A1(_06404_),
    .S(net4),
    .X(_00286_));
 sky130_fd_sc_hd__nand2b_2 _14922_ (.A_N(_06392_),
    .B(_06401_),
    .Y(_06405_));
 sky130_fd_sc_hd__a21o_1 _14923_ (.A1(_06262_),
    .A2(_06263_),
    .B1(_06265_),
    .X(_06406_));
 sky130_fd_sc_hd__or2_1 _14924_ (.A(_06289_),
    .B(_06291_),
    .X(_06407_));
 sky130_fd_sc_hd__nor2_1 _14925_ (.A(_06285_),
    .B(_06287_),
    .Y(_06408_));
 sky130_fd_sc_hd__a21bo_1 _14926_ (.A1(_06293_),
    .A2(_06327_),
    .B1_N(_06326_),
    .X(_06409_));
 sky130_fd_sc_hd__a22o_1 _14927_ (.A1(net538),
    .A2(net334),
    .B1(net331),
    .B2(net543),
    .X(_06410_));
 sky130_fd_sc_hd__nand4_2 _14928_ (.A(net538),
    .B(net543),
    .C(net334),
    .D(net331),
    .Y(_06411_));
 sky130_fd_sc_hd__a22o_1 _14929_ (.A1(net547),
    .A2(net329),
    .B1(_06410_),
    .B2(_06411_),
    .X(_06412_));
 sky130_fd_sc_hd__nand4_2 _14930_ (.A(net547),
    .B(net329),
    .C(_06410_),
    .D(_06411_),
    .Y(_06413_));
 sky130_fd_sc_hd__o21ai_2 _14931_ (.A1(_06253_),
    .A2(_06254_),
    .B1(_06252_),
    .Y(_06414_));
 sky130_fd_sc_hd__a21oi_1 _14932_ (.A1(_06412_),
    .A2(_06413_),
    .B1(_06414_),
    .Y(_06415_));
 sky130_fd_sc_hd__a21o_1 _14933_ (.A1(_06412_),
    .A2(_06413_),
    .B1(_06414_),
    .X(_06416_));
 sky130_fd_sc_hd__and3_1 _14934_ (.A(_06412_),
    .B(_06413_),
    .C(_06414_),
    .X(_06417_));
 sky130_fd_sc_hd__or2_1 _14935_ (.A(_06415_),
    .B(_06417_),
    .X(_06418_));
 sky130_fd_sc_hd__and4b_1 _14936_ (.A_N(net556),
    .B(net327),
    .C(net326),
    .D(net551),
    .X(_06419_));
 sky130_fd_sc_hd__inv_2 _14937_ (.A(_06419_),
    .Y(_06420_));
 sky130_fd_sc_hd__o2bb2a_1 _14938_ (.A1_N(\mul0.a[7] ),
    .A2_N(net327),
    .B1(net57),
    .B2(net556),
    .X(_06421_));
 sky130_fd_sc_hd__nor2_1 _14939_ (.A(_06419_),
    .B(_06421_),
    .Y(_06422_));
 sky130_fd_sc_hd__xnor2_2 _14940_ (.A(_06418_),
    .B(_06422_),
    .Y(_06423_));
 sky130_fd_sc_hd__o32ai_4 _14941_ (.A1(_06257_),
    .A2(_06258_),
    .A3(_06260_),
    .B1(_06256_),
    .B2(_06255_),
    .Y(_06424_));
 sky130_fd_sc_hd__xnor2_2 _14942_ (.A(_06423_),
    .B(_06424_),
    .Y(_06425_));
 sky130_fd_sc_hd__nor2_1 _14943_ (.A(_06259_),
    .B(_06425_),
    .Y(_06426_));
 sky130_fd_sc_hd__xnor2_2 _14944_ (.A(_06259_),
    .B(_06425_),
    .Y(_06427_));
 sky130_fd_sc_hd__a21o_1 _14945_ (.A1(_06298_),
    .A2(_06306_),
    .B1(_06305_),
    .X(_06428_));
 sky130_fd_sc_hd__nand2_1 _14946_ (.A(_06272_),
    .B(_06274_),
    .Y(_06429_));
 sky130_fd_sc_hd__a32o_1 _14947_ (.A1(net522),
    .A2(net349),
    .A3(_06294_),
    .B1(_06295_),
    .B2(net357),
    .X(_06430_));
 sky130_fd_sc_hd__a22o_1 _14948_ (.A1(net522),
    .A2(net346),
    .B1(net342),
    .B2(net528),
    .X(_06431_));
 sky130_fd_sc_hd__nand4_2 _14949_ (.A(net522),
    .B(net528),
    .C(net346),
    .D(net342),
    .Y(_06432_));
 sky130_fd_sc_hd__a22o_1 _14950_ (.A1(net534),
    .A2(net339),
    .B1(_06431_),
    .B2(_06432_),
    .X(_06433_));
 sky130_fd_sc_hd__nand4_2 _14951_ (.A(net534),
    .B(net339),
    .C(_06431_),
    .D(_06432_),
    .Y(_06434_));
 sky130_fd_sc_hd__nand3_2 _14952_ (.A(_06430_),
    .B(_06433_),
    .C(_06434_),
    .Y(_06435_));
 sky130_fd_sc_hd__a21o_1 _14953_ (.A1(_06433_),
    .A2(_06434_),
    .B1(_06430_),
    .X(_06436_));
 sky130_fd_sc_hd__nand3_2 _14954_ (.A(_06429_),
    .B(_06435_),
    .C(_06436_),
    .Y(_06437_));
 sky130_fd_sc_hd__a21o_1 _14955_ (.A1(_06435_),
    .A2(_06436_),
    .B1(_06429_),
    .X(_06438_));
 sky130_fd_sc_hd__and3_2 _14956_ (.A(_06428_),
    .B(_06437_),
    .C(_06438_),
    .X(_06439_));
 sky130_fd_sc_hd__a21oi_2 _14957_ (.A1(_06437_),
    .A2(_06438_),
    .B1(_06428_),
    .Y(_06440_));
 sky130_fd_sc_hd__a211oi_1 _14958_ (.A1(_06275_),
    .A2(_06277_),
    .B1(_06439_),
    .C1(_06440_),
    .Y(_06441_));
 sky130_fd_sc_hd__a211o_1 _14959_ (.A1(_06275_),
    .A2(_06277_),
    .B1(_06439_),
    .C1(_06440_),
    .X(_06442_));
 sky130_fd_sc_hd__o211ai_2 _14960_ (.A1(_06439_),
    .A2(_06440_),
    .B1(_06275_),
    .C1(_06277_),
    .Y(_06443_));
 sky130_fd_sc_hd__o211a_1 _14961_ (.A1(_06279_),
    .A2(_06281_),
    .B1(_06442_),
    .C1(_06443_),
    .X(_06444_));
 sky130_fd_sc_hd__inv_2 _14962_ (.A(_06444_),
    .Y(_06445_));
 sky130_fd_sc_hd__a211oi_1 _14963_ (.A1(_06442_),
    .A2(_06443_),
    .B1(_06279_),
    .C1(_06281_),
    .Y(_06446_));
 sky130_fd_sc_hd__or2_1 _14964_ (.A(_06444_),
    .B(_06446_),
    .X(_06447_));
 sky130_fd_sc_hd__or2_1 _14965_ (.A(_06427_),
    .B(_06447_),
    .X(_06448_));
 sky130_fd_sc_hd__nand2_1 _14966_ (.A(_06427_),
    .B(_06447_),
    .Y(_06449_));
 sky130_fd_sc_hd__xnor2_1 _14967_ (.A(_06427_),
    .B(_06447_),
    .Y(_06450_));
 sky130_fd_sc_hd__xnor2_1 _14968_ (.A(_06409_),
    .B(_06450_),
    .Y(_06451_));
 sky130_fd_sc_hd__and2b_1 _14969_ (.A_N(_06408_),
    .B(_06451_),
    .X(_06452_));
 sky130_fd_sc_hd__xnor2_1 _14970_ (.A(_06408_),
    .B(_06451_),
    .Y(_06453_));
 sky130_fd_sc_hd__and3_2 _14971_ (.A(_06058_),
    .B(_06333_),
    .C(_06334_),
    .X(_06454_));
 sky130_fd_sc_hd__inv_2 _14972_ (.A(_06454_),
    .Y(_06455_));
 sky130_fd_sc_hd__nor2_2 _14973_ (.A(_06058_),
    .B(_06333_),
    .Y(_06456_));
 sky130_fd_sc_hd__or2_1 _14974_ (.A(_06058_),
    .B(_06333_),
    .X(_06457_));
 sky130_fd_sc_hd__nor2_2 _14975_ (.A(_06454_),
    .B(_06456_),
    .Y(_06458_));
 sky130_fd_sc_hd__nand2_1 _14976_ (.A(_06341_),
    .B(_06343_),
    .Y(_06459_));
 sky130_fd_sc_hd__a21o_2 _14977_ (.A1(net429),
    .A2(_06199_),
    .B1(_06197_),
    .X(_06460_));
 sky130_fd_sc_hd__a22o_1 _14978_ (.A1(net420),
    .A2(net456),
    .B1(net453),
    .B2(net424),
    .X(_06461_));
 sky130_fd_sc_hd__nand4_2 _14979_ (.A(net424),
    .B(net420),
    .C(net456),
    .D(net453),
    .Y(_06462_));
 sky130_fd_sc_hd__a22o_1 _14980_ (.A1(net415),
    .A2(\mul0.a[29] ),
    .B1(_06461_),
    .B2(_06462_),
    .X(_06463_));
 sky130_fd_sc_hd__nand4_2 _14981_ (.A(\mul0.b[8] ),
    .B(\mul0.a[29] ),
    .C(_06461_),
    .D(_06462_),
    .Y(_06464_));
 sky130_fd_sc_hd__nand3_1 _14982_ (.A(_06460_),
    .B(_06463_),
    .C(_06464_),
    .Y(_06465_));
 sky130_fd_sc_hd__a21o_1 _14983_ (.A1(_06463_),
    .A2(_06464_),
    .B1(_06460_),
    .X(_06466_));
 sky130_fd_sc_hd__nand3_1 _14984_ (.A(_06459_),
    .B(_06465_),
    .C(_06466_),
    .Y(_06467_));
 sky130_fd_sc_hd__a21o_1 _14985_ (.A1(_06465_),
    .A2(_06466_),
    .B1(_06459_),
    .X(_06468_));
 sky130_fd_sc_hd__a2bb2o_1 _14986_ (.A1_N(_06454_),
    .A2_N(_06456_),
    .B1(_06467_),
    .B2(_06468_),
    .X(_06469_));
 sky130_fd_sc_hd__or4bb_1 _14987_ (.A(_06454_),
    .B(_06456_),
    .C_N(_06467_),
    .D_N(_06468_),
    .X(_06470_));
 sky130_fd_sc_hd__a31o_1 _14988_ (.A1(_06337_),
    .A2(_06346_),
    .A3(_06347_),
    .B1(_06335_),
    .X(_06471_));
 sky130_fd_sc_hd__a21oi_2 _14989_ (.A1(_06469_),
    .A2(_06470_),
    .B1(_06471_),
    .Y(_06472_));
 sky130_fd_sc_hd__and3_2 _14990_ (.A(_06469_),
    .B(_06470_),
    .C(_06471_),
    .X(_06473_));
 sky130_fd_sc_hd__a21bo_1 _14991_ (.A1(_06338_),
    .A2(_06345_),
    .B1_N(_06344_),
    .X(_06474_));
 sky130_fd_sc_hd__a22o_1 _14992_ (.A1(net393),
    .A2(net475),
    .B1(net471),
    .B2(net399),
    .X(_06475_));
 sky130_fd_sc_hd__nand4_1 _14993_ (.A(net399),
    .B(net394),
    .C(net475),
    .D(net471),
    .Y(_06476_));
 sky130_fd_sc_hd__nand2_1 _14994_ (.A(_06475_),
    .B(_06476_),
    .Y(_06477_));
 sky130_fd_sc_hd__and2_1 _14995_ (.A(net389),
    .B(net479),
    .X(_06478_));
 sky130_fd_sc_hd__xnor2_1 _14996_ (.A(_06477_),
    .B(_06478_),
    .Y(_06479_));
 sky130_fd_sc_hd__a22o_1 _14997_ (.A1(net406),
    .A2(net463),
    .B1(net461),
    .B2(net410),
    .X(_06480_));
 sky130_fd_sc_hd__and4_1 _14998_ (.A(net410),
    .B(net406),
    .C(net464),
    .D(net461),
    .X(_06481_));
 sky130_fd_sc_hd__nand4_2 _14999_ (.A(net410),
    .B(net406),
    .C(net463),
    .D(net461),
    .Y(_06482_));
 sky130_fd_sc_hd__a22oi_4 _15000_ (.A1(net402),
    .A2(net466),
    .B1(_06480_),
    .B2(_06482_),
    .Y(_06483_));
 sky130_fd_sc_hd__and4_2 _15001_ (.A(net402),
    .B(net467),
    .C(_06480_),
    .D(_06482_),
    .X(_06484_));
 sky130_fd_sc_hd__a211o_1 _15002_ (.A1(_06360_),
    .A2(_06362_),
    .B1(_06483_),
    .C1(_06484_),
    .X(_06485_));
 sky130_fd_sc_hd__o211ai_2 _15003_ (.A1(_06483_),
    .A2(_06484_),
    .B1(_06360_),
    .C1(_06362_),
    .Y(_06486_));
 sky130_fd_sc_hd__nand3_2 _15004_ (.A(_06479_),
    .B(_06485_),
    .C(_06486_),
    .Y(_06487_));
 sky130_fd_sc_hd__a21o_1 _15005_ (.A1(_06485_),
    .A2(_06486_),
    .B1(_06479_),
    .X(_06488_));
 sky130_fd_sc_hd__and3_2 _15006_ (.A(_06474_),
    .B(_06487_),
    .C(_06488_),
    .X(_06489_));
 sky130_fd_sc_hd__a21oi_2 _15007_ (.A1(_06487_),
    .A2(_06488_),
    .B1(_06474_),
    .Y(_06490_));
 sky130_fd_sc_hd__a211oi_4 _15008_ (.A1(_06363_),
    .A2(_06365_),
    .B1(_06489_),
    .C1(_06490_),
    .Y(_06491_));
 sky130_fd_sc_hd__o211a_1 _15009_ (.A1(_06489_),
    .A2(_06490_),
    .B1(_06363_),
    .C1(_06365_),
    .X(_06492_));
 sky130_fd_sc_hd__o22ai_2 _15010_ (.A1(_06472_),
    .A2(_06473_),
    .B1(_06491_),
    .B2(_06492_),
    .Y(_06493_));
 sky130_fd_sc_hd__nor4_1 _15011_ (.A(_06472_),
    .B(_06473_),
    .C(_06491_),
    .D(_06492_),
    .Y(_06494_));
 sky130_fd_sc_hd__or4_1 _15012_ (.A(_06472_),
    .B(_06473_),
    .C(_06491_),
    .D(_06492_),
    .X(_06495_));
 sky130_fd_sc_hd__o211a_1 _15013_ (.A1(_06352_),
    .A2(_06371_),
    .B1(_06493_),
    .C1(_06495_),
    .X(_06496_));
 sky130_fd_sc_hd__a211oi_1 _15014_ (.A1(_06493_),
    .A2(_06495_),
    .B1(_06352_),
    .C1(_06371_),
    .Y(_06497_));
 sky130_fd_sc_hd__a22o_1 _15015_ (.A1(net509),
    .A2(net357),
    .B1(net352),
    .B2(net513),
    .X(_06498_));
 sky130_fd_sc_hd__nand4_1 _15016_ (.A(net509),
    .B(net513),
    .C(net357),
    .D(net352),
    .Y(_06499_));
 sky130_fd_sc_hd__nand2_1 _15017_ (.A(_06498_),
    .B(_06499_),
    .Y(_06500_));
 sky130_fd_sc_hd__and2_1 _15018_ (.A(net518),
    .B(net349),
    .X(_06501_));
 sky130_fd_sc_hd__xnor2_2 _15019_ (.A(_06500_),
    .B(_06501_),
    .Y(_06502_));
 sky130_fd_sc_hd__a22o_1 _15020_ (.A1(net634),
    .A2(net496),
    .B1(net368),
    .B2(net500),
    .X(_06503_));
 sky130_fd_sc_hd__nand4_1 _15021_ (.A(net500),
    .B(net634),
    .C(net496),
    .D(net368),
    .Y(_06504_));
 sky130_fd_sc_hd__and2_1 _15022_ (.A(net505),
    .B(net361),
    .X(_06505_));
 sky130_fd_sc_hd__a21o_1 _15023_ (.A1(_06503_),
    .A2(_06504_),
    .B1(_06505_),
    .X(_06506_));
 sky130_fd_sc_hd__nand3_1 _15024_ (.A(_06503_),
    .B(_06504_),
    .C(_06505_),
    .Y(_06507_));
 sky130_fd_sc_hd__o211a_1 _15025_ (.A1(_06300_),
    .A2(_06303_),
    .B1(_06506_),
    .C1(_06507_),
    .X(_06508_));
 sky130_fd_sc_hd__a211o_1 _15026_ (.A1(_06506_),
    .A2(_06507_),
    .B1(_06300_),
    .C1(_06303_),
    .X(_06509_));
 sky130_fd_sc_hd__nand2b_1 _15027_ (.A_N(_06508_),
    .B(_06509_),
    .Y(_06510_));
 sky130_fd_sc_hd__xnor2_2 _15028_ (.A(_06502_),
    .B(_06510_),
    .Y(_06511_));
 sky130_fd_sc_hd__nand2_1 _15029_ (.A(_06312_),
    .B(_06314_),
    .Y(_06512_));
 sky130_fd_sc_hd__a32o_1 _15030_ (.A1(net389),
    .A2(net483),
    .A3(_06354_),
    .B1(_06355_),
    .B2(net475),
    .X(_06513_));
 sky130_fd_sc_hd__a22o_1 _15031_ (.A1(net378),
    .A2(net488),
    .B1(net484),
    .B2(net384),
    .X(_06514_));
 sky130_fd_sc_hd__nand4_1 _15032_ (.A(net384),
    .B(net378),
    .C(net488),
    .D(net484),
    .Y(_06515_));
 sky130_fd_sc_hd__a22o_1 _15033_ (.A1(net373),
    .A2(net493),
    .B1(_06514_),
    .B2(_06515_),
    .X(_06516_));
 sky130_fd_sc_hd__nand4_1 _15034_ (.A(net373),
    .B(net493),
    .C(_06514_),
    .D(_06515_),
    .Y(_06517_));
 sky130_fd_sc_hd__nand3_1 _15035_ (.A(_06513_),
    .B(_06516_),
    .C(_06517_),
    .Y(_06518_));
 sky130_fd_sc_hd__a21o_1 _15036_ (.A1(_06516_),
    .A2(_06517_),
    .B1(_06513_),
    .X(_06519_));
 sky130_fd_sc_hd__nand3_1 _15037_ (.A(_06512_),
    .B(_06518_),
    .C(_06519_),
    .Y(_06520_));
 sky130_fd_sc_hd__a21o_1 _15038_ (.A1(_06518_),
    .A2(_06519_),
    .B1(_06512_),
    .X(_06521_));
 sky130_fd_sc_hd__a21bo_1 _15039_ (.A1(_06309_),
    .A2(_06316_),
    .B1_N(_06315_),
    .X(_06522_));
 sky130_fd_sc_hd__nand3_2 _15040_ (.A(_06520_),
    .B(_06521_),
    .C(_06522_),
    .Y(_06523_));
 sky130_fd_sc_hd__inv_2 _15041_ (.A(_06523_),
    .Y(_06524_));
 sky130_fd_sc_hd__a21o_1 _15042_ (.A1(_06520_),
    .A2(_06521_),
    .B1(_06522_),
    .X(_06525_));
 sky130_fd_sc_hd__and3_1 _15043_ (.A(_06511_),
    .B(_06523_),
    .C(_06525_),
    .X(_06526_));
 sky130_fd_sc_hd__nand3_2 _15044_ (.A(_06511_),
    .B(_06523_),
    .C(_06525_),
    .Y(_06527_));
 sky130_fd_sc_hd__a21o_1 _15045_ (.A1(_06523_),
    .A2(_06525_),
    .B1(_06511_),
    .X(_06528_));
 sky130_fd_sc_hd__o211ai_4 _15046_ (.A1(_06367_),
    .A2(_06369_),
    .B1(_06527_),
    .C1(_06528_),
    .Y(_06529_));
 sky130_fd_sc_hd__a211o_1 _15047_ (.A1(_06527_),
    .A2(_06528_),
    .B1(_06367_),
    .C1(_06369_),
    .X(_06530_));
 sky130_fd_sc_hd__o211ai_4 _15048_ (.A1(_06321_),
    .A2(_06323_),
    .B1(_06529_),
    .C1(_06530_),
    .Y(_06531_));
 sky130_fd_sc_hd__a211o_1 _15049_ (.A1(_06529_),
    .A2(_06530_),
    .B1(_06321_),
    .C1(_06323_),
    .X(_06532_));
 sky130_fd_sc_hd__and4bb_1 _15050_ (.A_N(_06496_),
    .B_N(_06497_),
    .C(_06531_),
    .D(_06532_),
    .X(_06533_));
 sky130_fd_sc_hd__a2bb2o_1 _15051_ (.A1_N(_06496_),
    .A2_N(_06497_),
    .B1(_06531_),
    .B2(_06532_),
    .X(_06534_));
 sky130_fd_sc_hd__and2b_1 _15052_ (.A_N(_06533_),
    .B(_06534_),
    .X(_06535_));
 sky130_fd_sc_hd__a21o_1 _15053_ (.A1(_06330_),
    .A2(_06376_),
    .B1(_06375_),
    .X(_06536_));
 sky130_fd_sc_hd__nand2_1 _15054_ (.A(_06535_),
    .B(_06536_),
    .Y(_06537_));
 sky130_fd_sc_hd__xor2_2 _15055_ (.A(_06535_),
    .B(_06536_),
    .X(_06538_));
 sky130_fd_sc_hd__xor2_1 _15056_ (.A(_06453_),
    .B(_06538_),
    .X(_06539_));
 sky130_fd_sc_hd__a21oi_1 _15057_ (.A1(_06292_),
    .A2(_06380_),
    .B1(_06379_),
    .Y(_06540_));
 sky130_fd_sc_hd__nand2b_1 _15058_ (.A_N(_06540_),
    .B(_06539_),
    .Y(_06541_));
 sky130_fd_sc_hd__xnor2_1 _15059_ (.A(_06539_),
    .B(_06540_),
    .Y(_06542_));
 sky130_fd_sc_hd__xnor2_1 _15060_ (.A(_06407_),
    .B(_06542_),
    .Y(_06543_));
 sky130_fd_sc_hd__a21boi_1 _15061_ (.A1(_06248_),
    .A2(_06384_),
    .B1_N(_06383_),
    .Y(_06544_));
 sky130_fd_sc_hd__or2_1 _15062_ (.A(_06543_),
    .B(_06544_),
    .X(_06545_));
 sky130_fd_sc_hd__xor2_1 _15063_ (.A(_06543_),
    .B(_06544_),
    .X(_06546_));
 sky130_fd_sc_hd__nand2_1 _15064_ (.A(_06406_),
    .B(_06546_),
    .Y(_06547_));
 sky130_fd_sc_hd__xnor2_1 _15065_ (.A(_06406_),
    .B(_06546_),
    .Y(_06548_));
 sky130_fd_sc_hd__a21oi_1 _15066_ (.A1(_06387_),
    .A2(_06389_),
    .B1(_06548_),
    .Y(_06549_));
 sky130_fd_sc_hd__and3_1 _15067_ (.A(_06387_),
    .B(_06389_),
    .C(_06548_),
    .X(_06550_));
 sky130_fd_sc_hd__nor2_2 _15068_ (.A(_06549_),
    .B(_06550_),
    .Y(_06551_));
 sky130_fd_sc_hd__xnor2_4 _15069_ (.A(_06405_),
    .B(_06551_),
    .Y(_06552_));
 sky130_fd_sc_hd__nor2_1 _15070_ (.A(net9),
    .B(_06552_),
    .Y(_06553_));
 sky130_fd_sc_hd__a221o_1 _15071_ (.A1(\state[4] ),
    .A2(net733),
    .B1(_02677_),
    .B2(_03794_),
    .C1(_06553_),
    .X(_06554_));
 sky130_fd_sc_hd__mux2_1 _15072_ (.A0(net851),
    .A1(_06554_),
    .S(_03055_),
    .X(_00287_));
 sky130_fd_sc_hd__a21o_1 _15073_ (.A1(_06423_),
    .A2(_06424_),
    .B1(_06426_),
    .X(_06555_));
 sky130_fd_sc_hd__a31o_1 _15074_ (.A1(_06409_),
    .A2(_06448_),
    .A3(_06449_),
    .B1(_06452_),
    .X(_06556_));
 sky130_fd_sc_hd__nand2_1 _15075_ (.A(_06462_),
    .B(_06464_),
    .Y(_06557_));
 sky130_fd_sc_hd__nand3_4 _15076_ (.A(net424),
    .B(net420),
    .C(net453),
    .Y(_06558_));
 sky130_fd_sc_hd__o21a_1 _15077_ (.A1(net424),
    .A2(net420),
    .B1(net453),
    .X(_06559_));
 sky130_fd_sc_hd__a22o_1 _15078_ (.A1(net416),
    .A2(net456),
    .B1(_06558_),
    .B2(_06559_),
    .X(_06560_));
 sky130_fd_sc_hd__nand4_2 _15079_ (.A(net416),
    .B(net456),
    .C(_06558_),
    .D(_06559_),
    .Y(_06561_));
 sky130_fd_sc_hd__nand3_1 _15080_ (.A(_06460_),
    .B(_06560_),
    .C(_06561_),
    .Y(_06562_));
 sky130_fd_sc_hd__a21o_1 _15081_ (.A1(_06560_),
    .A2(_06561_),
    .B1(_06460_),
    .X(_06563_));
 sky130_fd_sc_hd__and3_1 _15082_ (.A(_06557_),
    .B(_06562_),
    .C(_06563_),
    .X(_06564_));
 sky130_fd_sc_hd__a21oi_1 _15083_ (.A1(_06562_),
    .A2(_06563_),
    .B1(_06557_),
    .Y(_06565_));
 sky130_fd_sc_hd__o22ai_1 _15084_ (.A1(_06454_),
    .A2(_06456_),
    .B1(_06564_),
    .B2(_06565_),
    .Y(_06566_));
 sky130_fd_sc_hd__or4_1 _15085_ (.A(_06454_),
    .B(_06456_),
    .C(_06564_),
    .D(_06565_),
    .X(_06567_));
 sky130_fd_sc_hd__a31o_1 _15086_ (.A1(_06457_),
    .A2(_06467_),
    .A3(_06468_),
    .B1(_06454_),
    .X(_06568_));
 sky130_fd_sc_hd__and3_1 _15087_ (.A(_06566_),
    .B(_06567_),
    .C(_06568_),
    .X(_06569_));
 sky130_fd_sc_hd__a21oi_1 _15088_ (.A1(_06566_),
    .A2(_06567_),
    .B1(_06568_),
    .Y(_06570_));
 sky130_fd_sc_hd__a21bo_1 _15089_ (.A1(_06459_),
    .A2(_06466_),
    .B1_N(_06465_),
    .X(_06571_));
 sky130_fd_sc_hd__a22o_1 _15090_ (.A1(net393),
    .A2(net473),
    .B1(net467),
    .B2(net398),
    .X(_06572_));
 sky130_fd_sc_hd__and3_1 _15091_ (.A(net398),
    .B(net393),
    .C(net473),
    .X(_06573_));
 sky130_fd_sc_hd__a21bo_1 _15092_ (.A1(net467),
    .A2(_06573_),
    .B1_N(_06572_),
    .X(_06574_));
 sky130_fd_sc_hd__nand2_1 _15093_ (.A(net388),
    .B(net477),
    .Y(_06575_));
 sky130_fd_sc_hd__xor2_1 _15094_ (.A(_06574_),
    .B(_06575_),
    .X(_06576_));
 sky130_fd_sc_hd__a22o_1 _15095_ (.A1(net406),
    .A2(net461),
    .B1(net459),
    .B2(net410),
    .X(_06577_));
 sky130_fd_sc_hd__nand4_4 _15096_ (.A(net410),
    .B(net406),
    .C(net461),
    .D(net459),
    .Y(_06578_));
 sky130_fd_sc_hd__a22o_1 _15097_ (.A1(net402),
    .A2(net463),
    .B1(_06577_),
    .B2(_06578_),
    .X(_06579_));
 sky130_fd_sc_hd__nand4_4 _15098_ (.A(net402),
    .B(net463),
    .C(_06577_),
    .D(_06578_),
    .Y(_06580_));
 sky130_fd_sc_hd__o211ai_4 _15099_ (.A1(_06481_),
    .A2(_06484_),
    .B1(_06579_),
    .C1(_06580_),
    .Y(_06581_));
 sky130_fd_sc_hd__a211o_1 _15100_ (.A1(_06579_),
    .A2(_06580_),
    .B1(_06481_),
    .C1(_06484_),
    .X(_06582_));
 sky130_fd_sc_hd__nand3_2 _15101_ (.A(_06576_),
    .B(_06581_),
    .C(_06582_),
    .Y(_06583_));
 sky130_fd_sc_hd__a21o_1 _15102_ (.A1(_06581_),
    .A2(_06582_),
    .B1(_06576_),
    .X(_06584_));
 sky130_fd_sc_hd__and3_1 _15103_ (.A(_06571_),
    .B(_06583_),
    .C(_06584_),
    .X(_06585_));
 sky130_fd_sc_hd__a21oi_2 _15104_ (.A1(_06583_),
    .A2(_06584_),
    .B1(_06571_),
    .Y(_06586_));
 sky130_fd_sc_hd__a211oi_2 _15105_ (.A1(_06485_),
    .A2(_06487_),
    .B1(_06585_),
    .C1(_06586_),
    .Y(_06587_));
 sky130_fd_sc_hd__o211a_1 _15106_ (.A1(_06585_),
    .A2(_06586_),
    .B1(_06485_),
    .C1(_06487_),
    .X(_06588_));
 sky130_fd_sc_hd__o22ai_2 _15107_ (.A1(_06569_),
    .A2(_06570_),
    .B1(_06587_),
    .B2(_06588_),
    .Y(_06589_));
 sky130_fd_sc_hd__or4_2 _15108_ (.A(_06569_),
    .B(_06570_),
    .C(_06587_),
    .D(_06588_),
    .X(_06590_));
 sky130_fd_sc_hd__a211oi_2 _15109_ (.A1(_06589_),
    .A2(_06590_),
    .B1(_06473_),
    .C1(_06494_),
    .Y(_06591_));
 sky130_fd_sc_hd__o211a_2 _15110_ (.A1(_06473_),
    .A2(_06494_),
    .B1(_06589_),
    .C1(_06590_),
    .X(_06592_));
 sky130_fd_sc_hd__a22o_1 _15111_ (.A1(net505),
    .A2(net357),
    .B1(net352),
    .B2(net509),
    .X(_06593_));
 sky130_fd_sc_hd__and4_1 _15112_ (.A(net505),
    .B(net509),
    .C(net357),
    .D(net352),
    .X(_06594_));
 sky130_fd_sc_hd__inv_2 _15113_ (.A(_06594_),
    .Y(_06595_));
 sky130_fd_sc_hd__a22oi_1 _15114_ (.A1(net513),
    .A2(net349),
    .B1(_06593_),
    .B2(_06595_),
    .Y(_06596_));
 sky130_fd_sc_hd__and4_1 _15115_ (.A(net513),
    .B(net349),
    .C(_06593_),
    .D(_06595_),
    .X(_06597_));
 sky130_fd_sc_hd__or2_1 _15116_ (.A(_06596_),
    .B(_06597_),
    .X(_06598_));
 sky130_fd_sc_hd__a22o_1 _15117_ (.A1(net496),
    .A2(net368),
    .B1(net492),
    .B2(net634),
    .X(_06599_));
 sky130_fd_sc_hd__nand4_2 _15118_ (.A(net634),
    .B(net496),
    .C(net368),
    .D(net492),
    .Y(_06600_));
 sky130_fd_sc_hd__a22o_1 _15119_ (.A1(net500),
    .A2(net361),
    .B1(_06599_),
    .B2(_06600_),
    .X(_06601_));
 sky130_fd_sc_hd__nand4_2 _15120_ (.A(net500),
    .B(net362),
    .C(_06599_),
    .D(_06600_),
    .Y(_06602_));
 sky130_fd_sc_hd__a21bo_1 _15121_ (.A1(_06503_),
    .A2(_06505_),
    .B1_N(_06504_),
    .X(_06603_));
 sky130_fd_sc_hd__nand3_2 _15122_ (.A(_06601_),
    .B(_06602_),
    .C(_06603_),
    .Y(_06604_));
 sky130_fd_sc_hd__a21o_1 _15123_ (.A1(_06601_),
    .A2(_06602_),
    .B1(_06603_),
    .X(_06605_));
 sky130_fd_sc_hd__nand2_1 _15124_ (.A(_06604_),
    .B(_06605_),
    .Y(_06606_));
 sky130_fd_sc_hd__or2_1 _15125_ (.A(_06598_),
    .B(_06606_),
    .X(_06607_));
 sky130_fd_sc_hd__xor2_2 _15126_ (.A(_06598_),
    .B(_06606_),
    .X(_06608_));
 sky130_fd_sc_hd__nand2_1 _15127_ (.A(_06515_),
    .B(_06517_),
    .Y(_06609_));
 sky130_fd_sc_hd__a21boi_1 _15128_ (.A1(_06475_),
    .A2(_06478_),
    .B1_N(_06476_),
    .Y(_06610_));
 sky130_fd_sc_hd__a22oi_1 _15129_ (.A1(net378),
    .A2(net484),
    .B1(net479),
    .B2(net384),
    .Y(_06611_));
 sky130_fd_sc_hd__and4_1 _15130_ (.A(net385),
    .B(net379),
    .C(net484),
    .D(net479),
    .X(_06612_));
 sky130_fd_sc_hd__o2bb2a_1 _15131_ (.A1_N(net373),
    .A2_N(net488),
    .B1(_06611_),
    .B2(_06612_),
    .X(_06613_));
 sky130_fd_sc_hd__and4bb_1 _15132_ (.A_N(_06611_),
    .B_N(_06612_),
    .C(net373),
    .D(net488),
    .X(_06614_));
 sky130_fd_sc_hd__or3_2 _15133_ (.A(_06610_),
    .B(_06613_),
    .C(_06614_),
    .X(_06615_));
 sky130_fd_sc_hd__o21ai_1 _15134_ (.A1(_06613_),
    .A2(_06614_),
    .B1(_06610_),
    .Y(_06616_));
 sky130_fd_sc_hd__nand3_1 _15135_ (.A(_06609_),
    .B(_06615_),
    .C(_06616_),
    .Y(_06617_));
 sky130_fd_sc_hd__a21o_1 _15136_ (.A1(_06615_),
    .A2(_06616_),
    .B1(_06609_),
    .X(_06618_));
 sky130_fd_sc_hd__a21bo_1 _15137_ (.A1(_06512_),
    .A2(_06519_),
    .B1_N(_06518_),
    .X(_06619_));
 sky130_fd_sc_hd__nand3_1 _15138_ (.A(_06617_),
    .B(_06618_),
    .C(_06619_),
    .Y(_06620_));
 sky130_fd_sc_hd__a21o_1 _15139_ (.A1(_06617_),
    .A2(_06618_),
    .B1(_06619_),
    .X(_06621_));
 sky130_fd_sc_hd__nand3_2 _15140_ (.A(_06608_),
    .B(_06620_),
    .C(_06621_),
    .Y(_06622_));
 sky130_fd_sc_hd__a21o_1 _15141_ (.A1(_06620_),
    .A2(_06621_),
    .B1(_06608_),
    .X(_06623_));
 sky130_fd_sc_hd__o211ai_4 _15142_ (.A1(_06489_),
    .A2(_06491_),
    .B1(_06622_),
    .C1(_06623_),
    .Y(_06624_));
 sky130_fd_sc_hd__a211o_1 _15143_ (.A1(_06622_),
    .A2(_06623_),
    .B1(_06489_),
    .C1(_06491_),
    .X(_06625_));
 sky130_fd_sc_hd__o211ai_2 _15144_ (.A1(_06524_),
    .A2(_06526_),
    .B1(_06624_),
    .C1(_06625_),
    .Y(_06626_));
 sky130_fd_sc_hd__a211o_1 _15145_ (.A1(_06624_),
    .A2(_06625_),
    .B1(_06524_),
    .C1(_06526_),
    .X(_06627_));
 sky130_fd_sc_hd__and4bb_1 _15146_ (.A_N(_06591_),
    .B_N(_06592_),
    .C(_06626_),
    .D(_06627_),
    .X(_06628_));
 sky130_fd_sc_hd__or4bb_1 _15147_ (.A(_06591_),
    .B(_06592_),
    .C_N(_06626_),
    .D_N(_06627_),
    .X(_06629_));
 sky130_fd_sc_hd__a2bb2o_1 _15148_ (.A1_N(_06591_),
    .A2_N(_06592_),
    .B1(_06626_),
    .B2(_06627_),
    .X(_06630_));
 sky130_fd_sc_hd__o211a_2 _15149_ (.A1(_06496_),
    .A2(_06533_),
    .B1(_06629_),
    .C1(_06630_),
    .X(_06631_));
 sky130_fd_sc_hd__a211oi_1 _15150_ (.A1(_06629_),
    .A2(_06630_),
    .B1(_06496_),
    .C1(_06533_),
    .Y(_06632_));
 sky130_fd_sc_hd__nor2_2 _15151_ (.A(_06631_),
    .B(_06632_),
    .Y(_06633_));
 sky130_fd_sc_hd__a22oi_1 _15152_ (.A1(net534),
    .A2(net334),
    .B1(net331),
    .B2(net538),
    .Y(_06634_));
 sky130_fd_sc_hd__and4_1 _15153_ (.A(net533),
    .B(net538),
    .C(net334),
    .D(net331),
    .X(_06635_));
 sky130_fd_sc_hd__o2bb2a_1 _15154_ (.A1_N(net543),
    .A2_N(net329),
    .B1(_06634_),
    .B2(_06635_),
    .X(_06636_));
 sky130_fd_sc_hd__and4bb_1 _15155_ (.A_N(_06634_),
    .B_N(_06635_),
    .C(net543),
    .D(net329),
    .X(_06637_));
 sky130_fd_sc_hd__o211a_1 _15156_ (.A1(_06636_),
    .A2(_06637_),
    .B1(_06411_),
    .C1(_06413_),
    .X(_06638_));
 sky130_fd_sc_hd__a211o_1 _15157_ (.A1(_06411_),
    .A2(_06413_),
    .B1(_06636_),
    .C1(_06637_),
    .X(_06639_));
 sky130_fd_sc_hd__nand2b_1 _15158_ (.A_N(_06638_),
    .B(_06639_),
    .Y(_06640_));
 sky130_fd_sc_hd__and4b_1 _15159_ (.A_N(\mul0.a[7] ),
    .B(net327),
    .C(net326),
    .D(net547),
    .X(_06641_));
 sky130_fd_sc_hd__inv_2 _15160_ (.A(_06641_),
    .Y(_06642_));
 sky130_fd_sc_hd__o2bb2a_1 _15161_ (.A1_N(\mul0.a[8] ),
    .A2_N(net327),
    .B1(net57),
    .B2(\mul0.a[7] ),
    .X(_06643_));
 sky130_fd_sc_hd__nor2_1 _15162_ (.A(_06641_),
    .B(_06643_),
    .Y(_06644_));
 sky130_fd_sc_hd__xnor2_2 _15163_ (.A(_06640_),
    .B(_06644_),
    .Y(_06645_));
 sky130_fd_sc_hd__a21o_1 _15164_ (.A1(_06416_),
    .A2(_06422_),
    .B1(_06417_),
    .X(_06646_));
 sky130_fd_sc_hd__nand2_1 _15165_ (.A(_06645_),
    .B(_06646_),
    .Y(_06647_));
 sky130_fd_sc_hd__xnor2_2 _15166_ (.A(_06645_),
    .B(_06646_),
    .Y(_06648_));
 sky130_fd_sc_hd__xnor2_1 _15167_ (.A(_06420_),
    .B(_06648_),
    .Y(_06649_));
 sky130_fd_sc_hd__a21o_1 _15168_ (.A1(_06502_),
    .A2(_06509_),
    .B1(_06508_),
    .X(_06650_));
 sky130_fd_sc_hd__nand2_1 _15169_ (.A(_06432_),
    .B(_06434_),
    .Y(_06651_));
 sky130_fd_sc_hd__a21boi_1 _15170_ (.A1(_06498_),
    .A2(_06501_),
    .B1_N(_06499_),
    .Y(_06652_));
 sky130_fd_sc_hd__a22oi_1 _15171_ (.A1(net518),
    .A2(net346),
    .B1(net342),
    .B2(net522),
    .Y(_06653_));
 sky130_fd_sc_hd__and4_1 _15172_ (.A(net518),
    .B(net522),
    .C(net346),
    .D(net342),
    .X(_06654_));
 sky130_fd_sc_hd__o2bb2a_1 _15173_ (.A1_N(net528),
    .A2_N(net339),
    .B1(_06653_),
    .B2(_06654_),
    .X(_06655_));
 sky130_fd_sc_hd__and4bb_1 _15174_ (.A_N(_06653_),
    .B_N(_06654_),
    .C(net528),
    .D(net339),
    .X(_06656_));
 sky130_fd_sc_hd__or3_2 _15175_ (.A(_06652_),
    .B(_06655_),
    .C(_06656_),
    .X(_06657_));
 sky130_fd_sc_hd__o21ai_1 _15176_ (.A1(_06655_),
    .A2(_06656_),
    .B1(_06652_),
    .Y(_06658_));
 sky130_fd_sc_hd__nand3_2 _15177_ (.A(_06651_),
    .B(_06657_),
    .C(_06658_),
    .Y(_06659_));
 sky130_fd_sc_hd__a21o_1 _15178_ (.A1(_06657_),
    .A2(_06658_),
    .B1(_06651_),
    .X(_06660_));
 sky130_fd_sc_hd__and3_1 _15179_ (.A(_06650_),
    .B(_06659_),
    .C(_06660_),
    .X(_06661_));
 sky130_fd_sc_hd__a21oi_1 _15180_ (.A1(_06659_),
    .A2(_06660_),
    .B1(_06650_),
    .Y(_06662_));
 sky130_fd_sc_hd__a211o_1 _15181_ (.A1(_06435_),
    .A2(_06437_),
    .B1(_06661_),
    .C1(_06662_),
    .X(_06663_));
 sky130_fd_sc_hd__o211ai_1 _15182_ (.A1(_06661_),
    .A2(_06662_),
    .B1(_06435_),
    .C1(_06437_),
    .Y(_06664_));
 sky130_fd_sc_hd__o211a_1 _15183_ (.A1(_06439_),
    .A2(_06441_),
    .B1(_06663_),
    .C1(_06664_),
    .X(_06665_));
 sky130_fd_sc_hd__a211oi_1 _15184_ (.A1(_06663_),
    .A2(_06664_),
    .B1(_06439_),
    .C1(_06441_),
    .Y(_06666_));
 sky130_fd_sc_hd__nor3_1 _15185_ (.A(_06649_),
    .B(_06665_),
    .C(_06666_),
    .Y(_06667_));
 sky130_fd_sc_hd__o21a_1 _15186_ (.A1(_06665_),
    .A2(_06666_),
    .B1(_06649_),
    .X(_06668_));
 sky130_fd_sc_hd__a211oi_2 _15187_ (.A1(_06529_),
    .A2(_06531_),
    .B1(_06667_),
    .C1(_06668_),
    .Y(_06669_));
 sky130_fd_sc_hd__o211a_1 _15188_ (.A1(_06667_),
    .A2(_06668_),
    .B1(_06529_),
    .C1(_06531_),
    .X(_06670_));
 sky130_fd_sc_hd__a211oi_1 _15189_ (.A1(_06445_),
    .A2(_06448_),
    .B1(_06669_),
    .C1(_06670_),
    .Y(_06671_));
 sky130_fd_sc_hd__o211a_1 _15190_ (.A1(_06669_),
    .A2(_06670_),
    .B1(_06445_),
    .C1(_06448_),
    .X(_06672_));
 sky130_fd_sc_hd__nor2_2 _15191_ (.A(_06671_),
    .B(_06672_),
    .Y(_06673_));
 sky130_fd_sc_hd__xnor2_1 _15192_ (.A(_06633_),
    .B(_06673_),
    .Y(_06674_));
 sky130_fd_sc_hd__a21boi_2 _15193_ (.A1(_06453_),
    .A2(_06538_),
    .B1_N(_06537_),
    .Y(_06675_));
 sky130_fd_sc_hd__nor2_1 _15194_ (.A(_06674_),
    .B(_06675_),
    .Y(_06676_));
 sky130_fd_sc_hd__xor2_1 _15195_ (.A(_06674_),
    .B(_06675_),
    .X(_06677_));
 sky130_fd_sc_hd__xnor2_1 _15196_ (.A(_06556_),
    .B(_06677_),
    .Y(_06678_));
 sky130_fd_sc_hd__a21boi_1 _15197_ (.A1(_06407_),
    .A2(_06542_),
    .B1_N(_06541_),
    .Y(_06679_));
 sky130_fd_sc_hd__nor2_1 _15198_ (.A(_06678_),
    .B(_06679_),
    .Y(_06680_));
 sky130_fd_sc_hd__and2_1 _15199_ (.A(_06678_),
    .B(_06679_),
    .X(_06681_));
 sky130_fd_sc_hd__nor2_1 _15200_ (.A(_06680_),
    .B(_06681_),
    .Y(_06682_));
 sky130_fd_sc_hd__xnor2_1 _15201_ (.A(_06555_),
    .B(_06682_),
    .Y(_06683_));
 sky130_fd_sc_hd__a21oi_2 _15202_ (.A1(_06545_),
    .A2(_06547_),
    .B1(_06683_),
    .Y(_06684_));
 sky130_fd_sc_hd__and3_1 _15203_ (.A(_06545_),
    .B(_06547_),
    .C(_06683_),
    .X(_06685_));
 sky130_fd_sc_hd__or2_2 _15204_ (.A(_06684_),
    .B(_06685_),
    .X(_06686_));
 sky130_fd_sc_hd__o21ba_1 _15205_ (.A1(_06392_),
    .A2(_06549_),
    .B1_N(_06550_),
    .X(_06687_));
 sky130_fd_sc_hd__and2_1 _15206_ (.A(_06394_),
    .B(_06551_),
    .X(_06688_));
 sky130_fd_sc_hd__inv_2 _15207_ (.A(_06688_),
    .Y(_06689_));
 sky130_fd_sc_hd__o21ba_2 _15208_ (.A1(_06400_),
    .A2(_06689_),
    .B1_N(_06687_),
    .X(_06690_));
 sky130_fd_sc_hd__xnor2_4 _15209_ (.A(_06686_),
    .B(_06690_),
    .Y(_06691_));
 sky130_fd_sc_hd__nor2_1 _15210_ (.A(net9),
    .B(_06691_),
    .Y(_06692_));
 sky130_fd_sc_hd__a221o_1 _15211_ (.A1(\state[4] ),
    .A2(net684),
    .B1(_02683_),
    .B2(net5),
    .C1(_06692_),
    .X(_06693_));
 sky130_fd_sc_hd__mux2_1 _15212_ (.A0(net666),
    .A1(net685),
    .S(net4),
    .X(_00288_));
 sky130_fd_sc_hd__a21o_2 _15213_ (.A1(_06555_),
    .A2(_06682_),
    .B1(_06680_),
    .X(_06694_));
 sky130_fd_sc_hd__o21ai_4 _15214_ (.A1(_06420_),
    .A2(_06648_),
    .B1(_06647_),
    .Y(_06695_));
 sky130_fd_sc_hd__nand2_1 _15215_ (.A(_06558_),
    .B(_06561_),
    .Y(_06696_));
 sky130_fd_sc_hd__a22o_1 _15216_ (.A1(net416),
    .A2(net454),
    .B1(_06558_),
    .B2(_06559_),
    .X(_06697_));
 sky130_fd_sc_hd__nand4_2 _15217_ (.A(net416),
    .B(net454),
    .C(_06558_),
    .D(_06559_),
    .Y(_06698_));
 sky130_fd_sc_hd__and3_1 _15218_ (.A(_06460_),
    .B(_06697_),
    .C(_06698_),
    .X(_06699_));
 sky130_fd_sc_hd__a21o_1 _15219_ (.A1(_06697_),
    .A2(_06698_),
    .B1(_06460_),
    .X(_06700_));
 sky130_fd_sc_hd__and2b_1 _15220_ (.A_N(_06699_),
    .B(_06700_),
    .X(_06701_));
 sky130_fd_sc_hd__xor2_2 _15221_ (.A(_06696_),
    .B(_06701_),
    .X(_06702_));
 sky130_fd_sc_hd__xnor2_2 _15222_ (.A(_06458_),
    .B(_06702_),
    .Y(_06703_));
 sky130_fd_sc_hd__nand2_1 _15223_ (.A(_06455_),
    .B(_06567_),
    .Y(_06704_));
 sky130_fd_sc_hd__nand2b_1 _15224_ (.A_N(_06703_),
    .B(_06704_),
    .Y(_06705_));
 sky130_fd_sc_hd__xnor2_2 _15225_ (.A(_06703_),
    .B(_06704_),
    .Y(_06706_));
 sky130_fd_sc_hd__nand2_2 _15226_ (.A(_06581_),
    .B(_06583_),
    .Y(_06707_));
 sky130_fd_sc_hd__a31o_1 _15227_ (.A1(_06460_),
    .A2(_06560_),
    .A3(_06561_),
    .B1(_06564_),
    .X(_06708_));
 sky130_fd_sc_hd__a22o_1 _15228_ (.A1(net393),
    .A2(net468),
    .B1(net465),
    .B2(net398),
    .X(_06709_));
 sky130_fd_sc_hd__nand4_2 _15229_ (.A(net398),
    .B(net393),
    .C(net466),
    .D(net465),
    .Y(_06710_));
 sky130_fd_sc_hd__a22o_1 _15230_ (.A1(net388),
    .A2(net470),
    .B1(_06709_),
    .B2(_06710_),
    .X(_06711_));
 sky130_fd_sc_hd__nand4_1 _15231_ (.A(net388),
    .B(net471),
    .C(_06709_),
    .D(_06710_),
    .Y(_06712_));
 sky130_fd_sc_hd__nand2_1 _15232_ (.A(_06711_),
    .B(_06712_),
    .Y(_06713_));
 sky130_fd_sc_hd__a22oi_1 _15233_ (.A1(net406),
    .A2(net458),
    .B1(net455),
    .B2(net410),
    .Y(_06714_));
 sky130_fd_sc_hd__and4_1 _15234_ (.A(net410),
    .B(net406),
    .C(net459),
    .D(net455),
    .X(_06715_));
 sky130_fd_sc_hd__o2bb2a_1 _15235_ (.A1_N(net402),
    .A2_N(net461),
    .B1(_06714_),
    .B2(_06715_),
    .X(_06716_));
 sky130_fd_sc_hd__and4bb_1 _15236_ (.A_N(_06714_),
    .B_N(_06715_),
    .C(net402),
    .D(net461),
    .X(_06717_));
 sky130_fd_sc_hd__nor2_1 _15237_ (.A(_06716_),
    .B(_06717_),
    .Y(_06718_));
 sky130_fd_sc_hd__nand2_1 _15238_ (.A(_06578_),
    .B(_06580_),
    .Y(_06719_));
 sky130_fd_sc_hd__nand2_1 _15239_ (.A(_06718_),
    .B(_06719_),
    .Y(_06720_));
 sky130_fd_sc_hd__xnor2_2 _15240_ (.A(_06718_),
    .B(_06719_),
    .Y(_06721_));
 sky130_fd_sc_hd__or2_1 _15241_ (.A(_06713_),
    .B(_06721_),
    .X(_06722_));
 sky130_fd_sc_hd__xor2_2 _15242_ (.A(_06713_),
    .B(_06721_),
    .X(_06723_));
 sky130_fd_sc_hd__and2_2 _15243_ (.A(_06708_),
    .B(_06723_),
    .X(_06724_));
 sky130_fd_sc_hd__xnor2_2 _15244_ (.A(_06708_),
    .B(_06723_),
    .Y(_06725_));
 sky130_fd_sc_hd__nand2b_2 _15245_ (.A_N(_06725_),
    .B(_06707_),
    .Y(_06726_));
 sky130_fd_sc_hd__inv_2 _15246_ (.A(_06726_),
    .Y(_06727_));
 sky130_fd_sc_hd__xnor2_2 _15247_ (.A(_06707_),
    .B(_06725_),
    .Y(_06728_));
 sky130_fd_sc_hd__nand2_1 _15248_ (.A(_06706_),
    .B(_06728_),
    .Y(_06729_));
 sky130_fd_sc_hd__xnor2_2 _15249_ (.A(_06706_),
    .B(_06728_),
    .Y(_06730_));
 sky130_fd_sc_hd__nand2b_2 _15250_ (.A_N(_06569_),
    .B(_06590_),
    .Y(_06731_));
 sky130_fd_sc_hd__nand2b_2 _15251_ (.A_N(_06730_),
    .B(_06731_),
    .Y(_06732_));
 sky130_fd_sc_hd__xnor2_1 _15252_ (.A(_06730_),
    .B(_06731_),
    .Y(_06733_));
 sky130_fd_sc_hd__and2_1 _15253_ (.A(_06620_),
    .B(_06622_),
    .X(_06734_));
 sky130_fd_sc_hd__nor2_1 _15254_ (.A(_06585_),
    .B(_06587_),
    .Y(_06735_));
 sky130_fd_sc_hd__a22o_1 _15255_ (.A1(net500),
    .A2(net357),
    .B1(net353),
    .B2(net506),
    .X(_06736_));
 sky130_fd_sc_hd__nand4_2 _15256_ (.A(net505),
    .B(net500),
    .C(net357),
    .D(net353),
    .Y(_06737_));
 sky130_fd_sc_hd__a22o_1 _15257_ (.A1(net509),
    .A2(net350),
    .B1(_06736_),
    .B2(_06737_),
    .X(_06738_));
 sky130_fd_sc_hd__nand4_1 _15258_ (.A(net509),
    .B(net350),
    .C(_06736_),
    .D(_06737_),
    .Y(_06739_));
 sky130_fd_sc_hd__nand2_1 _15259_ (.A(_06738_),
    .B(_06739_),
    .Y(_06740_));
 sky130_fd_sc_hd__a22o_1 _15260_ (.A1(net368),
    .A2(net492),
    .B1(net489),
    .B2(net634),
    .X(_06741_));
 sky130_fd_sc_hd__and4_1 _15261_ (.A(net634),
    .B(net368),
    .C(net492),
    .D(net489),
    .X(_06742_));
 sky130_fd_sc_hd__inv_2 _15262_ (.A(_06742_),
    .Y(_06743_));
 sky130_fd_sc_hd__a22oi_1 _15263_ (.A1(net496),
    .A2(net362),
    .B1(_06741_),
    .B2(_06743_),
    .Y(_06744_));
 sky130_fd_sc_hd__and4_1 _15264_ (.A(net497),
    .B(net362),
    .C(_06741_),
    .D(_06743_),
    .X(_06745_));
 sky130_fd_sc_hd__or2_1 _15265_ (.A(_06744_),
    .B(_06745_),
    .X(_06746_));
 sky130_fd_sc_hd__nand2_1 _15266_ (.A(_06600_),
    .B(_06602_),
    .Y(_06747_));
 sky130_fd_sc_hd__or3b_2 _15267_ (.A(_06744_),
    .B(_06745_),
    .C_N(_06747_),
    .X(_06748_));
 sky130_fd_sc_hd__xor2_2 _15268_ (.A(_06746_),
    .B(_06747_),
    .X(_06749_));
 sky130_fd_sc_hd__or2_1 _15269_ (.A(_06740_),
    .B(_06749_),
    .X(_06750_));
 sky130_fd_sc_hd__xor2_2 _15270_ (.A(_06740_),
    .B(_06749_),
    .X(_06751_));
 sky130_fd_sc_hd__or2_2 _15271_ (.A(_06612_),
    .B(_06614_),
    .X(_06752_));
 sky130_fd_sc_hd__o2bb2a_2 _15272_ (.A1_N(net467),
    .A2_N(_06573_),
    .B1(_06574_),
    .B2(_06575_),
    .X(_06753_));
 sky130_fd_sc_hd__a22oi_1 _15273_ (.A1(net378),
    .A2(net480),
    .B1(net476),
    .B2(net384),
    .Y(_06754_));
 sky130_fd_sc_hd__and4_1 _15274_ (.A(net384),
    .B(net378),
    .C(net480),
    .D(net476),
    .X(_06755_));
 sky130_fd_sc_hd__o2bb2a_1 _15275_ (.A1_N(net373),
    .A2_N(net485),
    .B1(_06754_),
    .B2(_06755_),
    .X(_06756_));
 sky130_fd_sc_hd__and4bb_1 _15276_ (.A_N(_06754_),
    .B_N(_06755_),
    .C(net372),
    .D(net485),
    .X(_06757_));
 sky130_fd_sc_hd__or2_2 _15277_ (.A(_06756_),
    .B(_06757_),
    .X(_06758_));
 sky130_fd_sc_hd__or2_1 _15278_ (.A(_06753_),
    .B(_06758_),
    .X(_06759_));
 sky130_fd_sc_hd__xor2_2 _15279_ (.A(_06753_),
    .B(_06758_),
    .X(_06760_));
 sky130_fd_sc_hd__nand2_1 _15280_ (.A(_06752_),
    .B(_06760_),
    .Y(_06761_));
 sky130_fd_sc_hd__xnor2_2 _15281_ (.A(_06752_),
    .B(_06760_),
    .Y(_06762_));
 sky130_fd_sc_hd__nand2_2 _15282_ (.A(_06615_),
    .B(_06617_),
    .Y(_06763_));
 sky130_fd_sc_hd__nand2b_1 _15283_ (.A_N(_06762_),
    .B(_06763_),
    .Y(_06764_));
 sky130_fd_sc_hd__xnor2_2 _15284_ (.A(_06762_),
    .B(_06763_),
    .Y(_06765_));
 sky130_fd_sc_hd__nand2_1 _15285_ (.A(_06751_),
    .B(_06765_),
    .Y(_06766_));
 sky130_fd_sc_hd__xor2_2 _15286_ (.A(_06751_),
    .B(_06765_),
    .X(_06767_));
 sky130_fd_sc_hd__nand2b_2 _15287_ (.A_N(_06735_),
    .B(_06767_),
    .Y(_06768_));
 sky130_fd_sc_hd__xnor2_1 _15288_ (.A(_06735_),
    .B(_06767_),
    .Y(_06769_));
 sky130_fd_sc_hd__nand2b_2 _15289_ (.A_N(_06734_),
    .B(_06769_),
    .Y(_06770_));
 sky130_fd_sc_hd__xnor2_1 _15290_ (.A(_06734_),
    .B(_06769_),
    .Y(_06771_));
 sky130_fd_sc_hd__nand2_2 _15291_ (.A(_06733_),
    .B(_06771_),
    .Y(_06772_));
 sky130_fd_sc_hd__or2_1 _15292_ (.A(_06733_),
    .B(_06771_),
    .X(_06773_));
 sky130_fd_sc_hd__o211a_2 _15293_ (.A1(_06592_),
    .A2(_06628_),
    .B1(_06772_),
    .C1(_06773_),
    .X(_06774_));
 sky130_fd_sc_hd__a211oi_1 _15294_ (.A1(_06772_),
    .A2(_06773_),
    .B1(_06592_),
    .C1(_06628_),
    .Y(_06775_));
 sky130_fd_sc_hd__or2_2 _15295_ (.A(_06774_),
    .B(_06775_),
    .X(_06776_));
 sky130_fd_sc_hd__or2_1 _15296_ (.A(_06665_),
    .B(_06667_),
    .X(_06777_));
 sky130_fd_sc_hd__inv_2 _15297_ (.A(_06777_),
    .Y(_06778_));
 sky130_fd_sc_hd__nand2_2 _15298_ (.A(_06624_),
    .B(_06626_),
    .Y(_06779_));
 sky130_fd_sc_hd__a22o_1 _15299_ (.A1(net528),
    .A2(net334),
    .B1(net331),
    .B2(net533),
    .X(_06780_));
 sky130_fd_sc_hd__and4_1 _15300_ (.A(net528),
    .B(net533),
    .C(net334),
    .D(net331),
    .X(_06781_));
 sky130_fd_sc_hd__inv_2 _15301_ (.A(_06781_),
    .Y(_06782_));
 sky130_fd_sc_hd__a22oi_1 _15302_ (.A1(net539),
    .A2(net329),
    .B1(_06780_),
    .B2(_06782_),
    .Y(_06783_));
 sky130_fd_sc_hd__and4_1 _15303_ (.A(net539),
    .B(net329),
    .C(_06780_),
    .D(_06782_),
    .X(_06784_));
 sky130_fd_sc_hd__or2_1 _15304_ (.A(_06783_),
    .B(_06784_),
    .X(_06785_));
 sky130_fd_sc_hd__or2_1 _15305_ (.A(_06635_),
    .B(_06637_),
    .X(_06786_));
 sky130_fd_sc_hd__or3b_1 _15306_ (.A(_06783_),
    .B(_06784_),
    .C_N(_06786_),
    .X(_06787_));
 sky130_fd_sc_hd__xor2_2 _15307_ (.A(_06785_),
    .B(_06786_),
    .X(_06788_));
 sky130_fd_sc_hd__and4b_2 _15308_ (.A_N(\mul0.a[8] ),
    .B(net327),
    .C(net326),
    .D(\mul0.a[9] ),
    .X(_06789_));
 sky130_fd_sc_hd__o2bb2a_1 _15309_ (.A1_N(\mul0.a[9] ),
    .A2_N(net327),
    .B1(net57),
    .B2(net547),
    .X(_06790_));
 sky130_fd_sc_hd__nor2_1 _15310_ (.A(_06789_),
    .B(_06790_),
    .Y(_06791_));
 sky130_fd_sc_hd__xnor2_1 _15311_ (.A(_06788_),
    .B(_06791_),
    .Y(_06792_));
 sky130_fd_sc_hd__o31ai_2 _15312_ (.A1(_06638_),
    .A2(_06641_),
    .A3(_06643_),
    .B1(_06639_),
    .Y(_06793_));
 sky130_fd_sc_hd__nand2_1 _15313_ (.A(_06792_),
    .B(_06793_),
    .Y(_06794_));
 sky130_fd_sc_hd__xnor2_1 _15314_ (.A(_06792_),
    .B(_06793_),
    .Y(_06795_));
 sky130_fd_sc_hd__xnor2_1 _15315_ (.A(_06642_),
    .B(_06795_),
    .Y(_06796_));
 sky130_fd_sc_hd__or2_1 _15316_ (.A(_06654_),
    .B(_06656_),
    .X(_06797_));
 sky130_fd_sc_hd__a31oi_4 _15317_ (.A1(net513),
    .A2(net349),
    .A3(_06593_),
    .B1(_06594_),
    .Y(_06798_));
 sky130_fd_sc_hd__a22oi_1 _15318_ (.A1(net513),
    .A2(net346),
    .B1(net342),
    .B2(net518),
    .Y(_06799_));
 sky130_fd_sc_hd__and4_1 _15319_ (.A(net513),
    .B(net518),
    .C(net346),
    .D(net342),
    .X(_06800_));
 sky130_fd_sc_hd__o2bb2a_1 _15320_ (.A1_N(net522),
    .A2_N(net338),
    .B1(_06799_),
    .B2(_06800_),
    .X(_06801_));
 sky130_fd_sc_hd__and4bb_1 _15321_ (.A_N(_06799_),
    .B_N(_06800_),
    .C(net522),
    .D(net338),
    .X(_06802_));
 sky130_fd_sc_hd__or2_1 _15322_ (.A(_06801_),
    .B(_06802_),
    .X(_06803_));
 sky130_fd_sc_hd__or2_1 _15323_ (.A(_06798_),
    .B(_06803_),
    .X(_06804_));
 sky130_fd_sc_hd__xor2_2 _15324_ (.A(_06798_),
    .B(_06803_),
    .X(_06805_));
 sky130_fd_sc_hd__nand2_1 _15325_ (.A(_06797_),
    .B(_06805_),
    .Y(_06806_));
 sky130_fd_sc_hd__xnor2_2 _15326_ (.A(_06797_),
    .B(_06805_),
    .Y(_06807_));
 sky130_fd_sc_hd__a21oi_4 _15327_ (.A1(_06604_),
    .A2(_06607_),
    .B1(_06807_),
    .Y(_06808_));
 sky130_fd_sc_hd__and3_1 _15328_ (.A(_06604_),
    .B(_06607_),
    .C(_06807_),
    .X(_06809_));
 sky130_fd_sc_hd__a211oi_4 _15329_ (.A1(_06657_),
    .A2(_06659_),
    .B1(_06808_),
    .C1(_06809_),
    .Y(_06810_));
 sky130_fd_sc_hd__o211a_1 _15330_ (.A1(_06808_),
    .A2(_06809_),
    .B1(_06657_),
    .C1(_06659_),
    .X(_06811_));
 sky130_fd_sc_hd__and2b_1 _15331_ (.A_N(_06661_),
    .B(_06663_),
    .X(_06812_));
 sky130_fd_sc_hd__nor3_1 _15332_ (.A(_06810_),
    .B(_06811_),
    .C(_06812_),
    .Y(_06813_));
 sky130_fd_sc_hd__o21a_1 _15333_ (.A1(_06810_),
    .A2(_06811_),
    .B1(_06812_),
    .X(_06814_));
 sky130_fd_sc_hd__or3_1 _15334_ (.A(_06796_),
    .B(_06813_),
    .C(_06814_),
    .X(_06815_));
 sky130_fd_sc_hd__o21ai_1 _15335_ (.A1(_06813_),
    .A2(_06814_),
    .B1(_06796_),
    .Y(_06816_));
 sky130_fd_sc_hd__and3_2 _15336_ (.A(_06779_),
    .B(_06815_),
    .C(_06816_),
    .X(_06817_));
 sky130_fd_sc_hd__a21oi_1 _15337_ (.A1(_06815_),
    .A2(_06816_),
    .B1(_06779_),
    .Y(_06818_));
 sky130_fd_sc_hd__nor3_2 _15338_ (.A(_06778_),
    .B(_06817_),
    .C(_06818_),
    .Y(_06819_));
 sky130_fd_sc_hd__o21a_1 _15339_ (.A1(_06817_),
    .A2(_06818_),
    .B1(_06778_),
    .X(_06820_));
 sky130_fd_sc_hd__nor2_2 _15340_ (.A(_06819_),
    .B(_06820_),
    .Y(_06821_));
 sky130_fd_sc_hd__and2b_1 _15341_ (.A_N(_06776_),
    .B(_06821_),
    .X(_06822_));
 sky130_fd_sc_hd__xnor2_4 _15342_ (.A(_06776_),
    .B(_06821_),
    .Y(_06823_));
 sky130_fd_sc_hd__a21oi_4 _15343_ (.A1(_06633_),
    .A2(_06673_),
    .B1(_06631_),
    .Y(_06824_));
 sky130_fd_sc_hd__and2b_1 _15344_ (.A_N(_06824_),
    .B(_06823_),
    .X(_06825_));
 sky130_fd_sc_hd__xnor2_4 _15345_ (.A(_06823_),
    .B(_06824_),
    .Y(_06826_));
 sky130_fd_sc_hd__or2_2 _15346_ (.A(_06669_),
    .B(_06671_),
    .X(_06827_));
 sky130_fd_sc_hd__xnor2_4 _15347_ (.A(_06826_),
    .B(_06827_),
    .Y(_06828_));
 sky130_fd_sc_hd__a21o_1 _15348_ (.A1(_06556_),
    .A2(_06677_),
    .B1(_06676_),
    .X(_06829_));
 sky130_fd_sc_hd__and2b_1 _15349_ (.A_N(_06828_),
    .B(_06829_),
    .X(_06830_));
 sky130_fd_sc_hd__xnor2_4 _15350_ (.A(_06828_),
    .B(_06829_),
    .Y(_06831_));
 sky130_fd_sc_hd__xnor2_4 _15351_ (.A(_06695_),
    .B(_06831_),
    .Y(_06832_));
 sky130_fd_sc_hd__nand2b_1 _15352_ (.A_N(_06694_),
    .B(_06832_),
    .Y(_06833_));
 sky130_fd_sc_hd__and2b_1 _15353_ (.A_N(_06832_),
    .B(_06694_),
    .X(_06834_));
 sky130_fd_sc_hd__xor2_4 _15354_ (.A(_06694_),
    .B(_06832_),
    .X(_06835_));
 sky130_fd_sc_hd__o21ba_1 _15355_ (.A1(_06686_),
    .A2(_06690_),
    .B1_N(_06684_),
    .X(_06836_));
 sky130_fd_sc_hd__xor2_4 _15356_ (.A(_06835_),
    .B(_06836_),
    .X(_06837_));
 sky130_fd_sc_hd__a22o_1 _15357_ (.A1(\state[4] ),
    .A2(\temp[22] ),
    .B1(_02690_),
    .B2(net5),
    .X(_06838_));
 sky130_fd_sc_hd__a21o_1 _15358_ (.A1(_03058_),
    .A2(_06837_),
    .B1(_06838_),
    .X(_06839_));
 sky130_fd_sc_hd__mux2_1 _15359_ (.A0(net755),
    .A1(_06839_),
    .S(net4),
    .X(_00289_));
 sky130_fd_sc_hd__a21o_1 _15360_ (.A1(_06458_),
    .A2(_06702_),
    .B1(_06454_),
    .X(_06840_));
 sky130_fd_sc_hd__nand2_2 _15361_ (.A(_06558_),
    .B(_06698_),
    .Y(_06841_));
 sky130_fd_sc_hd__xnor2_2 _15362_ (.A(_06701_),
    .B(_06841_),
    .Y(_06842_));
 sky130_fd_sc_hd__xor2_1 _15363_ (.A(_06458_),
    .B(_06842_),
    .X(_06843_));
 sky130_fd_sc_hd__inv_2 _15364_ (.A(_06843_),
    .Y(_06844_));
 sky130_fd_sc_hd__xnor2_1 _15365_ (.A(_06840_),
    .B(_06843_),
    .Y(_06845_));
 sky130_fd_sc_hd__a21o_1 _15366_ (.A1(_06696_),
    .A2(_06700_),
    .B1(_06699_),
    .X(_06846_));
 sky130_fd_sc_hd__a22o_1 _15367_ (.A1(net393),
    .A2(net464),
    .B1(net461),
    .B2(net398),
    .X(_06847_));
 sky130_fd_sc_hd__nand4_2 _15368_ (.A(net398),
    .B(net393),
    .C(net464),
    .D(net461),
    .Y(_06848_));
 sky130_fd_sc_hd__a22o_1 _15369_ (.A1(net388),
    .A2(net466),
    .B1(_06847_),
    .B2(_06848_),
    .X(_06849_));
 sky130_fd_sc_hd__nand4_2 _15370_ (.A(net388),
    .B(net466),
    .C(_06847_),
    .D(_06848_),
    .Y(_06850_));
 sky130_fd_sc_hd__nand2_2 _15371_ (.A(_06849_),
    .B(_06850_),
    .Y(_06851_));
 sky130_fd_sc_hd__a22oi_1 _15372_ (.A1(net406),
    .A2(net455),
    .B1(net454),
    .B2(net410),
    .Y(_06852_));
 sky130_fd_sc_hd__and4_1 _15373_ (.A(net410),
    .B(net406),
    .C(net455),
    .D(net454),
    .X(_06853_));
 sky130_fd_sc_hd__nor2_2 _15374_ (.A(_06852_),
    .B(_06853_),
    .Y(_06854_));
 sky130_fd_sc_hd__nand2_2 _15375_ (.A(net402),
    .B(net458),
    .Y(_06855_));
 sky130_fd_sc_hd__xor2_4 _15376_ (.A(_06854_),
    .B(_06855_),
    .X(_06856_));
 sky130_fd_sc_hd__nor2_2 _15377_ (.A(_06715_),
    .B(_06717_),
    .Y(_06857_));
 sky130_fd_sc_hd__nor2_1 _15378_ (.A(_06856_),
    .B(_06857_),
    .Y(_06858_));
 sky130_fd_sc_hd__xnor2_4 _15379_ (.A(_06856_),
    .B(_06857_),
    .Y(_06859_));
 sky130_fd_sc_hd__xor2_2 _15380_ (.A(_06851_),
    .B(_06859_),
    .X(_06860_));
 sky130_fd_sc_hd__nand2_2 _15381_ (.A(_06846_),
    .B(_06860_),
    .Y(_06861_));
 sky130_fd_sc_hd__xnor2_1 _15382_ (.A(_06846_),
    .B(_06860_),
    .Y(_06862_));
 sky130_fd_sc_hd__a21o_2 _15383_ (.A1(_06720_),
    .A2(_06722_),
    .B1(_06862_),
    .X(_06863_));
 sky130_fd_sc_hd__nand3_1 _15384_ (.A(_06720_),
    .B(_06722_),
    .C(_06862_),
    .Y(_06864_));
 sky130_fd_sc_hd__a21oi_2 _15385_ (.A1(_06863_),
    .A2(_06864_),
    .B1(_06845_),
    .Y(_06865_));
 sky130_fd_sc_hd__and3_1 _15386_ (.A(_06845_),
    .B(_06863_),
    .C(_06864_),
    .X(_06866_));
 sky130_fd_sc_hd__o211a_2 _15387_ (.A1(_06865_),
    .A2(_06866_),
    .B1(_06705_),
    .C1(_06729_),
    .X(_06867_));
 sky130_fd_sc_hd__a211oi_4 _15388_ (.A1(_06705_),
    .A2(_06729_),
    .B1(_06865_),
    .C1(_06866_),
    .Y(_06868_));
 sky130_fd_sc_hd__a22o_1 _15389_ (.A1(net496),
    .A2(net358),
    .B1(net353),
    .B2(net501),
    .X(_06869_));
 sky130_fd_sc_hd__nand4_2 _15390_ (.A(net501),
    .B(net496),
    .C(net358),
    .D(net353),
    .Y(_06870_));
 sky130_fd_sc_hd__a22o_1 _15391_ (.A1(net505),
    .A2(net350),
    .B1(_06869_),
    .B2(_06870_),
    .X(_06871_));
 sky130_fd_sc_hd__nand4_1 _15392_ (.A(net505),
    .B(net350),
    .C(_06869_),
    .D(_06870_),
    .Y(_06872_));
 sky130_fd_sc_hd__nand2_1 _15393_ (.A(_06871_),
    .B(_06872_),
    .Y(_06873_));
 sky130_fd_sc_hd__a22o_1 _15394_ (.A1(net368),
    .A2(net489),
    .B1(net485),
    .B2(net634),
    .X(_06874_));
 sky130_fd_sc_hd__and4_1 _15395_ (.A(net634),
    .B(net368),
    .C(net489),
    .D(net485),
    .X(_06875_));
 sky130_fd_sc_hd__inv_2 _15396_ (.A(_06875_),
    .Y(_06876_));
 sky130_fd_sc_hd__a22oi_1 _15397_ (.A1(net492),
    .A2(net362),
    .B1(_06874_),
    .B2(_06876_),
    .Y(_06877_));
 sky130_fd_sc_hd__and4_1 _15398_ (.A(net492),
    .B(net362),
    .C(_06874_),
    .D(_06876_),
    .X(_06878_));
 sky130_fd_sc_hd__or2_1 _15399_ (.A(_06877_),
    .B(_06878_),
    .X(_06879_));
 sky130_fd_sc_hd__or2_1 _15400_ (.A(_06742_),
    .B(_06745_),
    .X(_06880_));
 sky130_fd_sc_hd__nand2b_2 _15401_ (.A_N(_06879_),
    .B(_06880_),
    .Y(_06881_));
 sky130_fd_sc_hd__xor2_1 _15402_ (.A(_06879_),
    .B(_06880_),
    .X(_06882_));
 sky130_fd_sc_hd__or2_2 _15403_ (.A(_06873_),
    .B(_06882_),
    .X(_06883_));
 sky130_fd_sc_hd__nand2_1 _15404_ (.A(_06873_),
    .B(_06882_),
    .Y(_06884_));
 sky130_fd_sc_hd__and2_1 _15405_ (.A(_06883_),
    .B(_06884_),
    .X(_06885_));
 sky130_fd_sc_hd__or2_1 _15406_ (.A(_06755_),
    .B(_06757_),
    .X(_06886_));
 sky130_fd_sc_hd__nand2_2 _15407_ (.A(_06710_),
    .B(_06712_),
    .Y(_06887_));
 sky130_fd_sc_hd__a22o_1 _15408_ (.A1(net378),
    .A2(net476),
    .B1(net471),
    .B2(net384),
    .X(_06888_));
 sky130_fd_sc_hd__inv_2 _15409_ (.A(_06888_),
    .Y(_06889_));
 sky130_fd_sc_hd__and4_1 _15410_ (.A(net384),
    .B(net378),
    .C(net476),
    .D(net471),
    .X(_06890_));
 sky130_fd_sc_hd__o2bb2a_1 _15411_ (.A1_N(net372),
    .A2_N(net480),
    .B1(_06889_),
    .B2(_06890_),
    .X(_06891_));
 sky130_fd_sc_hd__and4b_1 _15412_ (.A_N(_06890_),
    .B(net480),
    .C(net373),
    .D(_06888_),
    .X(_06892_));
 sky130_fd_sc_hd__or2_1 _15413_ (.A(_06891_),
    .B(_06892_),
    .X(_06893_));
 sky130_fd_sc_hd__nand2b_1 _15414_ (.A_N(_06893_),
    .B(_06887_),
    .Y(_06894_));
 sky130_fd_sc_hd__xnor2_1 _15415_ (.A(_06887_),
    .B(_06893_),
    .Y(_06895_));
 sky130_fd_sc_hd__nand2_1 _15416_ (.A(_06886_),
    .B(_06895_),
    .Y(_06896_));
 sky130_fd_sc_hd__xnor2_1 _15417_ (.A(_06886_),
    .B(_06895_),
    .Y(_06897_));
 sky130_fd_sc_hd__a21o_2 _15418_ (.A1(_06759_),
    .A2(_06761_),
    .B1(_06897_),
    .X(_06898_));
 sky130_fd_sc_hd__nand3_1 _15419_ (.A(_06759_),
    .B(_06761_),
    .C(_06897_),
    .Y(_06899_));
 sky130_fd_sc_hd__nand3_2 _15420_ (.A(_06885_),
    .B(_06898_),
    .C(_06899_),
    .Y(_06900_));
 sky130_fd_sc_hd__a21o_1 _15421_ (.A1(_06898_),
    .A2(_06899_),
    .B1(_06885_),
    .X(_06901_));
 sky130_fd_sc_hd__o211a_2 _15422_ (.A1(_06724_),
    .A2(_06727_),
    .B1(_06900_),
    .C1(_06901_),
    .X(_06902_));
 sky130_fd_sc_hd__a211oi_2 _15423_ (.A1(_06900_),
    .A2(_06901_),
    .B1(_06724_),
    .C1(_06727_),
    .Y(_06903_));
 sky130_fd_sc_hd__a211oi_4 _15424_ (.A1(_06764_),
    .A2(_06766_),
    .B1(_06902_),
    .C1(_06903_),
    .Y(_06904_));
 sky130_fd_sc_hd__o211a_1 _15425_ (.A1(_06902_),
    .A2(_06903_),
    .B1(_06764_),
    .C1(_06766_),
    .X(_06905_));
 sky130_fd_sc_hd__nor4_4 _15426_ (.A(_06867_),
    .B(_06868_),
    .C(_06904_),
    .D(_06905_),
    .Y(_06906_));
 sky130_fd_sc_hd__o22a_1 _15427_ (.A1(_06867_),
    .A2(_06868_),
    .B1(_06904_),
    .B2(_06905_),
    .X(_06907_));
 sky130_fd_sc_hd__a211o_2 _15428_ (.A1(_06732_),
    .A2(_06772_),
    .B1(_06906_),
    .C1(_06907_),
    .X(_06908_));
 sky130_fd_sc_hd__o211ai_4 _15429_ (.A1(_06906_),
    .A2(_06907_),
    .B1(_06732_),
    .C1(_06772_),
    .Y(_06909_));
 sky130_fd_sc_hd__nand2b_2 _15430_ (.A_N(_06813_),
    .B(_06815_),
    .Y(_06910_));
 sky130_fd_sc_hd__a22o_1 _15431_ (.A1(net523),
    .A2(net334),
    .B1(net331),
    .B2(net528),
    .X(_06911_));
 sky130_fd_sc_hd__and4_1 _15432_ (.A(net522),
    .B(net528),
    .C(net334),
    .D(net331),
    .X(_06912_));
 sky130_fd_sc_hd__inv_2 _15433_ (.A(_06912_),
    .Y(_06913_));
 sky130_fd_sc_hd__a22oi_1 _15434_ (.A1(net533),
    .A2(net329),
    .B1(_06911_),
    .B2(_06913_),
    .Y(_06914_));
 sky130_fd_sc_hd__and4_1 _15435_ (.A(net533),
    .B(net329),
    .C(_06911_),
    .D(_06913_),
    .X(_06915_));
 sky130_fd_sc_hd__or2_2 _15436_ (.A(_06914_),
    .B(_06915_),
    .X(_06916_));
 sky130_fd_sc_hd__nor2_2 _15437_ (.A(_06781_),
    .B(_06784_),
    .Y(_06917_));
 sky130_fd_sc_hd__xnor2_2 _15438_ (.A(_06916_),
    .B(_06917_),
    .Y(_06918_));
 sky130_fd_sc_hd__and4b_2 _15439_ (.A_N(\mul0.a[9] ),
    .B(net327),
    .C(net326),
    .D(net539),
    .X(_06919_));
 sky130_fd_sc_hd__inv_2 _15440_ (.A(_06919_),
    .Y(_06920_));
 sky130_fd_sc_hd__o2bb2a_1 _15441_ (.A1_N(net539),
    .A2_N(net328),
    .B1(net57),
    .B2(\mul0.a[9] ),
    .X(_06921_));
 sky130_fd_sc_hd__nor2_1 _15442_ (.A(_06919_),
    .B(_06921_),
    .Y(_06922_));
 sky130_fd_sc_hd__xnor2_2 _15443_ (.A(_06918_),
    .B(_06922_),
    .Y(_06923_));
 sky130_fd_sc_hd__o31ai_2 _15444_ (.A1(_06788_),
    .A2(_06789_),
    .A3(_06790_),
    .B1(_06787_),
    .Y(_06924_));
 sky130_fd_sc_hd__nand2_1 _15445_ (.A(_06923_),
    .B(_06924_),
    .Y(_06925_));
 sky130_fd_sc_hd__xnor2_2 _15446_ (.A(_06923_),
    .B(_06924_),
    .Y(_06926_));
 sky130_fd_sc_hd__inv_2 _15447_ (.A(_06926_),
    .Y(_06927_));
 sky130_fd_sc_hd__nand2_1 _15448_ (.A(_06789_),
    .B(_06927_),
    .Y(_06928_));
 sky130_fd_sc_hd__xor2_2 _15449_ (.A(_06789_),
    .B(_06926_),
    .X(_06929_));
 sky130_fd_sc_hd__or2_1 _15450_ (.A(_06800_),
    .B(_06802_),
    .X(_06930_));
 sky130_fd_sc_hd__nand2_1 _15451_ (.A(_06737_),
    .B(_06739_),
    .Y(_06931_));
 sky130_fd_sc_hd__a22o_1 _15452_ (.A1(net509),
    .A2(net346),
    .B1(net342),
    .B2(net513),
    .X(_06932_));
 sky130_fd_sc_hd__inv_2 _15453_ (.A(_06932_),
    .Y(_06933_));
 sky130_fd_sc_hd__and4_1 _15454_ (.A(net509),
    .B(net514),
    .C(net346),
    .D(net342),
    .X(_06934_));
 sky130_fd_sc_hd__o2bb2a_1 _15455_ (.A1_N(net518),
    .A2_N(net338),
    .B1(_06933_),
    .B2(_06934_),
    .X(_06935_));
 sky130_fd_sc_hd__and4b_1 _15456_ (.A_N(_06934_),
    .B(net338),
    .C(net518),
    .D(_06932_),
    .X(_06936_));
 sky130_fd_sc_hd__or2_1 _15457_ (.A(_06935_),
    .B(_06936_),
    .X(_06937_));
 sky130_fd_sc_hd__nand2b_1 _15458_ (.A_N(_06937_),
    .B(_06931_),
    .Y(_06938_));
 sky130_fd_sc_hd__xnor2_1 _15459_ (.A(_06931_),
    .B(_06937_),
    .Y(_06939_));
 sky130_fd_sc_hd__nand2_1 _15460_ (.A(_06930_),
    .B(_06939_),
    .Y(_06940_));
 sky130_fd_sc_hd__xnor2_1 _15461_ (.A(_06930_),
    .B(_06939_),
    .Y(_06941_));
 sky130_fd_sc_hd__a21oi_1 _15462_ (.A1(_06748_),
    .A2(_06750_),
    .B1(_06941_),
    .Y(_06942_));
 sky130_fd_sc_hd__a21o_1 _15463_ (.A1(_06748_),
    .A2(_06750_),
    .B1(_06941_),
    .X(_06943_));
 sky130_fd_sc_hd__and3_1 _15464_ (.A(_06748_),
    .B(_06750_),
    .C(_06941_),
    .X(_06944_));
 sky130_fd_sc_hd__a211o_2 _15465_ (.A1(_06804_),
    .A2(_06806_),
    .B1(_06942_),
    .C1(_06944_),
    .X(_06945_));
 sky130_fd_sc_hd__o211ai_2 _15466_ (.A1(_06942_),
    .A2(_06944_),
    .B1(_06804_),
    .C1(_06806_),
    .Y(_06946_));
 sky130_fd_sc_hd__o211a_2 _15467_ (.A1(_06808_),
    .A2(_06810_),
    .B1(_06945_),
    .C1(_06946_),
    .X(_06947_));
 sky130_fd_sc_hd__a211oi_2 _15468_ (.A1(_06945_),
    .A2(_06946_),
    .B1(_06808_),
    .C1(_06810_),
    .Y(_06948_));
 sky130_fd_sc_hd__nor3_2 _15469_ (.A(_06929_),
    .B(_06947_),
    .C(_06948_),
    .Y(_06949_));
 sky130_fd_sc_hd__o21a_1 _15470_ (.A1(_06947_),
    .A2(_06948_),
    .B1(_06929_),
    .X(_06950_));
 sky130_fd_sc_hd__a211o_2 _15471_ (.A1(_06768_),
    .A2(_06770_),
    .B1(_06949_),
    .C1(_06950_),
    .X(_06951_));
 sky130_fd_sc_hd__o211ai_4 _15472_ (.A1(_06949_),
    .A2(_06950_),
    .B1(_06768_),
    .C1(_06770_),
    .Y(_06952_));
 sky130_fd_sc_hd__nand3_4 _15473_ (.A(_06910_),
    .B(_06951_),
    .C(_06952_),
    .Y(_06953_));
 sky130_fd_sc_hd__a21o_1 _15474_ (.A1(_06951_),
    .A2(_06952_),
    .B1(_06910_),
    .X(_06954_));
 sky130_fd_sc_hd__nand4_4 _15475_ (.A(_06908_),
    .B(_06909_),
    .C(_06953_),
    .D(_06954_),
    .Y(_06955_));
 sky130_fd_sc_hd__a22o_1 _15476_ (.A1(_06908_),
    .A2(_06909_),
    .B1(_06953_),
    .B2(_06954_),
    .X(_06956_));
 sky130_fd_sc_hd__o211ai_4 _15477_ (.A1(_06774_),
    .A2(_06822_),
    .B1(_06955_),
    .C1(_06956_),
    .Y(_06957_));
 sky130_fd_sc_hd__a211o_1 _15478_ (.A1(_06955_),
    .A2(_06956_),
    .B1(_06774_),
    .C1(_06822_),
    .X(_06958_));
 sky130_fd_sc_hd__o211ai_4 _15479_ (.A1(_06817_),
    .A2(_06819_),
    .B1(_06957_),
    .C1(_06958_),
    .Y(_06959_));
 sky130_fd_sc_hd__a211o_1 _15480_ (.A1(_06957_),
    .A2(_06958_),
    .B1(_06817_),
    .C1(_06819_),
    .X(_06960_));
 sky130_fd_sc_hd__and2_1 _15481_ (.A(_06959_),
    .B(_06960_),
    .X(_06961_));
 sky130_fd_sc_hd__a21oi_1 _15482_ (.A1(_06826_),
    .A2(_06827_),
    .B1(_06825_),
    .Y(_06962_));
 sky130_fd_sc_hd__nand2b_1 _15483_ (.A_N(_06962_),
    .B(_06961_),
    .Y(_06963_));
 sky130_fd_sc_hd__xnor2_1 _15484_ (.A(_06961_),
    .B(_06962_),
    .Y(_06964_));
 sky130_fd_sc_hd__o21ai_1 _15485_ (.A1(_06642_),
    .A2(_06795_),
    .B1(_06794_),
    .Y(_06965_));
 sky130_fd_sc_hd__nand2_1 _15486_ (.A(_06964_),
    .B(_06965_),
    .Y(_06966_));
 sky130_fd_sc_hd__xnor2_1 _15487_ (.A(_06964_),
    .B(_06965_),
    .Y(_06967_));
 sky130_fd_sc_hd__a21oi_1 _15488_ (.A1(_06695_),
    .A2(_06831_),
    .B1(_06830_),
    .Y(_06968_));
 sky130_fd_sc_hd__nor2_1 _15489_ (.A(_06967_),
    .B(_06968_),
    .Y(_06969_));
 sky130_fd_sc_hd__and2_1 _15490_ (.A(_06967_),
    .B(_06968_),
    .X(_06970_));
 sky130_fd_sc_hd__or2_1 _15491_ (.A(_06969_),
    .B(_06970_),
    .X(_06971_));
 sky130_fd_sc_hd__nor2_1 _15492_ (.A(_06686_),
    .B(_06835_),
    .Y(_06972_));
 sky130_fd_sc_hd__a2111o_1 _15493_ (.A1(_06398_),
    .A2(_06399_),
    .B1(_06686_),
    .C1(_06689_),
    .D1(_06835_),
    .X(_06973_));
 sky130_fd_sc_hd__a221oi_2 _15494_ (.A1(_06684_),
    .A2(_06833_),
    .B1(_06972_),
    .B2(_06687_),
    .C1(_06834_),
    .Y(_06974_));
 sky130_fd_sc_hd__a21oi_1 _15495_ (.A1(_06973_),
    .A2(_06974_),
    .B1(_06971_),
    .Y(_06975_));
 sky130_fd_sc_hd__and3_1 _15496_ (.A(_06971_),
    .B(_06973_),
    .C(_06974_),
    .X(_06976_));
 sky130_fd_sc_hd__nor2_2 _15497_ (.A(_06975_),
    .B(_06976_),
    .Y(_06977_));
 sky130_fd_sc_hd__a22o_1 _15498_ (.A1(\state[4] ),
    .A2(net741),
    .B1(_02696_),
    .B2(net5),
    .X(_06978_));
 sky130_fd_sc_hd__a21o_1 _15499_ (.A1(_03058_),
    .A2(_06977_),
    .B1(_06978_),
    .X(_06979_));
 sky130_fd_sc_hd__mux2_1 _15500_ (.A0(net725),
    .A1(_06979_),
    .S(net4),
    .X(_00290_));
 sky130_fd_sc_hd__nor2_4 _15501_ (.A(_06455_),
    .B(_06842_),
    .Y(_06980_));
 sky130_fd_sc_hd__and2_1 _15502_ (.A(_06456_),
    .B(_06842_),
    .X(_06981_));
 sky130_fd_sc_hd__nor2_2 _15503_ (.A(_06980_),
    .B(_06981_),
    .Y(_06982_));
 sky130_fd_sc_hd__or2_4 _15504_ (.A(_06980_),
    .B(_06981_),
    .X(_06983_));
 sky130_fd_sc_hd__o21bai_4 _15505_ (.A1(_06851_),
    .A2(_06859_),
    .B1_N(_06858_),
    .Y(_06984_));
 sky130_fd_sc_hd__a21o_4 _15506_ (.A1(_06700_),
    .A2(_06841_),
    .B1(_06699_),
    .X(_06985_));
 sky130_fd_sc_hd__a22o_1 _15507_ (.A1(net393),
    .A2(net462),
    .B1(net458),
    .B2(net398),
    .X(_06986_));
 sky130_fd_sc_hd__nand4_2 _15508_ (.A(net398),
    .B(net393),
    .C(net462),
    .D(net458),
    .Y(_06987_));
 sky130_fd_sc_hd__a22o_1 _15509_ (.A1(net388),
    .A2(net465),
    .B1(_06986_),
    .B2(_06987_),
    .X(_06988_));
 sky130_fd_sc_hd__nand4_2 _15510_ (.A(net388),
    .B(net464),
    .C(_06986_),
    .D(_06987_),
    .Y(_06989_));
 sky130_fd_sc_hd__nand2_1 _15511_ (.A(_06988_),
    .B(_06989_),
    .Y(_06990_));
 sky130_fd_sc_hd__a31o_1 _15512_ (.A1(net402),
    .A2(net458),
    .A3(_06854_),
    .B1(_06853_),
    .X(_06991_));
 sky130_fd_sc_hd__nand2_1 _15513_ (.A(net403),
    .B(net455),
    .Y(_06992_));
 sky130_fd_sc_hd__and3_1 _15514_ (.A(net411),
    .B(net407),
    .C(net453),
    .X(_06993_));
 sky130_fd_sc_hd__o21a_1 _15515_ (.A1(net411),
    .A2(net407),
    .B1(net453),
    .X(_06994_));
 sky130_fd_sc_hd__and2b_1 _15516_ (.A_N(_06993_),
    .B(_06994_),
    .X(_06995_));
 sky130_fd_sc_hd__xnor2_2 _15517_ (.A(_06992_),
    .B(_06995_),
    .Y(_06996_));
 sky130_fd_sc_hd__xor2_2 _15518_ (.A(_06991_),
    .B(_06996_),
    .X(_06997_));
 sky130_fd_sc_hd__xnor2_2 _15519_ (.A(_06990_),
    .B(_06997_),
    .Y(_06998_));
 sky130_fd_sc_hd__and2_1 _15520_ (.A(_06985_),
    .B(_06998_),
    .X(_06999_));
 sky130_fd_sc_hd__xnor2_1 _15521_ (.A(_06985_),
    .B(_06998_),
    .Y(_07000_));
 sky130_fd_sc_hd__and2b_1 _15522_ (.A_N(_07000_),
    .B(_06984_),
    .X(_07001_));
 sky130_fd_sc_hd__xor2_1 _15523_ (.A(_06984_),
    .B(_07000_),
    .X(_07002_));
 sky130_fd_sc_hd__and2_1 _15524_ (.A(_06983_),
    .B(_07002_),
    .X(_07003_));
 sky130_fd_sc_hd__nor2_1 _15525_ (.A(_06983_),
    .B(_07002_),
    .Y(_07004_));
 sky130_fd_sc_hd__nor2_1 _15526_ (.A(_07003_),
    .B(_07004_),
    .Y(_07005_));
 sky130_fd_sc_hd__a21o_1 _15527_ (.A1(_06840_),
    .A2(_06844_),
    .B1(_06866_),
    .X(_07006_));
 sky130_fd_sc_hd__nand2_1 _15528_ (.A(_07005_),
    .B(_07006_),
    .Y(_07007_));
 sky130_fd_sc_hd__xnor2_1 _15529_ (.A(_07005_),
    .B(_07006_),
    .Y(_07008_));
 sky130_fd_sc_hd__a22o_1 _15530_ (.A1(net492),
    .A2(net358),
    .B1(net353),
    .B2(net496),
    .X(_07009_));
 sky130_fd_sc_hd__nand4_2 _15531_ (.A(net497),
    .B(net492),
    .C(net358),
    .D(net353),
    .Y(_07010_));
 sky130_fd_sc_hd__a22o_1 _15532_ (.A1(net501),
    .A2(net350),
    .B1(_07009_),
    .B2(_07010_),
    .X(_07011_));
 sky130_fd_sc_hd__nand4_1 _15533_ (.A(net501),
    .B(net350),
    .C(_07009_),
    .D(_07010_),
    .Y(_07012_));
 sky130_fd_sc_hd__nand2_1 _15534_ (.A(_07011_),
    .B(_07012_),
    .Y(_07013_));
 sky130_fd_sc_hd__a22o_1 _15535_ (.A1(net369),
    .A2(net485),
    .B1(net479),
    .B2(net634),
    .X(_07014_));
 sky130_fd_sc_hd__and4_1 _15536_ (.A(net634),
    .B(net369),
    .C(net485),
    .D(net480),
    .X(_07015_));
 sky130_fd_sc_hd__inv_2 _15537_ (.A(_07015_),
    .Y(_07016_));
 sky130_fd_sc_hd__a22oi_1 _15538_ (.A1(net362),
    .A2(net489),
    .B1(_07014_),
    .B2(_07016_),
    .Y(_07017_));
 sky130_fd_sc_hd__and4_1 _15539_ (.A(net362),
    .B(net489),
    .C(_07014_),
    .D(_07016_),
    .X(_07018_));
 sky130_fd_sc_hd__or2_1 _15540_ (.A(_07017_),
    .B(_07018_),
    .X(_07019_));
 sky130_fd_sc_hd__or2_1 _15541_ (.A(_06875_),
    .B(_06878_),
    .X(_07020_));
 sky130_fd_sc_hd__nand2b_1 _15542_ (.A_N(_07019_),
    .B(_07020_),
    .Y(_07021_));
 sky130_fd_sc_hd__xor2_1 _15543_ (.A(_07019_),
    .B(_07020_),
    .X(_07022_));
 sky130_fd_sc_hd__or2_1 _15544_ (.A(_07013_),
    .B(_07022_),
    .X(_07023_));
 sky130_fd_sc_hd__nand2_1 _15545_ (.A(_07013_),
    .B(_07022_),
    .Y(_07024_));
 sky130_fd_sc_hd__and2_1 _15546_ (.A(_07023_),
    .B(_07024_),
    .X(_07025_));
 sky130_fd_sc_hd__or2_1 _15547_ (.A(_06890_),
    .B(_06892_),
    .X(_07026_));
 sky130_fd_sc_hd__nand2_2 _15548_ (.A(_06848_),
    .B(_06850_),
    .Y(_07027_));
 sky130_fd_sc_hd__a22o_1 _15549_ (.A1(net378),
    .A2(net471),
    .B1(net469),
    .B2(net384),
    .X(_07028_));
 sky130_fd_sc_hd__inv_2 _15550_ (.A(_07028_),
    .Y(_07029_));
 sky130_fd_sc_hd__and4_1 _15551_ (.A(net384),
    .B(net378),
    .C(net472),
    .D(net468),
    .X(_07030_));
 sky130_fd_sc_hd__o2bb2a_1 _15552_ (.A1_N(net372),
    .A2_N(net476),
    .B1(_07029_),
    .B2(_07030_),
    .X(_07031_));
 sky130_fd_sc_hd__and4b_1 _15553_ (.A_N(_07030_),
    .B(net476),
    .C(net372),
    .D(_07028_),
    .X(_07032_));
 sky130_fd_sc_hd__or2_1 _15554_ (.A(_07031_),
    .B(_07032_),
    .X(_07033_));
 sky130_fd_sc_hd__nand2b_1 _15555_ (.A_N(_07033_),
    .B(_07027_),
    .Y(_07034_));
 sky130_fd_sc_hd__xnor2_1 _15556_ (.A(_07027_),
    .B(_07033_),
    .Y(_07035_));
 sky130_fd_sc_hd__nand2_1 _15557_ (.A(_07026_),
    .B(_07035_),
    .Y(_07036_));
 sky130_fd_sc_hd__xnor2_1 _15558_ (.A(_07026_),
    .B(_07035_),
    .Y(_07037_));
 sky130_fd_sc_hd__a21o_1 _15559_ (.A1(_06894_),
    .A2(_06896_),
    .B1(_07037_),
    .X(_07038_));
 sky130_fd_sc_hd__nand3_2 _15560_ (.A(_06894_),
    .B(_06896_),
    .C(_07037_),
    .Y(_07039_));
 sky130_fd_sc_hd__and3_1 _15561_ (.A(_07025_),
    .B(_07038_),
    .C(_07039_),
    .X(_07040_));
 sky130_fd_sc_hd__a21oi_2 _15562_ (.A1(_07038_),
    .A2(_07039_),
    .B1(_07025_),
    .Y(_07041_));
 sky130_fd_sc_hd__a211oi_4 _15563_ (.A1(_06861_),
    .A2(_06863_),
    .B1(_07040_),
    .C1(_07041_),
    .Y(_07042_));
 sky130_fd_sc_hd__o211a_1 _15564_ (.A1(_07040_),
    .A2(_07041_),
    .B1(_06861_),
    .C1(_06863_),
    .X(_07043_));
 sky130_fd_sc_hd__a211oi_4 _15565_ (.A1(_06898_),
    .A2(_06900_),
    .B1(_07042_),
    .C1(_07043_),
    .Y(_07044_));
 sky130_fd_sc_hd__o211a_1 _15566_ (.A1(_07042_),
    .A2(_07043_),
    .B1(_06898_),
    .C1(_06900_),
    .X(_07045_));
 sky130_fd_sc_hd__or3_4 _15567_ (.A(_07008_),
    .B(_07044_),
    .C(_07045_),
    .X(_07046_));
 sky130_fd_sc_hd__o21ai_1 _15568_ (.A1(_07044_),
    .A2(_07045_),
    .B1(_07008_),
    .Y(_07047_));
 sky130_fd_sc_hd__o211a_2 _15569_ (.A1(_06868_),
    .A2(_06906_),
    .B1(_07046_),
    .C1(_07047_),
    .X(_07048_));
 sky130_fd_sc_hd__a211oi_2 _15570_ (.A1(_07046_),
    .A2(_07047_),
    .B1(_06868_),
    .C1(_06906_),
    .Y(_07049_));
 sky130_fd_sc_hd__a22o_1 _15571_ (.A1(net519),
    .A2(net335),
    .B1(net331),
    .B2(net522),
    .X(_07050_));
 sky130_fd_sc_hd__and4_1 _15572_ (.A(\mul0.a[14] ),
    .B(net522),
    .C(net335),
    .D(net332),
    .X(_07051_));
 sky130_fd_sc_hd__inv_2 _15573_ (.A(_07051_),
    .Y(_07052_));
 sky130_fd_sc_hd__a22oi_1 _15574_ (.A1(net528),
    .A2(net329),
    .B1(_07050_),
    .B2(_07052_),
    .Y(_07053_));
 sky130_fd_sc_hd__and4_1 _15575_ (.A(net528),
    .B(\mul0.b[29] ),
    .C(_07050_),
    .D(_07052_),
    .X(_07054_));
 sky130_fd_sc_hd__or2_2 _15576_ (.A(_07053_),
    .B(_07054_),
    .X(_07055_));
 sky130_fd_sc_hd__nor2_2 _15577_ (.A(_06912_),
    .B(_06915_),
    .Y(_07056_));
 sky130_fd_sc_hd__xnor2_4 _15578_ (.A(_07055_),
    .B(_07056_),
    .Y(_07057_));
 sky130_fd_sc_hd__and4b_2 _15579_ (.A_N(net539),
    .B(\mul0.b[30] ),
    .C(net326),
    .D(net534),
    .X(_07058_));
 sky130_fd_sc_hd__o2bb2a_1 _15580_ (.A1_N(net533),
    .A2_N(\mul0.b[30] ),
    .B1(net57),
    .B2(net539),
    .X(_07059_));
 sky130_fd_sc_hd__nor2_1 _15581_ (.A(_07058_),
    .B(_07059_),
    .Y(_07060_));
 sky130_fd_sc_hd__xnor2_2 _15582_ (.A(_07057_),
    .B(_07060_),
    .Y(_07061_));
 sky130_fd_sc_hd__o32ai_4 _15583_ (.A1(_06918_),
    .A2(_06919_),
    .A3(_06921_),
    .B1(_06917_),
    .B2(_06916_),
    .Y(_07062_));
 sky130_fd_sc_hd__nand2_1 _15584_ (.A(_07061_),
    .B(_07062_),
    .Y(_07063_));
 sky130_fd_sc_hd__xnor2_2 _15585_ (.A(_07061_),
    .B(_07062_),
    .Y(_07064_));
 sky130_fd_sc_hd__xnor2_2 _15586_ (.A(_06920_),
    .B(_07064_),
    .Y(_07065_));
 sky130_fd_sc_hd__or2_1 _15587_ (.A(_06934_),
    .B(_06936_),
    .X(_07066_));
 sky130_fd_sc_hd__nand2_1 _15588_ (.A(_06870_),
    .B(_06872_),
    .Y(_07067_));
 sky130_fd_sc_hd__a22o_1 _15589_ (.A1(net506),
    .A2(net346),
    .B1(net342),
    .B2(net509),
    .X(_07068_));
 sky130_fd_sc_hd__inv_2 _15590_ (.A(_07068_),
    .Y(_07069_));
 sky130_fd_sc_hd__and4_1 _15591_ (.A(net506),
    .B(net509),
    .C(net346),
    .D(net342),
    .X(_07070_));
 sky130_fd_sc_hd__o2bb2a_1 _15592_ (.A1_N(net514),
    .A2_N(net338),
    .B1(_07069_),
    .B2(_07070_),
    .X(_07071_));
 sky130_fd_sc_hd__and4b_1 _15593_ (.A_N(_07070_),
    .B(net338),
    .C(net513),
    .D(_07068_),
    .X(_07072_));
 sky130_fd_sc_hd__or2_1 _15594_ (.A(_07071_),
    .B(_07072_),
    .X(_07073_));
 sky130_fd_sc_hd__nand2b_1 _15595_ (.A_N(_07073_),
    .B(_07067_),
    .Y(_07074_));
 sky130_fd_sc_hd__xnor2_2 _15596_ (.A(_07067_),
    .B(_07073_),
    .Y(_07075_));
 sky130_fd_sc_hd__nand2_1 _15597_ (.A(_07066_),
    .B(_07075_),
    .Y(_07076_));
 sky130_fd_sc_hd__xnor2_2 _15598_ (.A(_07066_),
    .B(_07075_),
    .Y(_07077_));
 sky130_fd_sc_hd__a21oi_4 _15599_ (.A1(_06881_),
    .A2(_06883_),
    .B1(_07077_),
    .Y(_07078_));
 sky130_fd_sc_hd__and3_1 _15600_ (.A(_06881_),
    .B(_06883_),
    .C(_07077_),
    .X(_07079_));
 sky130_fd_sc_hd__a211oi_4 _15601_ (.A1(_06938_),
    .A2(_06940_),
    .B1(_07078_),
    .C1(_07079_),
    .Y(_07080_));
 sky130_fd_sc_hd__o211a_1 _15602_ (.A1(_07078_),
    .A2(_07079_),
    .B1(_06938_),
    .C1(_06940_),
    .X(_07081_));
 sky130_fd_sc_hd__a211oi_2 _15603_ (.A1(_06943_),
    .A2(_06945_),
    .B1(_07080_),
    .C1(_07081_),
    .Y(_07082_));
 sky130_fd_sc_hd__o211a_1 _15604_ (.A1(_07080_),
    .A2(_07081_),
    .B1(_06943_),
    .C1(_06945_),
    .X(_07083_));
 sky130_fd_sc_hd__or3_2 _15605_ (.A(_07065_),
    .B(_07082_),
    .C(_07083_),
    .X(_07084_));
 sky130_fd_sc_hd__o21ai_2 _15606_ (.A1(_07082_),
    .A2(_07083_),
    .B1(_07065_),
    .Y(_07085_));
 sky130_fd_sc_hd__o211a_1 _15607_ (.A1(_06902_),
    .A2(_06904_),
    .B1(_07084_),
    .C1(_07085_),
    .X(_07086_));
 sky130_fd_sc_hd__o211ai_2 _15608_ (.A1(_06902_),
    .A2(_06904_),
    .B1(_07084_),
    .C1(_07085_),
    .Y(_07087_));
 sky130_fd_sc_hd__a211o_1 _15609_ (.A1(_07084_),
    .A2(_07085_),
    .B1(_06902_),
    .C1(_06904_),
    .X(_07088_));
 sky130_fd_sc_hd__o211a_2 _15610_ (.A1(_06947_),
    .A2(_06949_),
    .B1(_07087_),
    .C1(_07088_),
    .X(_07089_));
 sky130_fd_sc_hd__a211oi_2 _15611_ (.A1(_07087_),
    .A2(_07088_),
    .B1(_06947_),
    .C1(_06949_),
    .Y(_07090_));
 sky130_fd_sc_hd__nor4_4 _15612_ (.A(_07048_),
    .B(_07049_),
    .C(_07089_),
    .D(_07090_),
    .Y(_07091_));
 sky130_fd_sc_hd__o22a_1 _15613_ (.A1(_07048_),
    .A2(_07049_),
    .B1(_07089_),
    .B2(_07090_),
    .X(_07092_));
 sky130_fd_sc_hd__a211oi_4 _15614_ (.A1(_06908_),
    .A2(_06955_),
    .B1(_07091_),
    .C1(_07092_),
    .Y(_07093_));
 sky130_fd_sc_hd__o211a_1 _15615_ (.A1(_07091_),
    .A2(_07092_),
    .B1(_06908_),
    .C1(_06955_),
    .X(_07094_));
 sky130_fd_sc_hd__a211oi_4 _15616_ (.A1(_06951_),
    .A2(_06953_),
    .B1(_07093_),
    .C1(_07094_),
    .Y(_07095_));
 sky130_fd_sc_hd__o211a_1 _15617_ (.A1(_07093_),
    .A2(_07094_),
    .B1(_06951_),
    .C1(_06953_),
    .X(_07096_));
 sky130_fd_sc_hd__a211oi_4 _15618_ (.A1(_06957_),
    .A2(_06959_),
    .B1(_07095_),
    .C1(_07096_),
    .Y(_07097_));
 sky130_fd_sc_hd__o211a_1 _15619_ (.A1(_07095_),
    .A2(_07096_),
    .B1(_06957_),
    .C1(_06959_),
    .X(_07098_));
 sky130_fd_sc_hd__a211oi_2 _15620_ (.A1(_06925_),
    .A2(_06928_),
    .B1(_07097_),
    .C1(_07098_),
    .Y(_07099_));
 sky130_fd_sc_hd__o211a_1 _15621_ (.A1(_07097_),
    .A2(_07098_),
    .B1(_06925_),
    .C1(_06928_),
    .X(_07100_));
 sky130_fd_sc_hd__a211oi_2 _15622_ (.A1(_06963_),
    .A2(_06966_),
    .B1(_07099_),
    .C1(_07100_),
    .Y(_07101_));
 sky130_fd_sc_hd__o211ai_2 _15623_ (.A1(_07099_),
    .A2(_07100_),
    .B1(_06963_),
    .C1(_06966_),
    .Y(_07102_));
 sky130_fd_sc_hd__nand2b_1 _15624_ (.A_N(_07101_),
    .B(_07102_),
    .Y(_07103_));
 sky130_fd_sc_hd__or2_2 _15625_ (.A(_06969_),
    .B(_06975_),
    .X(_07104_));
 sky130_fd_sc_hd__xnor2_2 _15626_ (.A(_07103_),
    .B(_07104_),
    .Y(_07105_));
 sky130_fd_sc_hd__a22o_1 _15627_ (.A1(net599),
    .A2(net831),
    .B1(_02700_),
    .B2(net5),
    .X(_07106_));
 sky130_fd_sc_hd__a21o_1 _15628_ (.A1(_03058_),
    .A2(_07105_),
    .B1(_07106_),
    .X(_07107_));
 sky130_fd_sc_hd__mux2_1 _15629_ (.A0(net909),
    .A1(_07107_),
    .S(net4),
    .X(_00291_));
 sky130_fd_sc_hd__a32o_2 _15630_ (.A1(_06988_),
    .A2(_06989_),
    .A3(_06997_),
    .B1(_06996_),
    .B2(_06991_),
    .X(_07108_));
 sky130_fd_sc_hd__a22o_1 _15631_ (.A1(net393),
    .A2(net458),
    .B1(net455),
    .B2(net398),
    .X(_07109_));
 sky130_fd_sc_hd__and4_1 _15632_ (.A(net398),
    .B(net393),
    .C(net458),
    .D(net456),
    .X(_07110_));
 sky130_fd_sc_hd__inv_2 _15633_ (.A(_07110_),
    .Y(_07111_));
 sky130_fd_sc_hd__a22oi_1 _15634_ (.A1(net388),
    .A2(net462),
    .B1(_07109_),
    .B2(_07111_),
    .Y(_07112_));
 sky130_fd_sc_hd__and4_1 _15635_ (.A(net388),
    .B(net462),
    .C(_07109_),
    .D(_07111_),
    .X(_07113_));
 sky130_fd_sc_hd__or2_2 _15636_ (.A(_07112_),
    .B(_07113_),
    .X(_07114_));
 sky130_fd_sc_hd__a21oi_2 _15637_ (.A1(net403),
    .A2(net454),
    .B1(_06994_),
    .Y(_07115_));
 sky130_fd_sc_hd__a21o_1 _15638_ (.A1(_06992_),
    .A2(_06994_),
    .B1(_06993_),
    .X(_07116_));
 sky130_fd_sc_hd__a21oi_2 _15639_ (.A1(net403),
    .A2(_07116_),
    .B1(_07115_),
    .Y(_07117_));
 sky130_fd_sc_hd__or3b_1 _15640_ (.A(_07112_),
    .B(_07113_),
    .C_N(_07117_),
    .X(_07118_));
 sky130_fd_sc_hd__xnor2_4 _15641_ (.A(_07114_),
    .B(_07117_),
    .Y(_07119_));
 sky130_fd_sc_hd__nand2_1 _15642_ (.A(_06985_),
    .B(_07119_),
    .Y(_07120_));
 sky130_fd_sc_hd__xor2_1 _15643_ (.A(_06985_),
    .B(_07119_),
    .X(_07121_));
 sky130_fd_sc_hd__nand2_1 _15644_ (.A(_07108_),
    .B(_07121_),
    .Y(_07122_));
 sky130_fd_sc_hd__xnor2_1 _15645_ (.A(_07108_),
    .B(_07121_),
    .Y(_07123_));
 sky130_fd_sc_hd__nor2_1 _15646_ (.A(_06983_),
    .B(_07123_),
    .Y(_07124_));
 sky130_fd_sc_hd__xnor2_1 _15647_ (.A(_06982_),
    .B(_07123_),
    .Y(_07125_));
 sky130_fd_sc_hd__nor3_1 _15648_ (.A(_06980_),
    .B(_07004_),
    .C(_07125_),
    .Y(_07126_));
 sky130_fd_sc_hd__o21a_1 _15649_ (.A1(_06980_),
    .A2(_07004_),
    .B1(_07125_),
    .X(_07127_));
 sky130_fd_sc_hd__or2_1 _15650_ (.A(_07126_),
    .B(_07127_),
    .X(_07128_));
 sky130_fd_sc_hd__a21boi_1 _15651_ (.A1(_07025_),
    .A2(_07039_),
    .B1_N(_07038_),
    .Y(_07129_));
 sky130_fd_sc_hd__a22o_1 _15652_ (.A1(net489),
    .A2(net358),
    .B1(net353),
    .B2(net492),
    .X(_07130_));
 sky130_fd_sc_hd__nand4_2 _15653_ (.A(net492),
    .B(net489),
    .C(net357),
    .D(net353),
    .Y(_07131_));
 sky130_fd_sc_hd__a22o_1 _15654_ (.A1(net497),
    .A2(net350),
    .B1(_07130_),
    .B2(_07131_),
    .X(_07132_));
 sky130_fd_sc_hd__nand4_1 _15655_ (.A(net497),
    .B(net350),
    .C(_07130_),
    .D(_07131_),
    .Y(_07133_));
 sky130_fd_sc_hd__nand2_1 _15656_ (.A(_07132_),
    .B(_07133_),
    .Y(_07134_));
 sky130_fd_sc_hd__a22o_1 _15657_ (.A1(net369),
    .A2(net480),
    .B1(net476),
    .B2(net634),
    .X(_07135_));
 sky130_fd_sc_hd__and4_1 _15658_ (.A(net634),
    .B(net369),
    .C(net480),
    .D(net476),
    .X(_07136_));
 sky130_fd_sc_hd__inv_2 _15659_ (.A(_07136_),
    .Y(_07137_));
 sky130_fd_sc_hd__a22oi_1 _15660_ (.A1(net362),
    .A2(net484),
    .B1(_07135_),
    .B2(_07137_),
    .Y(_07138_));
 sky130_fd_sc_hd__and4_1 _15661_ (.A(net362),
    .B(net484),
    .C(_07135_),
    .D(_07137_),
    .X(_07139_));
 sky130_fd_sc_hd__or2_1 _15662_ (.A(_07138_),
    .B(_07139_),
    .X(_07140_));
 sky130_fd_sc_hd__or2_1 _15663_ (.A(_07015_),
    .B(_07018_),
    .X(_07141_));
 sky130_fd_sc_hd__nand2b_1 _15664_ (.A_N(_07140_),
    .B(_07141_),
    .Y(_07142_));
 sky130_fd_sc_hd__xor2_1 _15665_ (.A(_07140_),
    .B(_07141_),
    .X(_07143_));
 sky130_fd_sc_hd__or2_1 _15666_ (.A(_07134_),
    .B(_07143_),
    .X(_07144_));
 sky130_fd_sc_hd__nand2_1 _15667_ (.A(_07134_),
    .B(_07143_),
    .Y(_07145_));
 sky130_fd_sc_hd__and2_1 _15668_ (.A(_07144_),
    .B(_07145_),
    .X(_07146_));
 sky130_fd_sc_hd__or2_1 _15669_ (.A(_07030_),
    .B(_07032_),
    .X(_07147_));
 sky130_fd_sc_hd__nand2_2 _15670_ (.A(_06987_),
    .B(_06989_),
    .Y(_07148_));
 sky130_fd_sc_hd__a22o_1 _15671_ (.A1(net378),
    .A2(net469),
    .B1(net465),
    .B2(net384),
    .X(_07149_));
 sky130_fd_sc_hd__inv_2 _15672_ (.A(_07149_),
    .Y(_07150_));
 sky130_fd_sc_hd__and4_1 _15673_ (.A(net384),
    .B(net378),
    .C(net468),
    .D(net465),
    .X(_07151_));
 sky130_fd_sc_hd__o2bb2a_1 _15674_ (.A1_N(net373),
    .A2_N(net472),
    .B1(_07150_),
    .B2(_07151_),
    .X(_07152_));
 sky130_fd_sc_hd__and4b_1 _15675_ (.A_N(_07151_),
    .B(net472),
    .C(net372),
    .D(_07149_),
    .X(_07153_));
 sky130_fd_sc_hd__or2_1 _15676_ (.A(_07152_),
    .B(_07153_),
    .X(_07154_));
 sky130_fd_sc_hd__nand2b_1 _15677_ (.A_N(_07154_),
    .B(_07148_),
    .Y(_07155_));
 sky130_fd_sc_hd__xnor2_1 _15678_ (.A(_07148_),
    .B(_07154_),
    .Y(_07156_));
 sky130_fd_sc_hd__nand2_1 _15679_ (.A(_07147_),
    .B(_07156_),
    .Y(_07157_));
 sky130_fd_sc_hd__xnor2_1 _15680_ (.A(_07147_),
    .B(_07156_),
    .Y(_07158_));
 sky130_fd_sc_hd__a21o_2 _15681_ (.A1(_07034_),
    .A2(_07036_),
    .B1(_07158_),
    .X(_07159_));
 sky130_fd_sc_hd__nand3_2 _15682_ (.A(_07034_),
    .B(_07036_),
    .C(_07158_),
    .Y(_07160_));
 sky130_fd_sc_hd__nand3_4 _15683_ (.A(_07146_),
    .B(_07159_),
    .C(_07160_),
    .Y(_07161_));
 sky130_fd_sc_hd__a21o_1 _15684_ (.A1(_07159_),
    .A2(_07160_),
    .B1(_07146_),
    .X(_07162_));
 sky130_fd_sc_hd__o211a_2 _15685_ (.A1(_06999_),
    .A2(_07001_),
    .B1(_07161_),
    .C1(_07162_),
    .X(_07163_));
 sky130_fd_sc_hd__a211oi_2 _15686_ (.A1(_07161_),
    .A2(_07162_),
    .B1(_06999_),
    .C1(_07001_),
    .Y(_07164_));
 sky130_fd_sc_hd__nor3_2 _15687_ (.A(_07129_),
    .B(_07163_),
    .C(_07164_),
    .Y(_07165_));
 sky130_fd_sc_hd__o21a_1 _15688_ (.A1(_07163_),
    .A2(_07164_),
    .B1(_07129_),
    .X(_07166_));
 sky130_fd_sc_hd__nor3_4 _15689_ (.A(_07128_),
    .B(_07165_),
    .C(_07166_),
    .Y(_07167_));
 sky130_fd_sc_hd__o21a_1 _15690_ (.A1(_07165_),
    .A2(_07166_),
    .B1(_07128_),
    .X(_07168_));
 sky130_fd_sc_hd__a211oi_4 _15691_ (.A1(_07007_),
    .A2(_07046_),
    .B1(_07167_),
    .C1(_07168_),
    .Y(_07169_));
 sky130_fd_sc_hd__o211a_1 _15692_ (.A1(_07167_),
    .A2(_07168_),
    .B1(_07007_),
    .C1(_07046_),
    .X(_07170_));
 sky130_fd_sc_hd__nand2b_1 _15693_ (.A_N(_07082_),
    .B(_07084_),
    .Y(_07171_));
 sky130_fd_sc_hd__a22o_1 _15694_ (.A1(net514),
    .A2(net335),
    .B1(net332),
    .B2(net518),
    .X(_07172_));
 sky130_fd_sc_hd__and4_1 _15695_ (.A(net514),
    .B(net518),
    .C(net335),
    .D(net332),
    .X(_07173_));
 sky130_fd_sc_hd__inv_2 _15696_ (.A(_07173_),
    .Y(_07174_));
 sky130_fd_sc_hd__a22oi_1 _15697_ (.A1(net522),
    .A2(net329),
    .B1(_07172_),
    .B2(_07174_),
    .Y(_07175_));
 sky130_fd_sc_hd__and4_1 _15698_ (.A(net522),
    .B(net329),
    .C(_07172_),
    .D(_07174_),
    .X(_07176_));
 sky130_fd_sc_hd__or2_2 _15699_ (.A(_07175_),
    .B(_07176_),
    .X(_07177_));
 sky130_fd_sc_hd__nor2_2 _15700_ (.A(_07051_),
    .B(_07054_),
    .Y(_07178_));
 sky130_fd_sc_hd__xnor2_2 _15701_ (.A(_07177_),
    .B(_07178_),
    .Y(_07179_));
 sky130_fd_sc_hd__and4b_2 _15702_ (.A_N(net533),
    .B(net327),
    .C(net326),
    .D(net528),
    .X(_07180_));
 sky130_fd_sc_hd__inv_2 _15703_ (.A(_07180_),
    .Y(_07181_));
 sky130_fd_sc_hd__o2bb2a_1 _15704_ (.A1_N(net528),
    .A2_N(net327),
    .B1(net57),
    .B2(net533),
    .X(_07182_));
 sky130_fd_sc_hd__nor2_1 _15705_ (.A(_07180_),
    .B(_07182_),
    .Y(_07183_));
 sky130_fd_sc_hd__xnor2_2 _15706_ (.A(_07179_),
    .B(_07183_),
    .Y(_07184_));
 sky130_fd_sc_hd__o32ai_4 _15707_ (.A1(_07057_),
    .A2(_07058_),
    .A3(_07059_),
    .B1(_07056_),
    .B2(_07055_),
    .Y(_07185_));
 sky130_fd_sc_hd__nand2_1 _15708_ (.A(_07184_),
    .B(_07185_),
    .Y(_07186_));
 sky130_fd_sc_hd__xnor2_2 _15709_ (.A(_07184_),
    .B(_07185_),
    .Y(_07187_));
 sky130_fd_sc_hd__inv_2 _15710_ (.A(_07187_),
    .Y(_07188_));
 sky130_fd_sc_hd__nand2_1 _15711_ (.A(_07058_),
    .B(_07188_),
    .Y(_07189_));
 sky130_fd_sc_hd__xor2_2 _15712_ (.A(_07058_),
    .B(_07187_),
    .X(_07190_));
 sky130_fd_sc_hd__or2_1 _15713_ (.A(_07070_),
    .B(_07072_),
    .X(_07191_));
 sky130_fd_sc_hd__nand2_1 _15714_ (.A(_07010_),
    .B(_07012_),
    .Y(_07192_));
 sky130_fd_sc_hd__a22o_1 _15715_ (.A1(net501),
    .A2(net346),
    .B1(net342),
    .B2(net505),
    .X(_07193_));
 sky130_fd_sc_hd__inv_2 _15716_ (.A(_07193_),
    .Y(_07194_));
 sky130_fd_sc_hd__and4_1 _15717_ (.A(net505),
    .B(net501),
    .C(net346),
    .D(net342),
    .X(_07195_));
 sky130_fd_sc_hd__o2bb2a_1 _15718_ (.A1_N(net509),
    .A2_N(net338),
    .B1(_07194_),
    .B2(_07195_),
    .X(_07196_));
 sky130_fd_sc_hd__and4b_1 _15719_ (.A_N(_07195_),
    .B(net338),
    .C(net509),
    .D(_07193_),
    .X(_07197_));
 sky130_fd_sc_hd__or2_1 _15720_ (.A(_07196_),
    .B(_07197_),
    .X(_07198_));
 sky130_fd_sc_hd__nand2b_1 _15721_ (.A_N(_07198_),
    .B(_07192_),
    .Y(_07199_));
 sky130_fd_sc_hd__xnor2_1 _15722_ (.A(_07192_),
    .B(_07198_),
    .Y(_07200_));
 sky130_fd_sc_hd__nand2_1 _15723_ (.A(_07191_),
    .B(_07200_),
    .Y(_07201_));
 sky130_fd_sc_hd__xnor2_1 _15724_ (.A(_07191_),
    .B(_07200_),
    .Y(_07202_));
 sky130_fd_sc_hd__a21oi_1 _15725_ (.A1(_07021_),
    .A2(_07023_),
    .B1(_07202_),
    .Y(_07203_));
 sky130_fd_sc_hd__a21o_1 _15726_ (.A1(_07021_),
    .A2(_07023_),
    .B1(_07202_),
    .X(_07204_));
 sky130_fd_sc_hd__and3_1 _15727_ (.A(_07021_),
    .B(_07023_),
    .C(_07202_),
    .X(_07205_));
 sky130_fd_sc_hd__a211o_1 _15728_ (.A1(_07074_),
    .A2(_07076_),
    .B1(_07203_),
    .C1(_07205_),
    .X(_07206_));
 sky130_fd_sc_hd__o211ai_2 _15729_ (.A1(_07203_),
    .A2(_07205_),
    .B1(_07074_),
    .C1(_07076_),
    .Y(_07207_));
 sky130_fd_sc_hd__o211a_1 _15730_ (.A1(_07078_),
    .A2(_07080_),
    .B1(_07206_),
    .C1(_07207_),
    .X(_07208_));
 sky130_fd_sc_hd__a211oi_2 _15731_ (.A1(_07206_),
    .A2(_07207_),
    .B1(_07078_),
    .C1(_07080_),
    .Y(_07209_));
 sky130_fd_sc_hd__nor3_1 _15732_ (.A(_07190_),
    .B(_07208_),
    .C(_07209_),
    .Y(_07210_));
 sky130_fd_sc_hd__or3_2 _15733_ (.A(_07190_),
    .B(_07208_),
    .C(_07209_),
    .X(_07211_));
 sky130_fd_sc_hd__o21ai_2 _15734_ (.A1(_07208_),
    .A2(_07209_),
    .B1(_07190_),
    .Y(_07212_));
 sky130_fd_sc_hd__o211ai_4 _15735_ (.A1(_07042_),
    .A2(_07044_),
    .B1(_07211_),
    .C1(_07212_),
    .Y(_07213_));
 sky130_fd_sc_hd__a211o_1 _15736_ (.A1(_07211_),
    .A2(_07212_),
    .B1(_07042_),
    .C1(_07044_),
    .X(_07214_));
 sky130_fd_sc_hd__and3_2 _15737_ (.A(_07171_),
    .B(_07213_),
    .C(_07214_),
    .X(_07215_));
 sky130_fd_sc_hd__inv_2 _15738_ (.A(_07215_),
    .Y(_07216_));
 sky130_fd_sc_hd__a21oi_2 _15739_ (.A1(_07213_),
    .A2(_07214_),
    .B1(_07171_),
    .Y(_07217_));
 sky130_fd_sc_hd__nor4_1 _15740_ (.A(_07169_),
    .B(_07170_),
    .C(_07215_),
    .D(_07217_),
    .Y(_07218_));
 sky130_fd_sc_hd__or4_2 _15741_ (.A(_07169_),
    .B(_07170_),
    .C(_07215_),
    .D(_07217_),
    .X(_07219_));
 sky130_fd_sc_hd__o22ai_4 _15742_ (.A1(_07169_),
    .A2(_07170_),
    .B1(_07215_),
    .B2(_07217_),
    .Y(_07220_));
 sky130_fd_sc_hd__o211ai_4 _15743_ (.A1(_07048_),
    .A2(_07091_),
    .B1(_07219_),
    .C1(_07220_),
    .Y(_07221_));
 sky130_fd_sc_hd__a211o_1 _15744_ (.A1(_07219_),
    .A2(_07220_),
    .B1(_07048_),
    .C1(_07091_),
    .X(_07222_));
 sky130_fd_sc_hd__o211ai_4 _15745_ (.A1(_07086_),
    .A2(_07089_),
    .B1(_07221_),
    .C1(_07222_),
    .Y(_07223_));
 sky130_fd_sc_hd__a211o_1 _15746_ (.A1(_07221_),
    .A2(_07222_),
    .B1(_07086_),
    .C1(_07089_),
    .X(_07224_));
 sky130_fd_sc_hd__o211ai_4 _15747_ (.A1(_07093_),
    .A2(_07095_),
    .B1(_07223_),
    .C1(_07224_),
    .Y(_07225_));
 sky130_fd_sc_hd__a211o_1 _15748_ (.A1(_07223_),
    .A2(_07224_),
    .B1(_07093_),
    .C1(_07095_),
    .X(_07226_));
 sky130_fd_sc_hd__nand2_1 _15749_ (.A(_07225_),
    .B(_07226_),
    .Y(_07227_));
 sky130_fd_sc_hd__o21a_1 _15750_ (.A1(_06920_),
    .A2(_07064_),
    .B1(_07063_),
    .X(_07228_));
 sky130_fd_sc_hd__or2_1 _15751_ (.A(_07227_),
    .B(_07228_),
    .X(_07229_));
 sky130_fd_sc_hd__xnor2_1 _15752_ (.A(_07227_),
    .B(_07228_),
    .Y(_07230_));
 sky130_fd_sc_hd__nor2_1 _15753_ (.A(_07097_),
    .B(_07099_),
    .Y(_07231_));
 sky130_fd_sc_hd__or2_1 _15754_ (.A(_07230_),
    .B(_07231_),
    .X(_07232_));
 sky130_fd_sc_hd__nand2_1 _15755_ (.A(_07230_),
    .B(_07231_),
    .Y(_07233_));
 sky130_fd_sc_hd__nand2_1 _15756_ (.A(_07232_),
    .B(_07233_),
    .Y(_07234_));
 sky130_fd_sc_hd__o21ai_2 _15757_ (.A1(_07101_),
    .A2(_07104_),
    .B1(_07102_),
    .Y(_07235_));
 sky130_fd_sc_hd__xnor2_2 _15758_ (.A(_07234_),
    .B(_07235_),
    .Y(_07236_));
 sky130_fd_sc_hd__nor2_1 _15759_ (.A(_03057_),
    .B(_07236_),
    .Y(_07237_));
 sky130_fd_sc_hd__a221o_1 _15760_ (.A1(net600),
    .A2(net758),
    .B1(_02703_),
    .B2(net5),
    .C1(_07237_),
    .X(_07238_));
 sky130_fd_sc_hd__mux2_1 _15761_ (.A0(net724),
    .A1(_07238_),
    .S(net2),
    .X(_00292_));
 sky130_fd_sc_hd__and2_2 _15762_ (.A(net403),
    .B(_06993_),
    .X(_07239_));
 sky130_fd_sc_hd__nand2_1 _15763_ (.A(net403),
    .B(_06993_),
    .Y(_07240_));
 sky130_fd_sc_hd__nand2_1 _15764_ (.A(_07118_),
    .B(_07240_),
    .Y(_07241_));
 sky130_fd_sc_hd__a22oi_1 _15765_ (.A1(net394),
    .A2(net455),
    .B1(net453),
    .B2(net398),
    .Y(_07242_));
 sky130_fd_sc_hd__and4_1 _15766_ (.A(net398),
    .B(net394),
    .C(net455),
    .D(net453),
    .X(_07243_));
 sky130_fd_sc_hd__nor2_1 _15767_ (.A(_07242_),
    .B(_07243_),
    .Y(_07244_));
 sky130_fd_sc_hd__nand2_1 _15768_ (.A(net389),
    .B(net458),
    .Y(_07245_));
 sky130_fd_sc_hd__xor2_1 _15769_ (.A(_07244_),
    .B(_07245_),
    .X(_07246_));
 sky130_fd_sc_hd__or2_2 _15770_ (.A(_07115_),
    .B(_07239_),
    .X(_07247_));
 sky130_fd_sc_hd__nor2_1 _15771_ (.A(_07246_),
    .B(_07247_),
    .Y(_07248_));
 sky130_fd_sc_hd__and2_1 _15772_ (.A(_07246_),
    .B(_07247_),
    .X(_07249_));
 sky130_fd_sc_hd__nor2_1 _15773_ (.A(_07248_),
    .B(_07249_),
    .Y(_07250_));
 sky130_fd_sc_hd__nand2_2 _15774_ (.A(_06985_),
    .B(_07250_),
    .Y(_07251_));
 sky130_fd_sc_hd__or2_1 _15775_ (.A(_06985_),
    .B(_07250_),
    .X(_07252_));
 sky130_fd_sc_hd__nand2_1 _15776_ (.A(_07251_),
    .B(_07252_),
    .Y(_07253_));
 sky130_fd_sc_hd__nand2b_1 _15777_ (.A_N(_07253_),
    .B(_07241_),
    .Y(_07254_));
 sky130_fd_sc_hd__xor2_1 _15778_ (.A(_07241_),
    .B(_07253_),
    .X(_07255_));
 sky130_fd_sc_hd__and2_1 _15779_ (.A(_06983_),
    .B(_07255_),
    .X(_07256_));
 sky130_fd_sc_hd__nor2_1 _15780_ (.A(_06983_),
    .B(_07255_),
    .Y(_07257_));
 sky130_fd_sc_hd__nor2_1 _15781_ (.A(_07256_),
    .B(_07257_),
    .Y(_07258_));
 sky130_fd_sc_hd__or3_1 _15782_ (.A(_06980_),
    .B(_07124_),
    .C(_07258_),
    .X(_07259_));
 sky130_fd_sc_hd__o21ai_2 _15783_ (.A1(_06980_),
    .A2(_07124_),
    .B1(_07258_),
    .Y(_07260_));
 sky130_fd_sc_hd__nand2_1 _15784_ (.A(_07259_),
    .B(_07260_),
    .Y(_07261_));
 sky130_fd_sc_hd__a22o_1 _15785_ (.A1(net357),
    .A2(net485),
    .B1(net353),
    .B2(net489),
    .X(_07262_));
 sky130_fd_sc_hd__nand4_1 _15786_ (.A(net488),
    .B(net358),
    .C(net485),
    .D(net353),
    .Y(_07263_));
 sky130_fd_sc_hd__a22o_1 _15787_ (.A1(net493),
    .A2(net349),
    .B1(_07262_),
    .B2(_07263_),
    .X(_07264_));
 sky130_fd_sc_hd__nand4_1 _15788_ (.A(net493),
    .B(net349),
    .C(_07262_),
    .D(_07263_),
    .Y(_07265_));
 sky130_fd_sc_hd__nand2_1 _15789_ (.A(_07264_),
    .B(_07265_),
    .Y(_07266_));
 sky130_fd_sc_hd__a22o_1 _15790_ (.A1(net369),
    .A2(net476),
    .B1(net472),
    .B2(net634),
    .X(_07267_));
 sky130_fd_sc_hd__and4_1 _15791_ (.A(net634),
    .B(net369),
    .C(net476),
    .D(net472),
    .X(_07268_));
 sky130_fd_sc_hd__inv_2 _15792_ (.A(_07268_),
    .Y(_07269_));
 sky130_fd_sc_hd__a22oi_1 _15793_ (.A1(net362),
    .A2(net480),
    .B1(_07267_),
    .B2(_07269_),
    .Y(_07270_));
 sky130_fd_sc_hd__and4_1 _15794_ (.A(net362),
    .B(net480),
    .C(_07267_),
    .D(_07269_),
    .X(_07271_));
 sky130_fd_sc_hd__or2_1 _15795_ (.A(_07270_),
    .B(_07271_),
    .X(_07272_));
 sky130_fd_sc_hd__or2_1 _15796_ (.A(_07136_),
    .B(_07139_),
    .X(_07273_));
 sky130_fd_sc_hd__nand2b_1 _15797_ (.A_N(_07272_),
    .B(_07273_),
    .Y(_07274_));
 sky130_fd_sc_hd__xor2_1 _15798_ (.A(_07272_),
    .B(_07273_),
    .X(_07275_));
 sky130_fd_sc_hd__or2_1 _15799_ (.A(_07266_),
    .B(_07275_),
    .X(_07276_));
 sky130_fd_sc_hd__nand2_1 _15800_ (.A(_07266_),
    .B(_07275_),
    .Y(_07277_));
 sky130_fd_sc_hd__and2_1 _15801_ (.A(_07276_),
    .B(_07277_),
    .X(_07278_));
 sky130_fd_sc_hd__or2_1 _15802_ (.A(_07151_),
    .B(_07153_),
    .X(_07279_));
 sky130_fd_sc_hd__nor2_1 _15803_ (.A(_07110_),
    .B(_07113_),
    .Y(_07280_));
 sky130_fd_sc_hd__a22o_1 _15804_ (.A1(net378),
    .A2(net465),
    .B1(net462),
    .B2(net384),
    .X(_07281_));
 sky130_fd_sc_hd__inv_2 _15805_ (.A(_07281_),
    .Y(_07282_));
 sky130_fd_sc_hd__and4_1 _15806_ (.A(net384),
    .B(net378),
    .C(net465),
    .D(net462),
    .X(_07283_));
 sky130_fd_sc_hd__o2bb2a_1 _15807_ (.A1_N(net372),
    .A2_N(net468),
    .B1(_07282_),
    .B2(_07283_),
    .X(_07284_));
 sky130_fd_sc_hd__and4b_1 _15808_ (.A_N(_07283_),
    .B(net468),
    .C(net372),
    .D(_07281_),
    .X(_07285_));
 sky130_fd_sc_hd__or2_1 _15809_ (.A(_07284_),
    .B(_07285_),
    .X(_07286_));
 sky130_fd_sc_hd__or2_1 _15810_ (.A(_07280_),
    .B(_07286_),
    .X(_07287_));
 sky130_fd_sc_hd__xor2_1 _15811_ (.A(_07280_),
    .B(_07286_),
    .X(_07288_));
 sky130_fd_sc_hd__nand2_1 _15812_ (.A(_07279_),
    .B(_07288_),
    .Y(_07289_));
 sky130_fd_sc_hd__xnor2_1 _15813_ (.A(_07279_),
    .B(_07288_),
    .Y(_07290_));
 sky130_fd_sc_hd__a21o_2 _15814_ (.A1(_07155_),
    .A2(_07157_),
    .B1(_07290_),
    .X(_07291_));
 sky130_fd_sc_hd__nand3_1 _15815_ (.A(_07155_),
    .B(_07157_),
    .C(_07290_),
    .Y(_07292_));
 sky130_fd_sc_hd__and3_2 _15816_ (.A(_07278_),
    .B(_07291_),
    .C(_07292_),
    .X(_07293_));
 sky130_fd_sc_hd__inv_2 _15817_ (.A(_07293_),
    .Y(_07294_));
 sky130_fd_sc_hd__a21oi_2 _15818_ (.A1(_07291_),
    .A2(_07292_),
    .B1(_07278_),
    .Y(_07295_));
 sky130_fd_sc_hd__a211oi_4 _15819_ (.A1(_07120_),
    .A2(_07122_),
    .B1(_07293_),
    .C1(_07295_),
    .Y(_07296_));
 sky130_fd_sc_hd__o211a_1 _15820_ (.A1(_07293_),
    .A2(_07295_),
    .B1(_07120_),
    .C1(_07122_),
    .X(_07297_));
 sky130_fd_sc_hd__a211oi_4 _15821_ (.A1(_07159_),
    .A2(_07161_),
    .B1(_07296_),
    .C1(_07297_),
    .Y(_07298_));
 sky130_fd_sc_hd__o211a_1 _15822_ (.A1(_07296_),
    .A2(_07297_),
    .B1(_07159_),
    .C1(_07161_),
    .X(_07299_));
 sky130_fd_sc_hd__or3_4 _15823_ (.A(_07261_),
    .B(_07298_),
    .C(_07299_),
    .X(_07300_));
 sky130_fd_sc_hd__o21ai_2 _15824_ (.A1(_07298_),
    .A2(_07299_),
    .B1(_07261_),
    .Y(_07301_));
 sky130_fd_sc_hd__o211a_1 _15825_ (.A1(_07127_),
    .A2(_07167_),
    .B1(_07300_),
    .C1(_07301_),
    .X(_07302_));
 sky130_fd_sc_hd__o211ai_2 _15826_ (.A1(_07127_),
    .A2(_07167_),
    .B1(_07300_),
    .C1(_07301_),
    .Y(_07303_));
 sky130_fd_sc_hd__a211oi_2 _15827_ (.A1(_07300_),
    .A2(_07301_),
    .B1(_07127_),
    .C1(_07167_),
    .Y(_07304_));
 sky130_fd_sc_hd__a22o_1 _15828_ (.A1(net509),
    .A2(net334),
    .B1(net332),
    .B2(net514),
    .X(_07305_));
 sky130_fd_sc_hd__and4_1 _15829_ (.A(net510),
    .B(net513),
    .C(net334),
    .D(net332),
    .X(_07306_));
 sky130_fd_sc_hd__inv_2 _15830_ (.A(_07306_),
    .Y(_07307_));
 sky130_fd_sc_hd__a22oi_1 _15831_ (.A1(net518),
    .A2(net330),
    .B1(_07305_),
    .B2(_07307_),
    .Y(_07308_));
 sky130_fd_sc_hd__and4_1 _15832_ (.A(net518),
    .B(net330),
    .C(_07305_),
    .D(_07307_),
    .X(_07309_));
 sky130_fd_sc_hd__or2_1 _15833_ (.A(_07308_),
    .B(_07309_),
    .X(_07310_));
 sky130_fd_sc_hd__or2_1 _15834_ (.A(_07173_),
    .B(_07176_),
    .X(_07311_));
 sky130_fd_sc_hd__and2b_1 _15835_ (.A_N(_07311_),
    .B(_07310_),
    .X(_07312_));
 sky130_fd_sc_hd__and2b_1 _15836_ (.A_N(_07310_),
    .B(_07311_),
    .X(_07313_));
 sky130_fd_sc_hd__or2_1 _15837_ (.A(_07312_),
    .B(_07313_),
    .X(_07314_));
 sky130_fd_sc_hd__and4b_2 _15838_ (.A_N(net528),
    .B(net327),
    .C(net326),
    .D(net522),
    .X(_07315_));
 sky130_fd_sc_hd__o2bb2a_1 _15839_ (.A1_N(net522),
    .A2_N(net327),
    .B1(_02567_),
    .B2(net529),
    .X(_07316_));
 sky130_fd_sc_hd__o21a_1 _15840_ (.A1(_07315_),
    .A2(_07316_),
    .B1(_07314_),
    .X(_07317_));
 sky130_fd_sc_hd__nor3_1 _15841_ (.A(_07314_),
    .B(_07315_),
    .C(_07316_),
    .Y(_07318_));
 sky130_fd_sc_hd__nor2_1 _15842_ (.A(_07317_),
    .B(_07318_),
    .Y(_07319_));
 sky130_fd_sc_hd__o32ai_4 _15843_ (.A1(_07179_),
    .A2(_07180_),
    .A3(_07182_),
    .B1(_07178_),
    .B2(_07177_),
    .Y(_07320_));
 sky130_fd_sc_hd__xnor2_1 _15844_ (.A(_07319_),
    .B(_07320_),
    .Y(_07321_));
 sky130_fd_sc_hd__nor2_1 _15845_ (.A(_07181_),
    .B(_07321_),
    .Y(_07322_));
 sky130_fd_sc_hd__and2_1 _15846_ (.A(_07181_),
    .B(_07321_),
    .X(_07323_));
 sky130_fd_sc_hd__or2_1 _15847_ (.A(_07322_),
    .B(_07323_),
    .X(_07324_));
 sky130_fd_sc_hd__or2_1 _15848_ (.A(_07195_),
    .B(_07197_),
    .X(_07325_));
 sky130_fd_sc_hd__nand2_1 _15849_ (.A(_07131_),
    .B(_07133_),
    .Y(_07326_));
 sky130_fd_sc_hd__a22o_1 _15850_ (.A1(net496),
    .A2(net347),
    .B1(net343),
    .B2(net500),
    .X(_07327_));
 sky130_fd_sc_hd__inv_2 _15851_ (.A(_07327_),
    .Y(_07328_));
 sky130_fd_sc_hd__and4_1 _15852_ (.A(net500),
    .B(net496),
    .C(net347),
    .D(net343),
    .X(_07329_));
 sky130_fd_sc_hd__o2bb2a_1 _15853_ (.A1_N(net505),
    .A2_N(net338),
    .B1(_07328_),
    .B2(_07329_),
    .X(_07330_));
 sky130_fd_sc_hd__and4b_1 _15854_ (.A_N(_07329_),
    .B(net338),
    .C(net505),
    .D(_07327_),
    .X(_07331_));
 sky130_fd_sc_hd__or2_1 _15855_ (.A(_07330_),
    .B(_07331_),
    .X(_07332_));
 sky130_fd_sc_hd__nand2b_1 _15856_ (.A_N(_07332_),
    .B(_07326_),
    .Y(_07333_));
 sky130_fd_sc_hd__xnor2_1 _15857_ (.A(_07326_),
    .B(_07332_),
    .Y(_07334_));
 sky130_fd_sc_hd__nand2_1 _15858_ (.A(_07325_),
    .B(_07334_),
    .Y(_07335_));
 sky130_fd_sc_hd__or2_1 _15859_ (.A(_07325_),
    .B(_07334_),
    .X(_07336_));
 sky130_fd_sc_hd__nand2_1 _15860_ (.A(_07335_),
    .B(_07336_),
    .Y(_07337_));
 sky130_fd_sc_hd__a21oi_2 _15861_ (.A1(_07142_),
    .A2(_07144_),
    .B1(_07337_),
    .Y(_07338_));
 sky130_fd_sc_hd__and3_1 _15862_ (.A(_07142_),
    .B(_07144_),
    .C(_07337_),
    .X(_07339_));
 sky130_fd_sc_hd__a211oi_2 _15863_ (.A1(_07199_),
    .A2(_07201_),
    .B1(_07338_),
    .C1(_07339_),
    .Y(_07340_));
 sky130_fd_sc_hd__o211a_1 _15864_ (.A1(_07338_),
    .A2(_07339_),
    .B1(_07199_),
    .C1(_07201_),
    .X(_07341_));
 sky130_fd_sc_hd__a211oi_1 _15865_ (.A1(_07204_),
    .A2(_07206_),
    .B1(_07340_),
    .C1(_07341_),
    .Y(_07342_));
 sky130_fd_sc_hd__o211a_1 _15866_ (.A1(_07340_),
    .A2(_07341_),
    .B1(_07204_),
    .C1(_07206_),
    .X(_07343_));
 sky130_fd_sc_hd__or3_1 _15867_ (.A(_07324_),
    .B(_07342_),
    .C(_07343_),
    .X(_07344_));
 sky130_fd_sc_hd__o21ai_1 _15868_ (.A1(_07342_),
    .A2(_07343_),
    .B1(_07324_),
    .Y(_07345_));
 sky130_fd_sc_hd__o211ai_2 _15869_ (.A1(_07163_),
    .A2(_07165_),
    .B1(_07344_),
    .C1(_07345_),
    .Y(_07346_));
 sky130_fd_sc_hd__inv_2 _15870_ (.A(_07346_),
    .Y(_07347_));
 sky130_fd_sc_hd__a211o_1 _15871_ (.A1(_07344_),
    .A2(_07345_),
    .B1(_07163_),
    .C1(_07165_),
    .X(_07348_));
 sky130_fd_sc_hd__o211a_2 _15872_ (.A1(_07208_),
    .A2(_07210_),
    .B1(_07346_),
    .C1(_07348_),
    .X(_07349_));
 sky130_fd_sc_hd__a211oi_1 _15873_ (.A1(_07346_),
    .A2(_07348_),
    .B1(_07208_),
    .C1(_07210_),
    .Y(_07350_));
 sky130_fd_sc_hd__or4_2 _15874_ (.A(_07302_),
    .B(_07304_),
    .C(_07349_),
    .D(_07350_),
    .X(_07351_));
 sky130_fd_sc_hd__o22ai_2 _15875_ (.A1(_07302_),
    .A2(_07304_),
    .B1(_07349_),
    .B2(_07350_),
    .Y(_07352_));
 sky130_fd_sc_hd__o211a_2 _15876_ (.A1(_07169_),
    .A2(_07218_),
    .B1(_07351_),
    .C1(_07352_),
    .X(_07353_));
 sky130_fd_sc_hd__a211oi_2 _15877_ (.A1(_07351_),
    .A2(_07352_),
    .B1(_07169_),
    .C1(_07218_),
    .Y(_07354_));
 sky130_fd_sc_hd__a211oi_4 _15878_ (.A1(_07213_),
    .A2(_07216_),
    .B1(_07353_),
    .C1(_07354_),
    .Y(_07355_));
 sky130_fd_sc_hd__o211a_1 _15879_ (.A1(_07353_),
    .A2(_07354_),
    .B1(_07213_),
    .C1(_07216_),
    .X(_07356_));
 sky130_fd_sc_hd__a211oi_4 _15880_ (.A1(_07221_),
    .A2(_07223_),
    .B1(_07355_),
    .C1(_07356_),
    .Y(_07357_));
 sky130_fd_sc_hd__o211a_1 _15881_ (.A1(_07355_),
    .A2(_07356_),
    .B1(_07221_),
    .C1(_07223_),
    .X(_07358_));
 sky130_fd_sc_hd__a211oi_2 _15882_ (.A1(_07186_),
    .A2(_07189_),
    .B1(_07357_),
    .C1(_07358_),
    .Y(_07359_));
 sky130_fd_sc_hd__o211a_1 _15883_ (.A1(_07357_),
    .A2(_07358_),
    .B1(_07186_),
    .C1(_07189_),
    .X(_07360_));
 sky130_fd_sc_hd__o211a_1 _15884_ (.A1(_07359_),
    .A2(_07360_),
    .B1(_07225_),
    .C1(_07229_),
    .X(_07361_));
 sky130_fd_sc_hd__a211oi_1 _15885_ (.A1(_07225_),
    .A2(_07229_),
    .B1(_07359_),
    .C1(_07360_),
    .Y(_07362_));
 sky130_fd_sc_hd__or2_1 _15886_ (.A(_07361_),
    .B(_07362_),
    .X(_07363_));
 sky130_fd_sc_hd__o21ai_1 _15887_ (.A1(_07234_),
    .A2(_07235_),
    .B1(_07232_),
    .Y(_07364_));
 sky130_fd_sc_hd__xnor2_2 _15888_ (.A(_07363_),
    .B(_07364_),
    .Y(_07365_));
 sky130_fd_sc_hd__a22o_1 _15889_ (.A1(net600),
    .A2(net770),
    .B1(_02711_),
    .B2(net5),
    .X(_07366_));
 sky130_fd_sc_hd__a21o_1 _15890_ (.A1(_03058_),
    .A2(_07365_),
    .B1(_07366_),
    .X(_07367_));
 sky130_fd_sc_hd__mux2_1 _15891_ (.A0(net854),
    .A1(_07367_),
    .S(net2),
    .X(_00293_));
 sky130_fd_sc_hd__and3_1 _15892_ (.A(net398),
    .B(net394),
    .C(net454),
    .X(_07368_));
 sky130_fd_sc_hd__o21ai_1 _15893_ (.A1(net398),
    .A2(net393),
    .B1(net454),
    .Y(_07369_));
 sky130_fd_sc_hd__nor2_2 _15894_ (.A(_07368_),
    .B(_07369_),
    .Y(_07370_));
 sky130_fd_sc_hd__nand2_1 _15895_ (.A(net388),
    .B(net456),
    .Y(_07371_));
 sky130_fd_sc_hd__xor2_1 _15896_ (.A(_07370_),
    .B(_07371_),
    .X(_07372_));
 sky130_fd_sc_hd__nor2_1 _15897_ (.A(_07247_),
    .B(_07372_),
    .Y(_07373_));
 sky130_fd_sc_hd__and2_1 _15898_ (.A(_07247_),
    .B(_07372_),
    .X(_07374_));
 sky130_fd_sc_hd__nor2_1 _15899_ (.A(_07373_),
    .B(_07374_),
    .Y(_07375_));
 sky130_fd_sc_hd__nand2_1 _15900_ (.A(_06985_),
    .B(_07375_),
    .Y(_07376_));
 sky130_fd_sc_hd__or2_1 _15901_ (.A(_06985_),
    .B(_07375_),
    .X(_07377_));
 sky130_fd_sc_hd__and2_1 _15902_ (.A(_07376_),
    .B(_07377_),
    .X(_07378_));
 sky130_fd_sc_hd__o21ai_2 _15903_ (.A1(_07239_),
    .A2(_07248_),
    .B1(_07378_),
    .Y(_07379_));
 sky130_fd_sc_hd__or3_1 _15904_ (.A(_07239_),
    .B(_07248_),
    .C(_07378_),
    .X(_07380_));
 sky130_fd_sc_hd__nand2_2 _15905_ (.A(_07379_),
    .B(_07380_),
    .Y(_07381_));
 sky130_fd_sc_hd__xnor2_1 _15906_ (.A(_06982_),
    .B(_07381_),
    .Y(_07382_));
 sky130_fd_sc_hd__nor3_1 _15907_ (.A(_06980_),
    .B(_07257_),
    .C(_07382_),
    .Y(_07383_));
 sky130_fd_sc_hd__o21a_1 _15908_ (.A1(_06980_),
    .A2(_07257_),
    .B1(_07382_),
    .X(_07384_));
 sky130_fd_sc_hd__or2_1 _15909_ (.A(_07383_),
    .B(_07384_),
    .X(_07385_));
 sky130_fd_sc_hd__a22o_1 _15910_ (.A1(net484),
    .A2(net353),
    .B1(net480),
    .B2(net358),
    .X(_07386_));
 sky130_fd_sc_hd__nand4_1 _15911_ (.A(net358),
    .B(net485),
    .C(net353),
    .D(net480),
    .Y(_07387_));
 sky130_fd_sc_hd__a22o_1 _15912_ (.A1(net488),
    .A2(net349),
    .B1(_07386_),
    .B2(_07387_),
    .X(_07388_));
 sky130_fd_sc_hd__nand4_1 _15913_ (.A(net489),
    .B(net350),
    .C(_07386_),
    .D(_07387_),
    .Y(_07389_));
 sky130_fd_sc_hd__nand2_1 _15914_ (.A(_07388_),
    .B(_07389_),
    .Y(_07390_));
 sky130_fd_sc_hd__a22o_1 _15915_ (.A1(net368),
    .A2(net472),
    .B1(net468),
    .B2(net635),
    .X(_07391_));
 sky130_fd_sc_hd__and4_1 _15916_ (.A(net635),
    .B(net369),
    .C(net472),
    .D(net468),
    .X(_07392_));
 sky130_fd_sc_hd__inv_2 _15917_ (.A(_07392_),
    .Y(_07393_));
 sky130_fd_sc_hd__a22oi_1 _15918_ (.A1(net362),
    .A2(net476),
    .B1(_07391_),
    .B2(_07393_),
    .Y(_07394_));
 sky130_fd_sc_hd__and4_1 _15919_ (.A(net362),
    .B(net476),
    .C(_07391_),
    .D(_07393_),
    .X(_07395_));
 sky130_fd_sc_hd__or2_1 _15920_ (.A(_07394_),
    .B(_07395_),
    .X(_07396_));
 sky130_fd_sc_hd__or2_1 _15921_ (.A(_07268_),
    .B(_07271_),
    .X(_07397_));
 sky130_fd_sc_hd__nand2b_1 _15922_ (.A_N(_07396_),
    .B(_07397_),
    .Y(_07398_));
 sky130_fd_sc_hd__xor2_1 _15923_ (.A(_07396_),
    .B(_07397_),
    .X(_07399_));
 sky130_fd_sc_hd__or2_1 _15924_ (.A(_07390_),
    .B(_07399_),
    .X(_07400_));
 sky130_fd_sc_hd__nand2_1 _15925_ (.A(_07390_),
    .B(_07399_),
    .Y(_07401_));
 sky130_fd_sc_hd__and2_1 _15926_ (.A(_07400_),
    .B(_07401_),
    .X(_07402_));
 sky130_fd_sc_hd__or2_1 _15927_ (.A(_07283_),
    .B(_07285_),
    .X(_07403_));
 sky130_fd_sc_hd__a31o_1 _15928_ (.A1(net388),
    .A2(net458),
    .A3(_07244_),
    .B1(_07243_),
    .X(_07404_));
 sky130_fd_sc_hd__a22o_1 _15929_ (.A1(net378),
    .A2(net462),
    .B1(net458),
    .B2(net384),
    .X(_07405_));
 sky130_fd_sc_hd__inv_2 _15930_ (.A(_07405_),
    .Y(_07406_));
 sky130_fd_sc_hd__and4_1 _15931_ (.A(net384),
    .B(net378),
    .C(net462),
    .D(net458),
    .X(_07407_));
 sky130_fd_sc_hd__o2bb2a_1 _15932_ (.A1_N(net373),
    .A2_N(net465),
    .B1(_07406_),
    .B2(_07407_),
    .X(_07408_));
 sky130_fd_sc_hd__and4b_1 _15933_ (.A_N(_07407_),
    .B(net465),
    .C(net373),
    .D(_07405_),
    .X(_07409_));
 sky130_fd_sc_hd__or2_1 _15934_ (.A(_07408_),
    .B(_07409_),
    .X(_07410_));
 sky130_fd_sc_hd__nand2b_1 _15935_ (.A_N(_07410_),
    .B(_07404_),
    .Y(_07411_));
 sky130_fd_sc_hd__xnor2_1 _15936_ (.A(_07404_),
    .B(_07410_),
    .Y(_07412_));
 sky130_fd_sc_hd__nand2_1 _15937_ (.A(_07403_),
    .B(_07412_),
    .Y(_07413_));
 sky130_fd_sc_hd__xnor2_1 _15938_ (.A(_07403_),
    .B(_07412_),
    .Y(_07414_));
 sky130_fd_sc_hd__a21o_1 _15939_ (.A1(_07287_),
    .A2(_07289_),
    .B1(_07414_),
    .X(_07415_));
 sky130_fd_sc_hd__nand3_1 _15940_ (.A(_07287_),
    .B(_07289_),
    .C(_07414_),
    .Y(_07416_));
 sky130_fd_sc_hd__and3_2 _15941_ (.A(_07402_),
    .B(_07415_),
    .C(_07416_),
    .X(_07417_));
 sky130_fd_sc_hd__inv_2 _15942_ (.A(_07417_),
    .Y(_07418_));
 sky130_fd_sc_hd__a21oi_2 _15943_ (.A1(_07415_),
    .A2(_07416_),
    .B1(_07402_),
    .Y(_07419_));
 sky130_fd_sc_hd__a211oi_4 _15944_ (.A1(_07251_),
    .A2(_07254_),
    .B1(_07417_),
    .C1(_07419_),
    .Y(_07420_));
 sky130_fd_sc_hd__o211a_1 _15945_ (.A1(_07417_),
    .A2(_07419_),
    .B1(_07251_),
    .C1(_07254_),
    .X(_07421_));
 sky130_fd_sc_hd__a211oi_4 _15946_ (.A1(_07291_),
    .A2(_07294_),
    .B1(_07420_),
    .C1(_07421_),
    .Y(_07422_));
 sky130_fd_sc_hd__o211a_1 _15947_ (.A1(_07420_),
    .A2(_07421_),
    .B1(_07291_),
    .C1(_07294_),
    .X(_07423_));
 sky130_fd_sc_hd__nor3_4 _15948_ (.A(_07385_),
    .B(_07422_),
    .C(_07423_),
    .Y(_07424_));
 sky130_fd_sc_hd__o21a_1 _15949_ (.A1(_07422_),
    .A2(_07423_),
    .B1(_07385_),
    .X(_07425_));
 sky130_fd_sc_hd__a211oi_4 _15950_ (.A1(_07260_),
    .A2(_07300_),
    .B1(_07424_),
    .C1(_07425_),
    .Y(_07426_));
 sky130_fd_sc_hd__o211a_1 _15951_ (.A1(_07424_),
    .A2(_07425_),
    .B1(_07260_),
    .C1(_07300_),
    .X(_07427_));
 sky130_fd_sc_hd__nand2b_1 _15952_ (.A_N(_07342_),
    .B(_07344_),
    .Y(_07428_));
 sky130_fd_sc_hd__a22o_1 _15953_ (.A1(net505),
    .A2(\mul0.b[27] ),
    .B1(net331),
    .B2(net510),
    .X(_07429_));
 sky130_fd_sc_hd__and4_1 _15954_ (.A(net505),
    .B(net510),
    .C(net335),
    .D(net331),
    .X(_07430_));
 sky130_fd_sc_hd__inv_2 _15955_ (.A(_07430_),
    .Y(_07431_));
 sky130_fd_sc_hd__a22oi_1 _15956_ (.A1(net513),
    .A2(\mul0.b[29] ),
    .B1(_07429_),
    .B2(_07431_),
    .Y(_07432_));
 sky130_fd_sc_hd__and4_1 _15957_ (.A(net513),
    .B(\mul0.b[29] ),
    .C(_07429_),
    .D(_07431_),
    .X(_07433_));
 sky130_fd_sc_hd__or2_2 _15958_ (.A(_07432_),
    .B(_07433_),
    .X(_07434_));
 sky130_fd_sc_hd__nor2_2 _15959_ (.A(_07306_),
    .B(_07309_),
    .Y(_07435_));
 sky130_fd_sc_hd__xnor2_2 _15960_ (.A(_07434_),
    .B(_07435_),
    .Y(_07436_));
 sky130_fd_sc_hd__and4b_2 _15961_ (.A_N(net523),
    .B(\mul0.b[30] ),
    .C(\mul0.b[31] ),
    .D(net518),
    .X(_07437_));
 sky130_fd_sc_hd__inv_2 _15962_ (.A(_07437_),
    .Y(_07438_));
 sky130_fd_sc_hd__o2bb2a_1 _15963_ (.A1_N(net519),
    .A2_N(\mul0.b[30] ),
    .B1(_02567_),
    .B2(net523),
    .X(_07439_));
 sky130_fd_sc_hd__nor2_1 _15964_ (.A(_07437_),
    .B(_07439_),
    .Y(_07440_));
 sky130_fd_sc_hd__xnor2_1 _15965_ (.A(_07436_),
    .B(_07440_),
    .Y(_07441_));
 sky130_fd_sc_hd__or3_1 _15966_ (.A(_07313_),
    .B(_07318_),
    .C(_07441_),
    .X(_07442_));
 sky130_fd_sc_hd__o21ai_2 _15967_ (.A1(_07313_),
    .A2(_07318_),
    .B1(_07441_),
    .Y(_07443_));
 sky130_fd_sc_hd__nand2_1 _15968_ (.A(_07442_),
    .B(_07443_),
    .Y(_07444_));
 sky130_fd_sc_hd__inv_2 _15969_ (.A(_07444_),
    .Y(_07445_));
 sky130_fd_sc_hd__nand2_1 _15970_ (.A(_07315_),
    .B(_07445_),
    .Y(_07446_));
 sky130_fd_sc_hd__xor2_2 _15971_ (.A(_07315_),
    .B(_07444_),
    .X(_07447_));
 sky130_fd_sc_hd__or2_1 _15972_ (.A(_07329_),
    .B(_07331_),
    .X(_07448_));
 sky130_fd_sc_hd__nand2_1 _15973_ (.A(_07263_),
    .B(_07265_),
    .Y(_07449_));
 sky130_fd_sc_hd__a22o_1 _15974_ (.A1(net492),
    .A2(net347),
    .B1(net343),
    .B2(net496),
    .X(_07450_));
 sky130_fd_sc_hd__inv_2 _15975_ (.A(_07450_),
    .Y(_07451_));
 sky130_fd_sc_hd__and4_1 _15976_ (.A(net496),
    .B(net492),
    .C(net347),
    .D(net342),
    .X(_07452_));
 sky130_fd_sc_hd__o2bb2a_1 _15977_ (.A1_N(net500),
    .A2_N(net338),
    .B1(_07451_),
    .B2(_07452_),
    .X(_07453_));
 sky130_fd_sc_hd__and4b_1 _15978_ (.A_N(_07452_),
    .B(net338),
    .C(net500),
    .D(_07450_),
    .X(_07454_));
 sky130_fd_sc_hd__or2_1 _15979_ (.A(_07453_),
    .B(_07454_),
    .X(_07455_));
 sky130_fd_sc_hd__nand2b_1 _15980_ (.A_N(_07455_),
    .B(_07449_),
    .Y(_07456_));
 sky130_fd_sc_hd__xnor2_1 _15981_ (.A(_07449_),
    .B(_07455_),
    .Y(_07457_));
 sky130_fd_sc_hd__nand2_1 _15982_ (.A(_07448_),
    .B(_07457_),
    .Y(_07458_));
 sky130_fd_sc_hd__xnor2_1 _15983_ (.A(_07448_),
    .B(_07457_),
    .Y(_07459_));
 sky130_fd_sc_hd__a21oi_1 _15984_ (.A1(_07274_),
    .A2(_07276_),
    .B1(_07459_),
    .Y(_07460_));
 sky130_fd_sc_hd__a21o_1 _15985_ (.A1(_07274_),
    .A2(_07276_),
    .B1(_07459_),
    .X(_07461_));
 sky130_fd_sc_hd__and3_1 _15986_ (.A(_07274_),
    .B(_07276_),
    .C(_07459_),
    .X(_07462_));
 sky130_fd_sc_hd__a211o_2 _15987_ (.A1(_07333_),
    .A2(_07335_),
    .B1(_07460_),
    .C1(_07462_),
    .X(_07463_));
 sky130_fd_sc_hd__o211ai_2 _15988_ (.A1(_07460_),
    .A2(_07462_),
    .B1(_07333_),
    .C1(_07335_),
    .Y(_07464_));
 sky130_fd_sc_hd__o211a_1 _15989_ (.A1(_07338_),
    .A2(_07340_),
    .B1(_07463_),
    .C1(_07464_),
    .X(_07465_));
 sky130_fd_sc_hd__a211oi_1 _15990_ (.A1(_07463_),
    .A2(_07464_),
    .B1(_07338_),
    .C1(_07340_),
    .Y(_07466_));
 sky130_fd_sc_hd__or3_2 _15991_ (.A(_07447_),
    .B(_07465_),
    .C(_07466_),
    .X(_07467_));
 sky130_fd_sc_hd__inv_2 _15992_ (.A(_07467_),
    .Y(_07468_));
 sky130_fd_sc_hd__o21ai_2 _15993_ (.A1(_07465_),
    .A2(_07466_),
    .B1(_07447_),
    .Y(_07469_));
 sky130_fd_sc_hd__o211ai_4 _15994_ (.A1(_07296_),
    .A2(_07298_),
    .B1(_07467_),
    .C1(_07469_),
    .Y(_07470_));
 sky130_fd_sc_hd__a211o_1 _15995_ (.A1(_07467_),
    .A2(_07469_),
    .B1(_07296_),
    .C1(_07298_),
    .X(_07471_));
 sky130_fd_sc_hd__and3_1 _15996_ (.A(_07428_),
    .B(_07470_),
    .C(_07471_),
    .X(_07472_));
 sky130_fd_sc_hd__inv_2 _15997_ (.A(_07472_),
    .Y(_07473_));
 sky130_fd_sc_hd__a21oi_1 _15998_ (.A1(_07470_),
    .A2(_07471_),
    .B1(_07428_),
    .Y(_07474_));
 sky130_fd_sc_hd__nor4_2 _15999_ (.A(_07426_),
    .B(_07427_),
    .C(_07472_),
    .D(_07474_),
    .Y(_07475_));
 sky130_fd_sc_hd__o22a_1 _16000_ (.A1(_07426_),
    .A2(_07427_),
    .B1(_07472_),
    .B2(_07474_),
    .X(_07476_));
 sky130_fd_sc_hd__a211o_2 _16001_ (.A1(_07303_),
    .A2(_07351_),
    .B1(_07475_),
    .C1(_07476_),
    .X(_07477_));
 sky130_fd_sc_hd__o211ai_2 _16002_ (.A1(_07475_),
    .A2(_07476_),
    .B1(_07303_),
    .C1(_07351_),
    .Y(_07478_));
 sky130_fd_sc_hd__o211ai_4 _16003_ (.A1(_07347_),
    .A2(_07349_),
    .B1(_07477_),
    .C1(_07478_),
    .Y(_07479_));
 sky130_fd_sc_hd__a211o_1 _16004_ (.A1(_07477_),
    .A2(_07478_),
    .B1(_07347_),
    .C1(_07349_),
    .X(_07480_));
 sky130_fd_sc_hd__o211ai_4 _16005_ (.A1(_07353_),
    .A2(_07355_),
    .B1(_07479_),
    .C1(_07480_),
    .Y(_07481_));
 sky130_fd_sc_hd__a211o_1 _16006_ (.A1(_07479_),
    .A2(_07480_),
    .B1(_07353_),
    .C1(_07355_),
    .X(_07482_));
 sky130_fd_sc_hd__nand2_1 _16007_ (.A(_07481_),
    .B(_07482_),
    .Y(_07483_));
 sky130_fd_sc_hd__a21oi_1 _16008_ (.A1(_07319_),
    .A2(_07320_),
    .B1(_07322_),
    .Y(_07484_));
 sky130_fd_sc_hd__or2_1 _16009_ (.A(_07483_),
    .B(_07484_),
    .X(_07485_));
 sky130_fd_sc_hd__xnor2_1 _16010_ (.A(_07483_),
    .B(_07484_),
    .Y(_07486_));
 sky130_fd_sc_hd__nor2_1 _16011_ (.A(_07357_),
    .B(_07359_),
    .Y(_07487_));
 sky130_fd_sc_hd__or2_1 _16012_ (.A(_07486_),
    .B(_07487_),
    .X(_07488_));
 sky130_fd_sc_hd__inv_2 _16013_ (.A(_07488_),
    .Y(_07489_));
 sky130_fd_sc_hd__nand2_1 _16014_ (.A(_07486_),
    .B(_07487_),
    .Y(_07490_));
 sky130_fd_sc_hd__nand2_1 _16015_ (.A(_07488_),
    .B(_07490_),
    .Y(_07491_));
 sky130_fd_sc_hd__or3_1 _16016_ (.A(_07234_),
    .B(_07361_),
    .C(_07362_),
    .X(_07492_));
 sky130_fd_sc_hd__a2111o_1 _16017_ (.A1(_06973_),
    .A2(_06974_),
    .B1(_07103_),
    .C1(_07492_),
    .D1(_06971_),
    .X(_07493_));
 sky130_fd_sc_hd__o21ai_1 _16018_ (.A1(_06969_),
    .A2(_07101_),
    .B1(_07102_),
    .Y(_07494_));
 sky130_fd_sc_hd__o21ba_1 _16019_ (.A1(_07232_),
    .A2(_07361_),
    .B1_N(_07362_),
    .X(_07495_));
 sky130_fd_sc_hd__o21a_1 _16020_ (.A1(_07492_),
    .A2(_07494_),
    .B1(_07495_),
    .X(_07496_));
 sky130_fd_sc_hd__and3_1 _16021_ (.A(_07491_),
    .B(_07493_),
    .C(_07496_),
    .X(_07497_));
 sky130_fd_sc_hd__a21oi_2 _16022_ (.A1(_07493_),
    .A2(_07496_),
    .B1(_07491_),
    .Y(_07498_));
 sky130_fd_sc_hd__or2_2 _16023_ (.A(_07497_),
    .B(_07498_),
    .X(_07499_));
 sky130_fd_sc_hd__nor2_1 _16024_ (.A(_03057_),
    .B(_07499_),
    .Y(_07500_));
 sky130_fd_sc_hd__a221o_1 _16025_ (.A1(net600),
    .A2(\temp[27] ),
    .B1(_02716_),
    .B2(net5),
    .C1(_07500_),
    .X(_07501_));
 sky130_fd_sc_hd__mux2_1 _16026_ (.A0(net682),
    .A1(_07501_),
    .S(net1),
    .X(_00294_));
 sky130_fd_sc_hd__nand2_1 _16027_ (.A(net388),
    .B(net454),
    .Y(_07502_));
 sky130_fd_sc_hd__xor2_2 _16028_ (.A(_07370_),
    .B(_07502_),
    .X(_07503_));
 sky130_fd_sc_hd__xor2_1 _16029_ (.A(_07247_),
    .B(_07503_),
    .X(_07504_));
 sky130_fd_sc_hd__nand2_1 _16030_ (.A(_06985_),
    .B(_07504_),
    .Y(_07505_));
 sky130_fd_sc_hd__or2_1 _16031_ (.A(_06985_),
    .B(_07504_),
    .X(_07506_));
 sky130_fd_sc_hd__and2_1 _16032_ (.A(_07505_),
    .B(_07506_),
    .X(_07507_));
 sky130_fd_sc_hd__o21ai_2 _16033_ (.A1(_07239_),
    .A2(_07373_),
    .B1(_07507_),
    .Y(_07508_));
 sky130_fd_sc_hd__or3_1 _16034_ (.A(_07239_),
    .B(_07373_),
    .C(_07507_),
    .X(_07509_));
 sky130_fd_sc_hd__nand2_1 _16035_ (.A(_07508_),
    .B(_07509_),
    .Y(_07510_));
 sky130_fd_sc_hd__xnor2_1 _16036_ (.A(_06983_),
    .B(_07510_),
    .Y(_07511_));
 sky130_fd_sc_hd__o21ba_1 _16037_ (.A1(_06983_),
    .A2(_07381_),
    .B1_N(_06980_),
    .X(_07512_));
 sky130_fd_sc_hd__xnor2_1 _16038_ (.A(_07511_),
    .B(_07512_),
    .Y(_07513_));
 sky130_fd_sc_hd__a22o_1 _16039_ (.A1(net354),
    .A2(net480),
    .B1(net475),
    .B2(net359),
    .X(_07514_));
 sky130_fd_sc_hd__nand4_2 _16040_ (.A(net359),
    .B(net354),
    .C(net480),
    .D(net475),
    .Y(_07515_));
 sky130_fd_sc_hd__a22o_1 _16041_ (.A1(net485),
    .A2(net351),
    .B1(_07514_),
    .B2(_07515_),
    .X(_07516_));
 sky130_fd_sc_hd__nand4_1 _16042_ (.A(net485),
    .B(net351),
    .C(_07514_),
    .D(_07515_),
    .Y(_07517_));
 sky130_fd_sc_hd__nand2_1 _16043_ (.A(_07516_),
    .B(_07517_),
    .Y(_07518_));
 sky130_fd_sc_hd__a22o_1 _16044_ (.A1(net368),
    .A2(net468),
    .B1(\mul0.a[27] ),
    .B2(net635),
    .X(_07519_));
 sky130_fd_sc_hd__and4_1 _16045_ (.A(net635),
    .B(net368),
    .C(net468),
    .D(net465),
    .X(_07520_));
 sky130_fd_sc_hd__inv_2 _16046_ (.A(_07520_),
    .Y(_07521_));
 sky130_fd_sc_hd__a22oi_1 _16047_ (.A1(net363),
    .A2(net472),
    .B1(_07519_),
    .B2(_07521_),
    .Y(_07522_));
 sky130_fd_sc_hd__and4_1 _16048_ (.A(net363),
    .B(net472),
    .C(_07519_),
    .D(_07521_),
    .X(_07523_));
 sky130_fd_sc_hd__or2_1 _16049_ (.A(_07522_),
    .B(_07523_),
    .X(_07524_));
 sky130_fd_sc_hd__or2_1 _16050_ (.A(_07392_),
    .B(_07395_),
    .X(_07525_));
 sky130_fd_sc_hd__nand2b_1 _16051_ (.A_N(_07524_),
    .B(_07525_),
    .Y(_07526_));
 sky130_fd_sc_hd__xor2_1 _16052_ (.A(_07524_),
    .B(_07525_),
    .X(_07527_));
 sky130_fd_sc_hd__or2_1 _16053_ (.A(_07518_),
    .B(_07527_),
    .X(_07528_));
 sky130_fd_sc_hd__nand2_1 _16054_ (.A(_07518_),
    .B(_07527_),
    .Y(_07529_));
 sky130_fd_sc_hd__and2_1 _16055_ (.A(_07528_),
    .B(_07529_),
    .X(_07530_));
 sky130_fd_sc_hd__or2_1 _16056_ (.A(_07407_),
    .B(_07409_),
    .X(_07531_));
 sky130_fd_sc_hd__a31o_1 _16057_ (.A1(net388),
    .A2(net455),
    .A3(_07370_),
    .B1(_07368_),
    .X(_07532_));
 sky130_fd_sc_hd__a22o_1 _16058_ (.A1(net379),
    .A2(net458),
    .B1(net455),
    .B2(net385),
    .X(_07533_));
 sky130_fd_sc_hd__and4_1 _16059_ (.A(net385),
    .B(net379),
    .C(net458),
    .D(net455),
    .X(_07534_));
 sky130_fd_sc_hd__inv_2 _16060_ (.A(_07534_),
    .Y(_07535_));
 sky130_fd_sc_hd__a22o_1 _16061_ (.A1(net374),
    .A2(net462),
    .B1(_07533_),
    .B2(_07535_),
    .X(_07536_));
 sky130_fd_sc_hd__and4b_1 _16062_ (.A_N(_07534_),
    .B(net462),
    .C(net374),
    .D(_07533_),
    .X(_07537_));
 sky130_fd_sc_hd__inv_2 _16063_ (.A(_07537_),
    .Y(_07538_));
 sky130_fd_sc_hd__and3_1 _16064_ (.A(_07532_),
    .B(_07536_),
    .C(_07538_),
    .X(_07539_));
 sky130_fd_sc_hd__a21o_1 _16065_ (.A1(_07536_),
    .A2(_07538_),
    .B1(_07532_),
    .X(_07540_));
 sky130_fd_sc_hd__and2b_1 _16066_ (.A_N(_07539_),
    .B(_07540_),
    .X(_07541_));
 sky130_fd_sc_hd__xnor2_1 _16067_ (.A(_07531_),
    .B(_07541_),
    .Y(_07542_));
 sky130_fd_sc_hd__a21o_1 _16068_ (.A1(_07411_),
    .A2(_07413_),
    .B1(_07542_),
    .X(_07543_));
 sky130_fd_sc_hd__nand3_1 _16069_ (.A(_07411_),
    .B(_07413_),
    .C(_07542_),
    .Y(_07544_));
 sky130_fd_sc_hd__and3_1 _16070_ (.A(_07530_),
    .B(_07543_),
    .C(_07544_),
    .X(_07545_));
 sky130_fd_sc_hd__inv_2 _16071_ (.A(_07545_),
    .Y(_07546_));
 sky130_fd_sc_hd__a21oi_1 _16072_ (.A1(_07543_),
    .A2(_07544_),
    .B1(_07530_),
    .Y(_07547_));
 sky130_fd_sc_hd__a211o_1 _16073_ (.A1(_07376_),
    .A2(_07379_),
    .B1(_07545_),
    .C1(_07547_),
    .X(_07548_));
 sky130_fd_sc_hd__o211ai_1 _16074_ (.A1(_07545_),
    .A2(_07547_),
    .B1(_07376_),
    .C1(_07379_),
    .Y(_07549_));
 sky130_fd_sc_hd__nand2_1 _16075_ (.A(_07548_),
    .B(_07549_),
    .Y(_07550_));
 sky130_fd_sc_hd__a21oi_1 _16076_ (.A1(_07415_),
    .A2(_07418_),
    .B1(_07550_),
    .Y(_07551_));
 sky130_fd_sc_hd__a21o_1 _16077_ (.A1(_07415_),
    .A2(_07418_),
    .B1(_07550_),
    .X(_07552_));
 sky130_fd_sc_hd__and3_1 _16078_ (.A(_07415_),
    .B(_07418_),
    .C(_07550_),
    .X(_07553_));
 sky130_fd_sc_hd__or3_2 _16079_ (.A(_07513_),
    .B(_07551_),
    .C(_07553_),
    .X(_07554_));
 sky130_fd_sc_hd__o21ai_2 _16080_ (.A1(_07551_),
    .A2(_07553_),
    .B1(_07513_),
    .Y(_07555_));
 sky130_fd_sc_hd__o211ai_4 _16081_ (.A1(_07384_),
    .A2(_07424_),
    .B1(_07554_),
    .C1(_07555_),
    .Y(_07556_));
 sky130_fd_sc_hd__a211o_1 _16082_ (.A1(_07554_),
    .A2(_07555_),
    .B1(_07384_),
    .C1(_07424_),
    .X(_07557_));
 sky130_fd_sc_hd__a22o_1 _16083_ (.A1(net500),
    .A2(net335),
    .B1(net332),
    .B2(net505),
    .X(_07558_));
 sky130_fd_sc_hd__and4_1 _16084_ (.A(net505),
    .B(net500),
    .C(net335),
    .D(net332),
    .X(_07559_));
 sky130_fd_sc_hd__inv_2 _16085_ (.A(_07559_),
    .Y(_07560_));
 sky130_fd_sc_hd__a22oi_1 _16086_ (.A1(net509),
    .A2(net330),
    .B1(_07558_),
    .B2(_07560_),
    .Y(_07561_));
 sky130_fd_sc_hd__and4_1 _16087_ (.A(net509),
    .B(\mul0.b[29] ),
    .C(_07558_),
    .D(_07560_),
    .X(_07562_));
 sky130_fd_sc_hd__or2_1 _16088_ (.A(_07561_),
    .B(_07562_),
    .X(_07563_));
 sky130_fd_sc_hd__or2_1 _16089_ (.A(_07430_),
    .B(_07433_),
    .X(_07564_));
 sky130_fd_sc_hd__and2b_1 _16090_ (.A_N(_07563_),
    .B(_07564_),
    .X(_07565_));
 sky130_fd_sc_hd__xor2_1 _16091_ (.A(_07563_),
    .B(_07564_),
    .X(_07566_));
 sky130_fd_sc_hd__and4b_2 _16092_ (.A_N(net519),
    .B(\mul0.b[30] ),
    .C(\mul0.b[31] ),
    .D(net513),
    .X(_07567_));
 sky130_fd_sc_hd__o2bb2a_1 _16093_ (.A1_N(net513),
    .A2_N(\mul0.b[30] ),
    .B1(net57),
    .B2(net519),
    .X(_07568_));
 sky130_fd_sc_hd__o21a_1 _16094_ (.A1(_07567_),
    .A2(_07568_),
    .B1(_07566_),
    .X(_07569_));
 sky130_fd_sc_hd__nor3_1 _16095_ (.A(_07566_),
    .B(_07567_),
    .C(_07568_),
    .Y(_07570_));
 sky130_fd_sc_hd__nor2_1 _16096_ (.A(_07569_),
    .B(_07570_),
    .Y(_07571_));
 sky130_fd_sc_hd__o32ai_4 _16097_ (.A1(_07436_),
    .A2(_07437_),
    .A3(_07439_),
    .B1(_07435_),
    .B2(_07434_),
    .Y(_07572_));
 sky130_fd_sc_hd__xnor2_2 _16098_ (.A(_07571_),
    .B(_07572_),
    .Y(_07573_));
 sky130_fd_sc_hd__nor2_1 _16099_ (.A(_07438_),
    .B(_07573_),
    .Y(_07574_));
 sky130_fd_sc_hd__xnor2_2 _16100_ (.A(_07438_),
    .B(_07573_),
    .Y(_07575_));
 sky130_fd_sc_hd__or2_1 _16101_ (.A(_07452_),
    .B(_07454_),
    .X(_07576_));
 sky130_fd_sc_hd__nand2_1 _16102_ (.A(_07387_),
    .B(_07389_),
    .Y(_07577_));
 sky130_fd_sc_hd__a22o_1 _16103_ (.A1(net489),
    .A2(net347),
    .B1(net343),
    .B2(net492),
    .X(_07578_));
 sky130_fd_sc_hd__inv_2 _16104_ (.A(_07578_),
    .Y(_07579_));
 sky130_fd_sc_hd__and4_1 _16105_ (.A(net492),
    .B(net489),
    .C(net347),
    .D(net343),
    .X(_07580_));
 sky130_fd_sc_hd__o2bb2a_1 _16106_ (.A1_N(net496),
    .A2_N(\mul0.b[26] ),
    .B1(_07579_),
    .B2(_07580_),
    .X(_07581_));
 sky130_fd_sc_hd__and4b_1 _16107_ (.A_N(_07580_),
    .B(\mul0.b[26] ),
    .C(net496),
    .D(_07578_),
    .X(_07582_));
 sky130_fd_sc_hd__or2_1 _16108_ (.A(_07581_),
    .B(_07582_),
    .X(_07583_));
 sky130_fd_sc_hd__nand2b_1 _16109_ (.A_N(_07583_),
    .B(_07577_),
    .Y(_07584_));
 sky130_fd_sc_hd__xnor2_1 _16110_ (.A(_07577_),
    .B(_07583_),
    .Y(_07585_));
 sky130_fd_sc_hd__nand2_1 _16111_ (.A(_07576_),
    .B(_07585_),
    .Y(_07586_));
 sky130_fd_sc_hd__xnor2_1 _16112_ (.A(_07576_),
    .B(_07585_),
    .Y(_07587_));
 sky130_fd_sc_hd__a21oi_2 _16113_ (.A1(_07398_),
    .A2(_07400_),
    .B1(_07587_),
    .Y(_07588_));
 sky130_fd_sc_hd__and3_1 _16114_ (.A(_07398_),
    .B(_07400_),
    .C(_07587_),
    .X(_07589_));
 sky130_fd_sc_hd__a211oi_4 _16115_ (.A1(_07456_),
    .A2(_07458_),
    .B1(_07588_),
    .C1(_07589_),
    .Y(_07590_));
 sky130_fd_sc_hd__o211a_1 _16116_ (.A1(_07588_),
    .A2(_07589_),
    .B1(_07456_),
    .C1(_07458_),
    .X(_07591_));
 sky130_fd_sc_hd__a211oi_2 _16117_ (.A1(_07461_),
    .A2(_07463_),
    .B1(_07590_),
    .C1(_07591_),
    .Y(_07592_));
 sky130_fd_sc_hd__o211a_1 _16118_ (.A1(_07590_),
    .A2(_07591_),
    .B1(_07461_),
    .C1(_07463_),
    .X(_07593_));
 sky130_fd_sc_hd__or3_2 _16119_ (.A(_07575_),
    .B(_07592_),
    .C(_07593_),
    .X(_07594_));
 sky130_fd_sc_hd__inv_2 _16120_ (.A(_07594_),
    .Y(_07595_));
 sky130_fd_sc_hd__o21ai_1 _16121_ (.A1(_07592_),
    .A2(_07593_),
    .B1(_07575_),
    .Y(_07596_));
 sky130_fd_sc_hd__o211a_1 _16122_ (.A1(_07420_),
    .A2(_07422_),
    .B1(_07594_),
    .C1(_07596_),
    .X(_07597_));
 sky130_fd_sc_hd__inv_2 _16123_ (.A(_07597_),
    .Y(_07598_));
 sky130_fd_sc_hd__a211o_1 _16124_ (.A1(_07594_),
    .A2(_07596_),
    .B1(_07420_),
    .C1(_07422_),
    .X(_07599_));
 sky130_fd_sc_hd__o211a_1 _16125_ (.A1(_07465_),
    .A2(_07468_),
    .B1(_07598_),
    .C1(_07599_),
    .X(_07600_));
 sky130_fd_sc_hd__a211oi_1 _16126_ (.A1(_07598_),
    .A2(_07599_),
    .B1(_07465_),
    .C1(_07468_),
    .Y(_07601_));
 sky130_fd_sc_hd__nor2_1 _16127_ (.A(_07600_),
    .B(_07601_),
    .Y(_07602_));
 sky130_fd_sc_hd__nand3_2 _16128_ (.A(_07556_),
    .B(_07557_),
    .C(_07602_),
    .Y(_07603_));
 sky130_fd_sc_hd__a21o_1 _16129_ (.A1(_07556_),
    .A2(_07557_),
    .B1(_07602_),
    .X(_07604_));
 sky130_fd_sc_hd__o211a_1 _16130_ (.A1(_07426_),
    .A2(_07475_),
    .B1(_07603_),
    .C1(_07604_),
    .X(_07605_));
 sky130_fd_sc_hd__a211oi_1 _16131_ (.A1(_07603_),
    .A2(_07604_),
    .B1(_07426_),
    .C1(_07475_),
    .Y(_07606_));
 sky130_fd_sc_hd__or2_1 _16132_ (.A(_07605_),
    .B(_07606_),
    .X(_07607_));
 sky130_fd_sc_hd__a21oi_4 _16133_ (.A1(_07470_),
    .A2(_07473_),
    .B1(_07607_),
    .Y(_07608_));
 sky130_fd_sc_hd__and3_1 _16134_ (.A(_07470_),
    .B(_07473_),
    .C(_07607_),
    .X(_07609_));
 sky130_fd_sc_hd__a211oi_4 _16135_ (.A1(_07477_),
    .A2(_07479_),
    .B1(_07608_),
    .C1(_07609_),
    .Y(_07610_));
 sky130_fd_sc_hd__o211a_1 _16136_ (.A1(_07608_),
    .A2(_07609_),
    .B1(_07477_),
    .C1(_07479_),
    .X(_07611_));
 sky130_fd_sc_hd__a211oi_4 _16137_ (.A1(_07443_),
    .A2(_07446_),
    .B1(_07610_),
    .C1(_07611_),
    .Y(_07612_));
 sky130_fd_sc_hd__o211a_1 _16138_ (.A1(_07610_),
    .A2(_07611_),
    .B1(_07443_),
    .C1(_07446_),
    .X(_07613_));
 sky130_fd_sc_hd__a211oi_4 _16139_ (.A1(_07481_),
    .A2(_07485_),
    .B1(_07612_),
    .C1(_07613_),
    .Y(_07614_));
 sky130_fd_sc_hd__o211a_1 _16140_ (.A1(_07612_),
    .A2(_07613_),
    .B1(_07481_),
    .C1(_07485_),
    .X(_07615_));
 sky130_fd_sc_hd__inv_2 _16141_ (.A(_07615_),
    .Y(_07616_));
 sky130_fd_sc_hd__nor2_1 _16142_ (.A(_07614_),
    .B(_07615_),
    .Y(_07617_));
 sky130_fd_sc_hd__or2_1 _16143_ (.A(_07489_),
    .B(_07498_),
    .X(_07618_));
 sky130_fd_sc_hd__xnor2_2 _16144_ (.A(_07617_),
    .B(_07618_),
    .Y(_07619_));
 sky130_fd_sc_hd__nor2_1 _16145_ (.A(_03057_),
    .B(_07619_),
    .Y(_07620_));
 sky130_fd_sc_hd__a221o_1 _16146_ (.A1(net600),
    .A2(net723),
    .B1(_02722_),
    .B2(net5),
    .C1(_07620_),
    .X(_07621_));
 sky130_fd_sc_hd__mux2_1 _16147_ (.A0(net722),
    .A1(_07621_),
    .S(net1),
    .X(_00295_));
 sky130_fd_sc_hd__o21ba_1 _16148_ (.A1(_06983_),
    .A2(_07510_),
    .B1_N(_06980_),
    .X(_07622_));
 sky130_fd_sc_hd__o21ai_4 _16149_ (.A1(_07247_),
    .A2(_07503_),
    .B1(_07240_),
    .Y(_07623_));
 sky130_fd_sc_hd__xor2_2 _16150_ (.A(_07507_),
    .B(_07623_),
    .X(_07624_));
 sky130_fd_sc_hd__xnor2_1 _16151_ (.A(_06982_),
    .B(_07624_),
    .Y(_07625_));
 sky130_fd_sc_hd__xnor2_1 _16152_ (.A(_07622_),
    .B(_07625_),
    .Y(_07626_));
 sky130_fd_sc_hd__a22o_1 _16153_ (.A1(net354),
    .A2(net475),
    .B1(net471),
    .B2(net359),
    .X(_07627_));
 sky130_fd_sc_hd__and4_1 _16154_ (.A(net359),
    .B(net354),
    .C(net475),
    .D(net471),
    .X(_07628_));
 sky130_fd_sc_hd__inv_2 _16155_ (.A(_07628_),
    .Y(_07629_));
 sky130_fd_sc_hd__a22oi_1 _16156_ (.A1(net479),
    .A2(net351),
    .B1(_07627_),
    .B2(_07629_),
    .Y(_07630_));
 sky130_fd_sc_hd__and4_1 _16157_ (.A(net479),
    .B(net351),
    .C(_07627_),
    .D(_07629_),
    .X(_07631_));
 sky130_fd_sc_hd__or2_1 _16158_ (.A(_07630_),
    .B(_07631_),
    .X(_07632_));
 sky130_fd_sc_hd__a22o_1 _16159_ (.A1(net368),
    .A2(net465),
    .B1(\mul0.a[28] ),
    .B2(net635),
    .X(_07633_));
 sky130_fd_sc_hd__and4_1 _16160_ (.A(net635),
    .B(net368),
    .C(\mul0.a[27] ),
    .D(net462),
    .X(_07634_));
 sky130_fd_sc_hd__inv_2 _16161_ (.A(_07634_),
    .Y(_07635_));
 sky130_fd_sc_hd__a22oi_1 _16162_ (.A1(net363),
    .A2(net469),
    .B1(_07633_),
    .B2(_07635_),
    .Y(_07636_));
 sky130_fd_sc_hd__and4_1 _16163_ (.A(net363),
    .B(net468),
    .C(_07633_),
    .D(_07635_),
    .X(_07637_));
 sky130_fd_sc_hd__or2_1 _16164_ (.A(_07636_),
    .B(_07637_),
    .X(_07638_));
 sky130_fd_sc_hd__or2_1 _16165_ (.A(_07520_),
    .B(_07523_),
    .X(_07639_));
 sky130_fd_sc_hd__nand2b_1 _16166_ (.A_N(_07638_),
    .B(_07639_),
    .Y(_07640_));
 sky130_fd_sc_hd__xor2_1 _16167_ (.A(_07638_),
    .B(_07639_),
    .X(_07641_));
 sky130_fd_sc_hd__or2_1 _16168_ (.A(_07632_),
    .B(_07641_),
    .X(_07642_));
 sky130_fd_sc_hd__nand2_1 _16169_ (.A(_07632_),
    .B(_07641_),
    .Y(_07643_));
 sky130_fd_sc_hd__and2_1 _16170_ (.A(_07642_),
    .B(_07643_),
    .X(_07644_));
 sky130_fd_sc_hd__or2_1 _16171_ (.A(_07534_),
    .B(_07537_),
    .X(_07645_));
 sky130_fd_sc_hd__o21ba_1 _16172_ (.A1(_07369_),
    .A2(_07502_),
    .B1_N(_07368_),
    .X(_07646_));
 sky130_fd_sc_hd__and2_1 _16173_ (.A(net385),
    .B(net453),
    .X(_07647_));
 sky130_fd_sc_hd__a21oi_1 _16174_ (.A1(net379),
    .A2(net455),
    .B1(_07647_),
    .Y(_07648_));
 sky130_fd_sc_hd__and3_1 _16175_ (.A(net379),
    .B(net455),
    .C(_07647_),
    .X(_07649_));
 sky130_fd_sc_hd__or2_1 _16176_ (.A(_07648_),
    .B(_07649_),
    .X(_07650_));
 sky130_fd_sc_hd__nand2_1 _16177_ (.A(net374),
    .B(net458),
    .Y(_07651_));
 sky130_fd_sc_hd__xnor2_1 _16178_ (.A(_07650_),
    .B(_07651_),
    .Y(_07652_));
 sky130_fd_sc_hd__or2_1 _16179_ (.A(_07646_),
    .B(_07652_),
    .X(_07653_));
 sky130_fd_sc_hd__xor2_1 _16180_ (.A(_07646_),
    .B(_07652_),
    .X(_07654_));
 sky130_fd_sc_hd__xnor2_1 _16181_ (.A(_07645_),
    .B(_07654_),
    .Y(_07655_));
 sky130_fd_sc_hd__a21oi_1 _16182_ (.A1(_07531_),
    .A2(_07541_),
    .B1(_07539_),
    .Y(_07656_));
 sky130_fd_sc_hd__xor2_1 _16183_ (.A(_07655_),
    .B(_07656_),
    .X(_07657_));
 sky130_fd_sc_hd__and2_1 _16184_ (.A(_07644_),
    .B(_07657_),
    .X(_07658_));
 sky130_fd_sc_hd__nor2_1 _16185_ (.A(_07644_),
    .B(_07657_),
    .Y(_07659_));
 sky130_fd_sc_hd__a211oi_2 _16186_ (.A1(_07505_),
    .A2(_07508_),
    .B1(_07658_),
    .C1(_07659_),
    .Y(_07660_));
 sky130_fd_sc_hd__o211a_1 _16187_ (.A1(_07658_),
    .A2(_07659_),
    .B1(_07505_),
    .C1(_07508_),
    .X(_07661_));
 sky130_fd_sc_hd__a211oi_2 _16188_ (.A1(_07543_),
    .A2(_07546_),
    .B1(_07660_),
    .C1(_07661_),
    .Y(_07662_));
 sky130_fd_sc_hd__o211a_1 _16189_ (.A1(_07660_),
    .A2(_07661_),
    .B1(_07543_),
    .C1(_07546_),
    .X(_07663_));
 sky130_fd_sc_hd__o21ai_2 _16190_ (.A1(_07662_),
    .A2(_07663_),
    .B1(_07626_),
    .Y(_07664_));
 sky130_fd_sc_hd__or3_2 _16191_ (.A(_07626_),
    .B(_07662_),
    .C(_07663_),
    .X(_07665_));
 sky130_fd_sc_hd__o21ai_1 _16192_ (.A1(_07511_),
    .A2(_07512_),
    .B1(_07554_),
    .Y(_07666_));
 sky130_fd_sc_hd__and3_1 _16193_ (.A(_07664_),
    .B(_07665_),
    .C(_07666_),
    .X(_07667_));
 sky130_fd_sc_hd__a21oi_1 _16194_ (.A1(_07664_),
    .A2(_07665_),
    .B1(_07666_),
    .Y(_07668_));
 sky130_fd_sc_hd__a22o_1 _16195_ (.A1(net496),
    .A2(net336),
    .B1(net333),
    .B2(net500),
    .X(_07669_));
 sky130_fd_sc_hd__and4_1 _16196_ (.A(net500),
    .B(net496),
    .C(net336),
    .D(net333),
    .X(_07670_));
 sky130_fd_sc_hd__inv_2 _16197_ (.A(_07670_),
    .Y(_07671_));
 sky130_fd_sc_hd__a22oi_1 _16198_ (.A1(net506),
    .A2(net330),
    .B1(_07669_),
    .B2(_07671_),
    .Y(_07672_));
 sky130_fd_sc_hd__and4_1 _16199_ (.A(net506),
    .B(net330),
    .C(_07669_),
    .D(_07671_),
    .X(_07673_));
 sky130_fd_sc_hd__or2_2 _16200_ (.A(_07672_),
    .B(_07673_),
    .X(_07674_));
 sky130_fd_sc_hd__nor2_2 _16201_ (.A(_07559_),
    .B(_07562_),
    .Y(_07675_));
 sky130_fd_sc_hd__xnor2_4 _16202_ (.A(_07674_),
    .B(_07675_),
    .Y(_07676_));
 sky130_fd_sc_hd__and4b_2 _16203_ (.A_N(net514),
    .B(net328),
    .C(net326),
    .D(net510),
    .X(_07677_));
 sky130_fd_sc_hd__o2bb2a_1 _16204_ (.A1_N(net510),
    .A2_N(net328),
    .B1(net57),
    .B2(net514),
    .X(_07678_));
 sky130_fd_sc_hd__nor2_1 _16205_ (.A(_07677_),
    .B(_07678_),
    .Y(_07679_));
 sky130_fd_sc_hd__xnor2_2 _16206_ (.A(_07676_),
    .B(_07679_),
    .Y(_07680_));
 sky130_fd_sc_hd__nor3_1 _16207_ (.A(_07565_),
    .B(_07570_),
    .C(_07680_),
    .Y(_07681_));
 sky130_fd_sc_hd__o21a_1 _16208_ (.A1(_07565_),
    .A2(_07570_),
    .B1(_07680_),
    .X(_07682_));
 sky130_fd_sc_hd__or2_1 _16209_ (.A(_07681_),
    .B(_07682_),
    .X(_07683_));
 sky130_fd_sc_hd__inv_2 _16210_ (.A(_07683_),
    .Y(_07684_));
 sky130_fd_sc_hd__xor2_2 _16211_ (.A(_07567_),
    .B(_07683_),
    .X(_07685_));
 sky130_fd_sc_hd__or2_1 _16212_ (.A(_07580_),
    .B(_07582_),
    .X(_07686_));
 sky130_fd_sc_hd__nand2_1 _16213_ (.A(_07515_),
    .B(_07517_),
    .Y(_07687_));
 sky130_fd_sc_hd__a22o_1 _16214_ (.A1(net484),
    .A2(net347),
    .B1(net343),
    .B2(net488),
    .X(_07688_));
 sky130_fd_sc_hd__and4_1 _16215_ (.A(net488),
    .B(net484),
    .C(net347),
    .D(net343),
    .X(_07689_));
 sky130_fd_sc_hd__inv_2 _16216_ (.A(_07689_),
    .Y(_07690_));
 sky130_fd_sc_hd__a22oi_1 _16217_ (.A1(net493),
    .A2(\mul0.b[26] ),
    .B1(_07688_),
    .B2(_07690_),
    .Y(_07691_));
 sky130_fd_sc_hd__and4_1 _16218_ (.A(net493),
    .B(net337),
    .C(_07688_),
    .D(_07690_),
    .X(_07692_));
 sky130_fd_sc_hd__or2_1 _16219_ (.A(_07691_),
    .B(_07692_),
    .X(_07693_));
 sky130_fd_sc_hd__nand2b_1 _16220_ (.A_N(_07693_),
    .B(_07687_),
    .Y(_07694_));
 sky130_fd_sc_hd__xnor2_1 _16221_ (.A(_07687_),
    .B(_07693_),
    .Y(_07695_));
 sky130_fd_sc_hd__nand2_1 _16222_ (.A(_07686_),
    .B(_07695_),
    .Y(_07696_));
 sky130_fd_sc_hd__or2_1 _16223_ (.A(_07686_),
    .B(_07695_),
    .X(_07697_));
 sky130_fd_sc_hd__nand2_1 _16224_ (.A(_07696_),
    .B(_07697_),
    .Y(_07698_));
 sky130_fd_sc_hd__a21oi_2 _16225_ (.A1(_07526_),
    .A2(_07528_),
    .B1(_07698_),
    .Y(_07699_));
 sky130_fd_sc_hd__and3_1 _16226_ (.A(_07526_),
    .B(_07528_),
    .C(_07698_),
    .X(_07700_));
 sky130_fd_sc_hd__a211oi_1 _16227_ (.A1(_07584_),
    .A2(_07586_),
    .B1(_07699_),
    .C1(_07700_),
    .Y(_07701_));
 sky130_fd_sc_hd__a211o_1 _16228_ (.A1(_07584_),
    .A2(_07586_),
    .B1(_07699_),
    .C1(_07700_),
    .X(_07702_));
 sky130_fd_sc_hd__o211ai_2 _16229_ (.A1(_07699_),
    .A2(_07700_),
    .B1(_07584_),
    .C1(_07586_),
    .Y(_07703_));
 sky130_fd_sc_hd__o211a_1 _16230_ (.A1(_07588_),
    .A2(_07590_),
    .B1(_07702_),
    .C1(_07703_),
    .X(_07704_));
 sky130_fd_sc_hd__a211oi_1 _16231_ (.A1(_07702_),
    .A2(_07703_),
    .B1(_07588_),
    .C1(_07590_),
    .Y(_07705_));
 sky130_fd_sc_hd__nor3_1 _16232_ (.A(_07685_),
    .B(_07704_),
    .C(_07705_),
    .Y(_07706_));
 sky130_fd_sc_hd__o21a_1 _16233_ (.A1(_07704_),
    .A2(_07705_),
    .B1(_07685_),
    .X(_07707_));
 sky130_fd_sc_hd__a211o_1 _16234_ (.A1(_07548_),
    .A2(_07552_),
    .B1(_07706_),
    .C1(_07707_),
    .X(_07708_));
 sky130_fd_sc_hd__inv_2 _16235_ (.A(_07708_),
    .Y(_07709_));
 sky130_fd_sc_hd__o211a_1 _16236_ (.A1(_07706_),
    .A2(_07707_),
    .B1(_07548_),
    .C1(_07552_),
    .X(_07710_));
 sky130_fd_sc_hd__inv_2 _16237_ (.A(_07710_),
    .Y(_07711_));
 sky130_fd_sc_hd__o211a_1 _16238_ (.A1(_07592_),
    .A2(_07595_),
    .B1(_07708_),
    .C1(_07711_),
    .X(_07712_));
 sky130_fd_sc_hd__a211oi_2 _16239_ (.A1(_07708_),
    .A2(_07711_),
    .B1(_07592_),
    .C1(_07595_),
    .Y(_07713_));
 sky130_fd_sc_hd__nor4_2 _16240_ (.A(_07667_),
    .B(_07668_),
    .C(_07712_),
    .D(_07713_),
    .Y(_07714_));
 sky130_fd_sc_hd__o22a_1 _16241_ (.A1(_07667_),
    .A2(_07668_),
    .B1(_07712_),
    .B2(_07713_),
    .X(_07715_));
 sky130_fd_sc_hd__a211o_1 _16242_ (.A1(_07556_),
    .A2(_07603_),
    .B1(_07714_),
    .C1(_07715_),
    .X(_07716_));
 sky130_fd_sc_hd__o211ai_2 _16243_ (.A1(_07714_),
    .A2(_07715_),
    .B1(_07556_),
    .C1(_07603_),
    .Y(_07717_));
 sky130_fd_sc_hd__o211ai_2 _16244_ (.A1(_07597_),
    .A2(_07600_),
    .B1(_07716_),
    .C1(_07717_),
    .Y(_07718_));
 sky130_fd_sc_hd__a211o_1 _16245_ (.A1(_07716_),
    .A2(_07717_),
    .B1(_07597_),
    .C1(_07600_),
    .X(_07719_));
 sky130_fd_sc_hd__o211ai_2 _16246_ (.A1(_07605_),
    .A2(_07608_),
    .B1(_07718_),
    .C1(_07719_),
    .Y(_07720_));
 sky130_fd_sc_hd__a211o_1 _16247_ (.A1(_07718_),
    .A2(_07719_),
    .B1(_07605_),
    .C1(_07608_),
    .X(_07721_));
 sky130_fd_sc_hd__nand2_1 _16248_ (.A(_07720_),
    .B(_07721_),
    .Y(_07722_));
 sky130_fd_sc_hd__a21oi_2 _16249_ (.A1(_07571_),
    .A2(_07572_),
    .B1(_07574_),
    .Y(_07723_));
 sky130_fd_sc_hd__xnor2_2 _16250_ (.A(_07722_),
    .B(_07723_),
    .Y(_07724_));
 sky130_fd_sc_hd__or2_1 _16251_ (.A(_07610_),
    .B(_07612_),
    .X(_07725_));
 sky130_fd_sc_hd__and2b_1 _16252_ (.A_N(_07724_),
    .B(_07725_),
    .X(_07726_));
 sky130_fd_sc_hd__xnor2_2 _16253_ (.A(_07724_),
    .B(_07725_),
    .Y(_07727_));
 sky130_fd_sc_hd__o31ai_2 _16254_ (.A1(_07489_),
    .A2(_07498_),
    .A3(_07614_),
    .B1(_07616_),
    .Y(_07728_));
 sky130_fd_sc_hd__o311a_1 _16255_ (.A1(_07489_),
    .A2(_07498_),
    .A3(_07614_),
    .B1(_07616_),
    .C1(_07727_),
    .X(_07729_));
 sky130_fd_sc_hd__xor2_2 _16256_ (.A(_07727_),
    .B(_07728_),
    .X(_07730_));
 sky130_fd_sc_hd__nor2_1 _16257_ (.A(_03057_),
    .B(_07730_),
    .Y(_07731_));
 sky130_fd_sc_hd__a221o_1 _16258_ (.A1(net600),
    .A2(\temp[29] ),
    .B1(_02727_),
    .B2(net5),
    .C1(_07731_),
    .X(_07732_));
 sky130_fd_sc_hd__mux2_1 _16259_ (.A0(net774),
    .A1(_07732_),
    .S(net1),
    .X(_00296_));
 sky130_fd_sc_hd__o21ai_1 _16260_ (.A1(_07622_),
    .A2(_07625_),
    .B1(_07665_),
    .Y(_07733_));
 sky130_fd_sc_hd__and2b_1 _16261_ (.A_N(_07624_),
    .B(_06981_),
    .X(_07734_));
 sky130_fd_sc_hd__a21o_1 _16262_ (.A1(_06980_),
    .A2(_07624_),
    .B1(_07734_),
    .X(_07735_));
 sky130_fd_sc_hd__o21ba_1 _16263_ (.A1(_07655_),
    .A2(_07656_),
    .B1_N(_07658_),
    .X(_07736_));
 sky130_fd_sc_hd__a21boi_4 _16264_ (.A1(_07506_),
    .A2(_07623_),
    .B1_N(_07505_),
    .Y(_07737_));
 sky130_fd_sc_hd__a22o_1 _16265_ (.A1(net354),
    .A2(net471),
    .B1(net468),
    .B2(net359),
    .X(_07738_));
 sky130_fd_sc_hd__and3_1 _16266_ (.A(net359),
    .B(net354),
    .C(net471),
    .X(_07739_));
 sky130_fd_sc_hd__a21bo_1 _16267_ (.A1(net468),
    .A2(_07739_),
    .B1_N(_07738_),
    .X(_07740_));
 sky130_fd_sc_hd__nand2_1 _16268_ (.A(net351),
    .B(net475),
    .Y(_07741_));
 sky130_fd_sc_hd__xnor2_1 _16269_ (.A(_07740_),
    .B(_07741_),
    .Y(_07742_));
 sky130_fd_sc_hd__a22o_1 _16270_ (.A1(net368),
    .A2(net462),
    .B1(\mul0.a[29] ),
    .B2(net635),
    .X(_07743_));
 sky130_fd_sc_hd__and3_1 _16271_ (.A(net635),
    .B(net368),
    .C(net462),
    .X(_07744_));
 sky130_fd_sc_hd__a21bo_1 _16272_ (.A1(net458),
    .A2(_07744_),
    .B1_N(_07743_),
    .X(_07745_));
 sky130_fd_sc_hd__nand2_1 _16273_ (.A(net363),
    .B(net465),
    .Y(_07746_));
 sky130_fd_sc_hd__xnor2_1 _16274_ (.A(_07745_),
    .B(_07746_),
    .Y(_07747_));
 sky130_fd_sc_hd__or2_1 _16275_ (.A(_07634_),
    .B(_07637_),
    .X(_07748_));
 sky130_fd_sc_hd__nand2b_1 _16276_ (.A_N(_07747_),
    .B(_07748_),
    .Y(_07749_));
 sky130_fd_sc_hd__xor2_1 _16277_ (.A(_07747_),
    .B(_07748_),
    .X(_07750_));
 sky130_fd_sc_hd__xor2_1 _16278_ (.A(_07742_),
    .B(_07750_),
    .X(_07751_));
 sky130_fd_sc_hd__inv_2 _16279_ (.A(_07751_),
    .Y(_07752_));
 sky130_fd_sc_hd__a21bo_1 _16280_ (.A1(_07645_),
    .A2(_07654_),
    .B1_N(_07653_),
    .X(_07753_));
 sky130_fd_sc_hd__o21ba_1 _16281_ (.A1(_07648_),
    .A2(_07651_),
    .B1_N(_07649_),
    .X(_07754_));
 sky130_fd_sc_hd__o21ai_1 _16282_ (.A1(net385),
    .A2(net379),
    .B1(net454),
    .Y(_07755_));
 sky130_fd_sc_hd__inv_2 _16283_ (.A(_07755_),
    .Y(_07756_));
 sky130_fd_sc_hd__nand2_1 _16284_ (.A(net379),
    .B(_07647_),
    .Y(_07757_));
 sky130_fd_sc_hd__a22o_1 _16285_ (.A1(net374),
    .A2(net455),
    .B1(_07756_),
    .B2(_07757_),
    .X(_07758_));
 sky130_fd_sc_hd__nand4_1 _16286_ (.A(net374),
    .B(net455),
    .C(_07756_),
    .D(_07757_),
    .Y(_07759_));
 sky130_fd_sc_hd__and3_1 _16287_ (.A(_07646_),
    .B(_07758_),
    .C(_07759_),
    .X(_07760_));
 sky130_fd_sc_hd__a21oi_1 _16288_ (.A1(_07758_),
    .A2(_07759_),
    .B1(_07646_),
    .Y(_07761_));
 sky130_fd_sc_hd__nor2_1 _16289_ (.A(_07760_),
    .B(_07761_),
    .Y(_07762_));
 sky130_fd_sc_hd__xor2_1 _16290_ (.A(_07754_),
    .B(_07762_),
    .X(_07763_));
 sky130_fd_sc_hd__xnor2_1 _16291_ (.A(_07753_),
    .B(_07763_),
    .Y(_07764_));
 sky130_fd_sc_hd__nor2_1 _16292_ (.A(_07752_),
    .B(_07764_),
    .Y(_07765_));
 sky130_fd_sc_hd__and2_1 _16293_ (.A(_07752_),
    .B(_07764_),
    .X(_07766_));
 sky130_fd_sc_hd__nor2_1 _16294_ (.A(_07765_),
    .B(_07766_),
    .Y(_07767_));
 sky130_fd_sc_hd__xnor2_1 _16295_ (.A(_07737_),
    .B(_07767_),
    .Y(_07768_));
 sky130_fd_sc_hd__nand2b_1 _16296_ (.A_N(_07736_),
    .B(_07768_),
    .Y(_07769_));
 sky130_fd_sc_hd__xnor2_1 _16297_ (.A(_07736_),
    .B(_07768_),
    .Y(_07770_));
 sky130_fd_sc_hd__xnor2_1 _16298_ (.A(_07735_),
    .B(_07770_),
    .Y(_07771_));
 sky130_fd_sc_hd__and2_1 _16299_ (.A(_07733_),
    .B(_07771_),
    .X(_07772_));
 sky130_fd_sc_hd__nor2_1 _16300_ (.A(_07733_),
    .B(_07771_),
    .Y(_07773_));
 sky130_fd_sc_hd__nor2_1 _16301_ (.A(_07772_),
    .B(_07773_),
    .Y(_07774_));
 sky130_fd_sc_hd__or2_1 _16302_ (.A(_07704_),
    .B(_07706_),
    .X(_07775_));
 sky130_fd_sc_hd__nor2_1 _16303_ (.A(_07660_),
    .B(_07662_),
    .Y(_07776_));
 sky130_fd_sc_hd__a22oi_1 _16304_ (.A1(net492),
    .A2(net336),
    .B1(net333),
    .B2(net497),
    .Y(_07777_));
 sky130_fd_sc_hd__and4_1 _16305_ (.A(net497),
    .B(net492),
    .C(net336),
    .D(net333),
    .X(_07778_));
 sky130_fd_sc_hd__nor2_1 _16306_ (.A(_07777_),
    .B(_07778_),
    .Y(_07779_));
 sky130_fd_sc_hd__nand2_1 _16307_ (.A(net502),
    .B(net330),
    .Y(_07780_));
 sky130_fd_sc_hd__xor2_1 _16308_ (.A(_07779_),
    .B(_07780_),
    .X(_07781_));
 sky130_fd_sc_hd__or2_1 _16309_ (.A(_07670_),
    .B(_07673_),
    .X(_07782_));
 sky130_fd_sc_hd__and2b_1 _16310_ (.A_N(_07782_),
    .B(_07781_),
    .X(_07783_));
 sky130_fd_sc_hd__and2b_1 _16311_ (.A_N(_07781_),
    .B(_07782_),
    .X(_07784_));
 sky130_fd_sc_hd__nor2_1 _16312_ (.A(_07783_),
    .B(_07784_),
    .Y(_07785_));
 sky130_fd_sc_hd__a22o_1 _16313_ (.A1(net506),
    .A2(net328),
    .B1(net326),
    .B2(_02563_),
    .X(_07786_));
 sky130_fd_sc_hd__nand4_2 _16314_ (.A(net506),
    .B(_02563_),
    .C(net328),
    .D(net326),
    .Y(_07787_));
 sky130_fd_sc_hd__nand2_1 _16315_ (.A(_07786_),
    .B(_07787_),
    .Y(_07788_));
 sky130_fd_sc_hd__xnor2_2 _16316_ (.A(_07785_),
    .B(_07788_),
    .Y(_07789_));
 sky130_fd_sc_hd__o32ai_4 _16317_ (.A1(_07676_),
    .A2(_07677_),
    .A3(_07678_),
    .B1(_07675_),
    .B2(_07674_),
    .Y(_07790_));
 sky130_fd_sc_hd__and2_1 _16318_ (.A(_07789_),
    .B(_07790_),
    .X(_07791_));
 sky130_fd_sc_hd__xnor2_2 _16319_ (.A(_07789_),
    .B(_07790_),
    .Y(_07792_));
 sky130_fd_sc_hd__inv_2 _16320_ (.A(_07792_),
    .Y(_07793_));
 sky130_fd_sc_hd__xor2_2 _16321_ (.A(_07677_),
    .B(_07792_),
    .X(_07794_));
 sky130_fd_sc_hd__nand2_1 _16322_ (.A(_07640_),
    .B(_07642_),
    .Y(_07795_));
 sky130_fd_sc_hd__or2_1 _16323_ (.A(_07689_),
    .B(_07692_),
    .X(_07796_));
 sky130_fd_sc_hd__nor2_1 _16324_ (.A(_07628_),
    .B(_07631_),
    .Y(_07797_));
 sky130_fd_sc_hd__a22oi_1 _16325_ (.A1(net479),
    .A2(net347),
    .B1(net343),
    .B2(net484),
    .Y(_07798_));
 sky130_fd_sc_hd__and4_1 _16326_ (.A(net484),
    .B(net479),
    .C(net347),
    .D(net343),
    .X(_07799_));
 sky130_fd_sc_hd__nor2_1 _16327_ (.A(_07798_),
    .B(_07799_),
    .Y(_07800_));
 sky130_fd_sc_hd__nand2_1 _16328_ (.A(net488),
    .B(net337),
    .Y(_07801_));
 sky130_fd_sc_hd__xor2_1 _16329_ (.A(_07800_),
    .B(_07801_),
    .X(_07802_));
 sky130_fd_sc_hd__nor2_1 _16330_ (.A(_07797_),
    .B(_07802_),
    .Y(_07803_));
 sky130_fd_sc_hd__nand2_1 _16331_ (.A(_07797_),
    .B(_07802_),
    .Y(_07804_));
 sky130_fd_sc_hd__and2b_1 _16332_ (.A_N(_07803_),
    .B(_07804_),
    .X(_07805_));
 sky130_fd_sc_hd__xnor2_1 _16333_ (.A(_07796_),
    .B(_07805_),
    .Y(_07806_));
 sky130_fd_sc_hd__nand2b_1 _16334_ (.A_N(_07806_),
    .B(_07795_),
    .Y(_07807_));
 sky130_fd_sc_hd__xor2_1 _16335_ (.A(_07795_),
    .B(_07806_),
    .X(_07808_));
 sky130_fd_sc_hd__a21o_1 _16336_ (.A1(_07694_),
    .A2(_07696_),
    .B1(_07808_),
    .X(_07809_));
 sky130_fd_sc_hd__nand3_1 _16337_ (.A(_07694_),
    .B(_07696_),
    .C(_07808_),
    .Y(_07810_));
 sky130_fd_sc_hd__o211a_1 _16338_ (.A1(_07699_),
    .A2(_07701_),
    .B1(_07809_),
    .C1(_07810_),
    .X(_07811_));
 sky130_fd_sc_hd__a211oi_1 _16339_ (.A1(_07809_),
    .A2(_07810_),
    .B1(_07699_),
    .C1(_07701_),
    .Y(_07812_));
 sky130_fd_sc_hd__nor2_1 _16340_ (.A(_07811_),
    .B(_07812_),
    .Y(_07813_));
 sky130_fd_sc_hd__xnor2_2 _16341_ (.A(_07794_),
    .B(_07813_),
    .Y(_07814_));
 sky130_fd_sc_hd__and2b_1 _16342_ (.A_N(_07776_),
    .B(_07814_),
    .X(_07815_));
 sky130_fd_sc_hd__xnor2_1 _16343_ (.A(_07776_),
    .B(_07814_),
    .Y(_07816_));
 sky130_fd_sc_hd__xor2_1 _16344_ (.A(_07775_),
    .B(_07816_),
    .X(_07817_));
 sky130_fd_sc_hd__xor2_1 _16345_ (.A(_07774_),
    .B(_07817_),
    .X(_07818_));
 sky130_fd_sc_hd__o21a_1 _16346_ (.A1(_07667_),
    .A2(_07714_),
    .B1(_07818_),
    .X(_07819_));
 sky130_fd_sc_hd__nor3_1 _16347_ (.A(_07667_),
    .B(_07714_),
    .C(_07818_),
    .Y(_07820_));
 sky130_fd_sc_hd__nor2_1 _16348_ (.A(_07709_),
    .B(_07712_),
    .Y(_07821_));
 sky130_fd_sc_hd__or3_1 _16349_ (.A(_07819_),
    .B(_07820_),
    .C(_07821_),
    .X(_07822_));
 sky130_fd_sc_hd__o21ai_1 _16350_ (.A1(_07819_),
    .A2(_07820_),
    .B1(_07821_),
    .Y(_07823_));
 sky130_fd_sc_hd__nand2_2 _16351_ (.A(_07822_),
    .B(_07823_),
    .Y(_07824_));
 sky130_fd_sc_hd__and2_1 _16352_ (.A(_07716_),
    .B(_07718_),
    .X(_07825_));
 sky130_fd_sc_hd__or2_1 _16353_ (.A(_07824_),
    .B(_07825_),
    .X(_07826_));
 sky130_fd_sc_hd__xnor2_2 _16354_ (.A(_07824_),
    .B(_07825_),
    .Y(_07827_));
 sky130_fd_sc_hd__a21oi_2 _16355_ (.A1(_07567_),
    .A2(_07684_),
    .B1(_07682_),
    .Y(_07828_));
 sky130_fd_sc_hd__xnor2_2 _16356_ (.A(_07827_),
    .B(_07828_),
    .Y(_07829_));
 sky130_fd_sc_hd__o21a_1 _16357_ (.A1(_07722_),
    .A2(_07723_),
    .B1(_07720_),
    .X(_07830_));
 sky130_fd_sc_hd__and2_1 _16358_ (.A(_07829_),
    .B(_07830_),
    .X(_07831_));
 sky130_fd_sc_hd__nor2_1 _16359_ (.A(_07829_),
    .B(_07830_),
    .Y(_07832_));
 sky130_fd_sc_hd__nor2_1 _16360_ (.A(_07831_),
    .B(_07832_),
    .Y(_07833_));
 sky130_fd_sc_hd__nor2_1 _16361_ (.A(_07726_),
    .B(_07729_),
    .Y(_07834_));
 sky130_fd_sc_hd__xnor2_2 _16362_ (.A(_07833_),
    .B(_07834_),
    .Y(_07835_));
 sky130_fd_sc_hd__and2_1 _16363_ (.A(net600),
    .B(\temp[30] ),
    .X(_07836_));
 sky130_fd_sc_hd__a221o_1 _16364_ (.A1(_02732_),
    .A2(net5),
    .B1(_07835_),
    .B2(_03058_),
    .C1(_07836_),
    .X(_07837_));
 sky130_fd_sc_hd__mux2_1 _16365_ (.A0(net738),
    .A1(_07837_),
    .S(net1),
    .X(_00297_));
 sky130_fd_sc_hd__and2b_1 _16366_ (.A_N(_07831_),
    .B(_07726_),
    .X(_07838_));
 sky130_fd_sc_hd__a211o_1 _16367_ (.A1(_07729_),
    .A2(_07833_),
    .B1(_07838_),
    .C1(_07832_),
    .X(_07839_));
 sky130_fd_sc_hd__and2b_1 _16368_ (.A_N(_07819_),
    .B(_07822_),
    .X(_07840_));
 sky130_fd_sc_hd__nand2_1 _16369_ (.A(net362),
    .B(net462),
    .Y(_07841_));
 sky130_fd_sc_hd__xor2_1 _16370_ (.A(_07840_),
    .B(_07841_),
    .X(_07842_));
 sky130_fd_sc_hd__nand2_1 _16371_ (.A(net368),
    .B(\mul0.a[29] ),
    .Y(_07843_));
 sky130_fd_sc_hd__xnor2_2 _16372_ (.A(_07737_),
    .B(_07843_),
    .Y(_07844_));
 sky130_fd_sc_hd__xnor2_2 _16373_ (.A(_07842_),
    .B(_07844_),
    .Y(_07845_));
 sky130_fd_sc_hd__or2_1 _16374_ (.A(net506),
    .B(net57),
    .X(_07846_));
 sky130_fd_sc_hd__a21oi_1 _16375_ (.A1(_07796_),
    .A2(_07804_),
    .B1(_07803_),
    .Y(_07847_));
 sky130_fd_sc_hd__xnor2_1 _16376_ (.A(_07846_),
    .B(_07847_),
    .Y(_07848_));
 sky130_fd_sc_hd__nand2_1 _16377_ (.A(net351),
    .B(net472),
    .Y(_07849_));
 sky130_fd_sc_hd__xnor2_1 _16378_ (.A(_07848_),
    .B(_07849_),
    .Y(_07850_));
 sky130_fd_sc_hd__xnor2_2 _16379_ (.A(_07845_),
    .B(_07850_),
    .Y(_07851_));
 sky130_fd_sc_hd__nand2_1 _16380_ (.A(net635),
    .B(net456),
    .Y(_07852_));
 sky130_fd_sc_hd__a21oi_1 _16381_ (.A1(_07774_),
    .A2(_07817_),
    .B1(_07772_),
    .Y(_07853_));
 sky130_fd_sc_hd__xnor2_1 _16382_ (.A(_07852_),
    .B(_07853_),
    .Y(_07854_));
 sky130_fd_sc_hd__mux2_1 _16383_ (.A0(_07760_),
    .A1(_07761_),
    .S(_07754_),
    .X(_07855_));
 sky130_fd_sc_hd__xnor2_2 _16384_ (.A(_07854_),
    .B(_07855_),
    .Y(_07856_));
 sky130_fd_sc_hd__o21a_1 _16385_ (.A1(_07827_),
    .A2(_07828_),
    .B1(_07826_),
    .X(_07857_));
 sky130_fd_sc_hd__a32o_1 _16386_ (.A1(net363),
    .A2(net465),
    .A3(_07743_),
    .B1(_07744_),
    .B2(net458),
    .X(_07858_));
 sky130_fd_sc_hd__xor2_1 _16387_ (.A(_07857_),
    .B(_07858_),
    .X(_07859_));
 sky130_fd_sc_hd__nand2_1 _16388_ (.A(_07807_),
    .B(_07809_),
    .Y(_07860_));
 sky130_fd_sc_hd__a21oi_1 _16389_ (.A1(_07677_),
    .A2(_07793_),
    .B1(_07791_),
    .Y(_07861_));
 sky130_fd_sc_hd__xnor2_1 _16390_ (.A(_07860_),
    .B(_07861_),
    .Y(_07862_));
 sky130_fd_sc_hd__nand2_1 _16391_ (.A(net359),
    .B(net465),
    .Y(_07863_));
 sky130_fd_sc_hd__xnor2_1 _16392_ (.A(_07862_),
    .B(_07863_),
    .Y(_07864_));
 sky130_fd_sc_hd__xnor2_1 _16393_ (.A(_07859_),
    .B(_07864_),
    .Y(_07865_));
 sky130_fd_sc_hd__xnor2_2 _16394_ (.A(_07856_),
    .B(_07865_),
    .Y(_07866_));
 sky130_fd_sc_hd__a31o_1 _16395_ (.A1(_07785_),
    .A2(_07786_),
    .A3(_07787_),
    .B1(_07784_),
    .X(_07867_));
 sky130_fd_sc_hd__nand2_1 _16396_ (.A(net476),
    .B(net347),
    .Y(_07868_));
 sky130_fd_sc_hd__o21ba_1 _16397_ (.A1(_07794_),
    .A2(_07812_),
    .B1_N(_07811_),
    .X(_07869_));
 sky130_fd_sc_hd__xnor2_1 _16398_ (.A(_07868_),
    .B(_07869_),
    .Y(_07870_));
 sky130_fd_sc_hd__nand2_1 _16399_ (.A(net489),
    .B(net336),
    .Y(_07871_));
 sky130_fd_sc_hd__xor2_1 _16400_ (.A(_07787_),
    .B(_07871_),
    .X(_07872_));
 sky130_fd_sc_hd__a32o_1 _16401_ (.A1(net351),
    .A2(net475),
    .A3(_07738_),
    .B1(_07739_),
    .B2(net468),
    .X(_07873_));
 sky130_fd_sc_hd__a31o_1 _16402_ (.A1(net502),
    .A2(net330),
    .A3(_07779_),
    .B1(_07778_),
    .X(_07874_));
 sky130_fd_sc_hd__xnor2_1 _16403_ (.A(_07873_),
    .B(_07874_),
    .Y(_07875_));
 sky130_fd_sc_hd__nand2_1 _16404_ (.A(net497),
    .B(net330),
    .Y(_07876_));
 sky130_fd_sc_hd__o31a_1 _16405_ (.A1(_07737_),
    .A2(_07765_),
    .A3(_07766_),
    .B1(_07769_),
    .X(_07877_));
 sky130_fd_sc_hd__nand2_1 _16406_ (.A(net502),
    .B(net328),
    .Y(_07878_));
 sky130_fd_sc_hd__xnor2_1 _16407_ (.A(_07877_),
    .B(_07878_),
    .Y(_07879_));
 sky130_fd_sc_hd__xnor2_1 _16408_ (.A(_07876_),
    .B(_07879_),
    .Y(_07880_));
 sky130_fd_sc_hd__nand2_1 _16409_ (.A(net493),
    .B(net333),
    .Y(_07881_));
 sky130_fd_sc_hd__xnor2_1 _16410_ (.A(_07880_),
    .B(_07881_),
    .Y(_07882_));
 sky130_fd_sc_hd__xnor2_1 _16411_ (.A(_07875_),
    .B(_07882_),
    .Y(_07883_));
 sky130_fd_sc_hd__xnor2_1 _16412_ (.A(_07872_),
    .B(_07883_),
    .Y(_07884_));
 sky130_fd_sc_hd__xnor2_1 _16413_ (.A(_07870_),
    .B(_07884_),
    .Y(_07885_));
 sky130_fd_sc_hd__nand2_1 _16414_ (.A(net354),
    .B(net468),
    .Y(_07886_));
 sky130_fd_sc_hd__a2bb2o_1 _16415_ (.A1_N(_07734_),
    .A2_N(_07770_),
    .B1(_06980_),
    .B2(_07624_),
    .X(_07887_));
 sky130_fd_sc_hd__xnor2_1 _16416_ (.A(_07886_),
    .B(_07887_),
    .Y(_07888_));
 sky130_fd_sc_hd__a31o_1 _16417_ (.A1(net488),
    .A2(\mul0.b[26] ),
    .A3(_07800_),
    .B1(_07799_),
    .X(_07889_));
 sky130_fd_sc_hd__nand2_1 _16418_ (.A(net479),
    .B(net343),
    .Y(_07890_));
 sky130_fd_sc_hd__o21a_1 _16419_ (.A1(_07742_),
    .A2(_07750_),
    .B1(_07749_),
    .X(_07891_));
 sky130_fd_sc_hd__xnor2_1 _16420_ (.A(_07890_),
    .B(_07891_),
    .Y(_07892_));
 sky130_fd_sc_hd__xnor2_1 _16421_ (.A(_07889_),
    .B(_07892_),
    .Y(_07893_));
 sky130_fd_sc_hd__xnor2_1 _16422_ (.A(_07888_),
    .B(_07893_),
    .Y(_07894_));
 sky130_fd_sc_hd__xnor2_1 _16423_ (.A(_07885_),
    .B(_07894_),
    .Y(_07895_));
 sky130_fd_sc_hd__nand2_1 _16424_ (.A(net485),
    .B(\mul0.b[26] ),
    .Y(_07896_));
 sky130_fd_sc_hd__a21o_1 _16425_ (.A1(_07775_),
    .A2(_07816_),
    .B1(_07815_),
    .X(_07897_));
 sky130_fd_sc_hd__a21oi_1 _16426_ (.A1(_07753_),
    .A2(_07763_),
    .B1(_07765_),
    .Y(_07898_));
 sky130_fd_sc_hd__o2111a_1 _16427_ (.A1(net455),
    .A2(_07755_),
    .B1(_07757_),
    .C1(net454),
    .D1(net374),
    .X(_07899_));
 sky130_fd_sc_hd__o211a_1 _16428_ (.A1(net385),
    .A2(net379),
    .B1(_02564_),
    .C1(net454),
    .X(_07900_));
 sky130_fd_sc_hd__nor2_1 _16429_ (.A(_07899_),
    .B(_07900_),
    .Y(_07901_));
 sky130_fd_sc_hd__xnor2_1 _16430_ (.A(_07898_),
    .B(_07901_),
    .Y(_07902_));
 sky130_fd_sc_hd__xnor2_1 _16431_ (.A(_07897_),
    .B(_07902_),
    .Y(_07903_));
 sky130_fd_sc_hd__xnor2_1 _16432_ (.A(_07896_),
    .B(_07903_),
    .Y(_07904_));
 sky130_fd_sc_hd__xnor2_1 _16433_ (.A(_07895_),
    .B(_07904_),
    .Y(_07905_));
 sky130_fd_sc_hd__xnor2_1 _16434_ (.A(_07867_),
    .B(_07905_),
    .Y(_07906_));
 sky130_fd_sc_hd__xnor2_2 _16435_ (.A(_07866_),
    .B(_07906_),
    .Y(_07907_));
 sky130_fd_sc_hd__xnor2_4 _16436_ (.A(_07851_),
    .B(_07907_),
    .Y(_07908_));
 sky130_fd_sc_hd__xnor2_2 _16437_ (.A(_07839_),
    .B(_07908_),
    .Y(_07909_));
 sky130_fd_sc_hd__a22o_1 _16438_ (.A1(net600),
    .A2(net833),
    .B1(_03058_),
    .B2(_07909_),
    .X(_07910_));
 sky130_fd_sc_hd__a21o_1 _16439_ (.A1(_02735_),
    .A2(net5),
    .B1(_07910_),
    .X(_07911_));
 sky130_fd_sc_hd__mux2_1 _16440_ (.A0(net878),
    .A1(_07911_),
    .S(net1),
    .X(_00298_));
 sky130_fd_sc_hd__and4_1 _16441_ (.A(net182),
    .B(net177),
    .C(net273),
    .D(net278),
    .X(_07912_));
 sky130_fd_sc_hd__a22oi_1 _16442_ (.A1(net182),
    .A2(net273),
    .B1(net278),
    .B2(net177),
    .Y(_07913_));
 sky130_fd_sc_hd__and4bb_1 _16443_ (.A_N(_07912_),
    .B_N(_07913_),
    .C(net172),
    .D(net283),
    .X(_07914_));
 sky130_fd_sc_hd__nor2_1 _16444_ (.A(_07912_),
    .B(_07914_),
    .Y(_07915_));
 sky130_fd_sc_hd__nand2_1 _16445_ (.A(net155),
    .B(net293),
    .Y(_07916_));
 sky130_fd_sc_hd__a22o_1 _16446_ (.A1(net165),
    .A2(net283),
    .B1(net288),
    .B2(net159),
    .X(_07917_));
 sky130_fd_sc_hd__and3_1 _16447_ (.A(net166),
    .B(net159),
    .C(net288),
    .X(_07918_));
 sky130_fd_sc_hd__a21bo_1 _16448_ (.A1(net283),
    .A2(_07918_),
    .B1_N(_07917_),
    .X(_07919_));
 sky130_fd_sc_hd__xor2_2 _16449_ (.A(_07916_),
    .B(_07919_),
    .X(_07920_));
 sky130_fd_sc_hd__nand2b_1 _16450_ (.A_N(_07915_),
    .B(_07920_),
    .Y(_07921_));
 sky130_fd_sc_hd__and4_1 _16451_ (.A(net165),
    .B(net159),
    .C(net288),
    .D(net294),
    .X(_07922_));
 sky130_fd_sc_hd__nand2_1 _16452_ (.A(net155),
    .B(net298),
    .Y(_07923_));
 sky130_fd_sc_hd__a22o_1 _16453_ (.A1(net165),
    .A2(net288),
    .B1(net294),
    .B2(net159),
    .X(_07924_));
 sky130_fd_sc_hd__and2b_1 _16454_ (.A_N(_07922_),
    .B(_07924_),
    .X(_07925_));
 sky130_fd_sc_hd__a31o_1 _16455_ (.A1(net155),
    .A2(net299),
    .A3(_07924_),
    .B1(_07922_),
    .X(_07926_));
 sky130_fd_sc_hd__xnor2_2 _16456_ (.A(_07915_),
    .B(_07920_),
    .Y(_07927_));
 sky130_fd_sc_hd__nand2_1 _16457_ (.A(_07926_),
    .B(_07927_),
    .Y(_07928_));
 sky130_fd_sc_hd__nand2_1 _16458_ (.A(net141),
    .B(net303),
    .Y(_07929_));
 sky130_fd_sc_hd__a22o_1 _16459_ (.A1(net150),
    .A2(net293),
    .B1(net298),
    .B2(net145),
    .X(_07930_));
 sky130_fd_sc_hd__and3_1 _16460_ (.A(net150),
    .B(net145),
    .C(net298),
    .X(_07931_));
 sky130_fd_sc_hd__a21bo_1 _16461_ (.A1(net294),
    .A2(_07931_),
    .B1_N(_07930_),
    .X(_07932_));
 sky130_fd_sc_hd__xor2_1 _16462_ (.A(_07929_),
    .B(_07932_),
    .X(_07933_));
 sky130_fd_sc_hd__and4_1 _16463_ (.A(net150),
    .B(net145),
    .C(net298),
    .D(net303),
    .X(_07934_));
 sky130_fd_sc_hd__nand2_1 _16464_ (.A(net141),
    .B(net308),
    .Y(_07935_));
 sky130_fd_sc_hd__a22o_1 _16465_ (.A1(net150),
    .A2(net298),
    .B1(net303),
    .B2(net145),
    .X(_07936_));
 sky130_fd_sc_hd__and2b_1 _16466_ (.A_N(_07934_),
    .B(_07936_),
    .X(_07937_));
 sky130_fd_sc_hd__a31o_1 _16467_ (.A1(net141),
    .A2(net308),
    .A3(_07936_),
    .B1(_07934_),
    .X(_07938_));
 sky130_fd_sc_hd__xor2_1 _16468_ (.A(_07933_),
    .B(_07938_),
    .X(_07939_));
 sky130_fd_sc_hd__a22o_1 _16469_ (.A1(net136),
    .A2(net308),
    .B1(net315),
    .B2(net131),
    .X(_07940_));
 sky130_fd_sc_hd__and4_1 _16470_ (.A(net136),
    .B(net131),
    .C(net308),
    .D(net315),
    .X(_07941_));
 sky130_fd_sc_hd__inv_2 _16471_ (.A(_07941_),
    .Y(_07942_));
 sky130_fd_sc_hd__and4_1 _16472_ (.A(net127),
    .B(net319),
    .C(_07940_),
    .D(_07942_),
    .X(_07943_));
 sky130_fd_sc_hd__a22oi_1 _16473_ (.A1(net127),
    .A2(net320),
    .B1(_07940_),
    .B2(_07942_),
    .Y(_07944_));
 sky130_fd_sc_hd__nor2_1 _16474_ (.A(_07943_),
    .B(_07944_),
    .Y(_07945_));
 sky130_fd_sc_hd__and2_1 _16475_ (.A(_07939_),
    .B(_07945_),
    .X(_07946_));
 sky130_fd_sc_hd__xnor2_1 _16476_ (.A(_07939_),
    .B(_07945_),
    .Y(_07947_));
 sky130_fd_sc_hd__a21o_1 _16477_ (.A1(_07921_),
    .A2(_07928_),
    .B1(_07947_),
    .X(_07948_));
 sky130_fd_sc_hd__xnor2_1 _16478_ (.A(_07935_),
    .B(_07937_),
    .Y(_07949_));
 sky130_fd_sc_hd__and4_1 _16479_ (.A(net150),
    .B(net145),
    .C(net303),
    .D(net309),
    .X(_07950_));
 sky130_fd_sc_hd__nand2_1 _16480_ (.A(net141),
    .B(net314),
    .Y(_07951_));
 sky130_fd_sc_hd__a22o_1 _16481_ (.A1(net150),
    .A2(net303),
    .B1(net309),
    .B2(net145),
    .X(_07952_));
 sky130_fd_sc_hd__and2b_1 _16482_ (.A_N(_07950_),
    .B(_07952_),
    .X(_07953_));
 sky130_fd_sc_hd__a31o_1 _16483_ (.A1(net141),
    .A2(net314),
    .A3(_07952_),
    .B1(_07950_),
    .X(_07954_));
 sky130_fd_sc_hd__and2_1 _16484_ (.A(_07949_),
    .B(_07954_),
    .X(_07955_));
 sky130_fd_sc_hd__xor2_1 _16485_ (.A(_07949_),
    .B(_07954_),
    .X(_07956_));
 sky130_fd_sc_hd__a22o_1 _16486_ (.A1(net136),
    .A2(net315),
    .B1(net319),
    .B2(net131),
    .X(_07957_));
 sky130_fd_sc_hd__and4_1 _16487_ (.A(net136),
    .B(net131),
    .C(net315),
    .D(net319),
    .X(_07958_));
 sky130_fd_sc_hd__inv_2 _16488_ (.A(_07958_),
    .Y(_07959_));
 sky130_fd_sc_hd__and4_1 _16489_ (.A(net127),
    .B(net323),
    .C(_07957_),
    .D(_07959_),
    .X(_07960_));
 sky130_fd_sc_hd__a22oi_1 _16490_ (.A1(net127),
    .A2(net323),
    .B1(_07957_),
    .B2(_07959_),
    .Y(_07961_));
 sky130_fd_sc_hd__nor2_1 _16491_ (.A(_07960_),
    .B(_07961_),
    .Y(_07962_));
 sky130_fd_sc_hd__and2_1 _16492_ (.A(_07956_),
    .B(_07962_),
    .X(_07963_));
 sky130_fd_sc_hd__nand3_2 _16493_ (.A(_07921_),
    .B(_07928_),
    .C(_07947_),
    .Y(_07964_));
 sky130_fd_sc_hd__o211ai_4 _16494_ (.A1(_07955_),
    .A2(_07963_),
    .B1(_07964_),
    .C1(_07948_),
    .Y(_07965_));
 sky130_fd_sc_hd__nor2_1 _16495_ (.A(_07958_),
    .B(_07960_),
    .Y(_07966_));
 sky130_fd_sc_hd__nand2_1 _16496_ (.A(net122),
    .B(net323),
    .Y(_07967_));
 sky130_fd_sc_hd__or2_1 _16497_ (.A(_07966_),
    .B(_07967_),
    .X(_07968_));
 sky130_fd_sc_hd__a22o_1 _16498_ (.A1(net319),
    .A2(net122),
    .B1(net117),
    .B2(net323),
    .X(_07969_));
 sky130_fd_sc_hd__and4_1 _16499_ (.A(net319),
    .B(net122),
    .C(net117),
    .D(net323),
    .X(_07970_));
 sky130_fd_sc_hd__nand4_1 _16500_ (.A(net320),
    .B(net122),
    .C(net117),
    .D(net323),
    .Y(_07971_));
 sky130_fd_sc_hd__o211a_2 _16501_ (.A1(_07941_),
    .A2(_07943_),
    .B1(_07969_),
    .C1(_07971_),
    .X(_07972_));
 sky130_fd_sc_hd__a211oi_1 _16502_ (.A1(_07969_),
    .A2(_07971_),
    .B1(_07941_),
    .C1(_07943_),
    .Y(_07973_));
 sky130_fd_sc_hd__or3_2 _16503_ (.A(_07968_),
    .B(_07972_),
    .C(_07973_),
    .X(_07974_));
 sky130_fd_sc_hd__o21ai_1 _16504_ (.A1(_07972_),
    .A2(_07973_),
    .B1(_07968_),
    .Y(_07975_));
 sky130_fd_sc_hd__nand2_1 _16505_ (.A(_07974_),
    .B(_07975_),
    .Y(_07976_));
 sky130_fd_sc_hd__a21oi_2 _16506_ (.A1(_07948_),
    .A2(_07965_),
    .B1(_07976_),
    .Y(_07977_));
 sky130_fd_sc_hd__and4_1 _16507_ (.A(net181),
    .B(net177),
    .C(net268),
    .D(net273),
    .X(_07978_));
 sky130_fd_sc_hd__a22oi_1 _16508_ (.A1(net181),
    .A2(net268),
    .B1(net273),
    .B2(net176),
    .Y(_07979_));
 sky130_fd_sc_hd__and4bb_1 _16509_ (.A_N(_07978_),
    .B_N(_07979_),
    .C(net171),
    .D(net278),
    .X(_07980_));
 sky130_fd_sc_hd__a22o_1 _16510_ (.A1(net165),
    .A2(net278),
    .B1(net283),
    .B2(net160),
    .X(_07981_));
 sky130_fd_sc_hd__nand4_2 _16511_ (.A(net165),
    .B(net159),
    .C(net278),
    .D(net283),
    .Y(_07982_));
 sky130_fd_sc_hd__nand4_1 _16512_ (.A(net155),
    .B(net289),
    .C(_07981_),
    .D(_07982_),
    .Y(_07983_));
 sky130_fd_sc_hd__a22o_1 _16513_ (.A1(net155),
    .A2(net289),
    .B1(_07981_),
    .B2(_07982_),
    .X(_07984_));
 sky130_fd_sc_hd__o211a_1 _16514_ (.A1(_07978_),
    .A2(_07980_),
    .B1(_07983_),
    .C1(_07984_),
    .X(_07985_));
 sky130_fd_sc_hd__a32o_1 _16515_ (.A1(net155),
    .A2(net293),
    .A3(_07917_),
    .B1(_07918_),
    .B2(net283),
    .X(_07986_));
 sky130_fd_sc_hd__a211o_1 _16516_ (.A1(_07983_),
    .A2(_07984_),
    .B1(_07978_),
    .C1(_07980_),
    .X(_07987_));
 sky130_fd_sc_hd__nand2b_1 _16517_ (.A_N(_07985_),
    .B(_07987_),
    .Y(_07988_));
 sky130_fd_sc_hd__a21o_1 _16518_ (.A1(_07986_),
    .A2(_07987_),
    .B1(_07985_),
    .X(_07989_));
 sky130_fd_sc_hd__and2_1 _16519_ (.A(net141),
    .B(net300),
    .X(_07990_));
 sky130_fd_sc_hd__a22o_1 _16520_ (.A1(net289),
    .A2(net150),
    .B1(net145),
    .B2(net293),
    .X(_07991_));
 sky130_fd_sc_hd__nand4_1 _16521_ (.A(net289),
    .B(net150),
    .C(net145),
    .D(net295),
    .Y(_07992_));
 sky130_fd_sc_hd__nand3_1 _16522_ (.A(_07990_),
    .B(_07991_),
    .C(_07992_),
    .Y(_07993_));
 sky130_fd_sc_hd__a21o_1 _16523_ (.A1(_07991_),
    .A2(_07992_),
    .B1(_07990_),
    .X(_07994_));
 sky130_fd_sc_hd__a32o_1 _16524_ (.A1(net141),
    .A2(net305),
    .A3(_07930_),
    .B1(_07931_),
    .B2(net294),
    .X(_07995_));
 sky130_fd_sc_hd__nand3_2 _16525_ (.A(_07993_),
    .B(_07994_),
    .C(_07995_),
    .Y(_07996_));
 sky130_fd_sc_hd__a21o_1 _16526_ (.A1(_07993_),
    .A2(_07994_),
    .B1(_07995_),
    .X(_07997_));
 sky130_fd_sc_hd__nand2_1 _16527_ (.A(net127),
    .B(net315),
    .Y(_07998_));
 sky130_fd_sc_hd__a22oi_1 _16528_ (.A1(net136),
    .A2(net305),
    .B1(net310),
    .B2(net131),
    .Y(_07999_));
 sky130_fd_sc_hd__and4_1 _16529_ (.A(net136),
    .B(net131),
    .C(net305),
    .D(net310),
    .X(_08000_));
 sky130_fd_sc_hd__nor2_1 _16530_ (.A(_07999_),
    .B(_08000_),
    .Y(_08001_));
 sky130_fd_sc_hd__xnor2_1 _16531_ (.A(_07998_),
    .B(_08001_),
    .Y(_08002_));
 sky130_fd_sc_hd__nand3_2 _16532_ (.A(_07996_),
    .B(_07997_),
    .C(_08002_),
    .Y(_08003_));
 sky130_fd_sc_hd__a21o_1 _16533_ (.A1(_07996_),
    .A2(_07997_),
    .B1(_08002_),
    .X(_08004_));
 sky130_fd_sc_hd__nand3_1 _16534_ (.A(_07989_),
    .B(_08003_),
    .C(_08004_),
    .Y(_08005_));
 sky130_fd_sc_hd__a21oi_1 _16535_ (.A1(_07933_),
    .A2(_07938_),
    .B1(_07946_),
    .Y(_08006_));
 sky130_fd_sc_hd__a21o_1 _16536_ (.A1(_08003_),
    .A2(_08004_),
    .B1(_07989_),
    .X(_08007_));
 sky130_fd_sc_hd__nand2_1 _16537_ (.A(_08005_),
    .B(_08007_),
    .Y(_08008_));
 sky130_fd_sc_hd__o21ai_1 _16538_ (.A1(_08006_),
    .A2(_08008_),
    .B1(_08005_),
    .Y(_08009_));
 sky130_fd_sc_hd__a31o_1 _16539_ (.A1(net127),
    .A2(net315),
    .A3(_08001_),
    .B1(_08000_),
    .X(_08010_));
 sky130_fd_sc_hd__nand2_1 _16540_ (.A(net114),
    .B(net323),
    .Y(_08011_));
 sky130_fd_sc_hd__and4_1 _16541_ (.A(net315),
    .B(net319),
    .C(net122),
    .D(net117),
    .X(_08012_));
 sky130_fd_sc_hd__a22o_1 _16542_ (.A1(net315),
    .A2(net122),
    .B1(net117),
    .B2(net319),
    .X(_08013_));
 sky130_fd_sc_hd__and2b_1 _16543_ (.A_N(_08012_),
    .B(_08013_),
    .X(_08014_));
 sky130_fd_sc_hd__xnor2_1 _16544_ (.A(_08011_),
    .B(_08014_),
    .Y(_08015_));
 sky130_fd_sc_hd__or2_1 _16545_ (.A(_08010_),
    .B(_08015_),
    .X(_08016_));
 sky130_fd_sc_hd__inv_2 _16546_ (.A(_08016_),
    .Y(_08017_));
 sky130_fd_sc_hd__and2_1 _16547_ (.A(_08010_),
    .B(_08015_),
    .X(_08018_));
 sky130_fd_sc_hd__nor2_2 _16548_ (.A(_08017_),
    .B(_08018_),
    .Y(_08019_));
 sky130_fd_sc_hd__nor2_1 _16549_ (.A(_07970_),
    .B(_07972_),
    .Y(_08020_));
 sky130_fd_sc_hd__xnor2_1 _16550_ (.A(_08019_),
    .B(_08020_),
    .Y(_08021_));
 sky130_fd_sc_hd__nand2_1 _16551_ (.A(_08009_),
    .B(_08021_),
    .Y(_08022_));
 sky130_fd_sc_hd__xnor2_1 _16552_ (.A(_08009_),
    .B(_08021_),
    .Y(_08023_));
 sky130_fd_sc_hd__xor2_1 _16553_ (.A(_07974_),
    .B(_08023_),
    .X(_08024_));
 sky130_fd_sc_hd__and4_1 _16554_ (.A(\mul1.b[3] ),
    .B(net177),
    .C(net263),
    .D(net268),
    .X(_08025_));
 sky130_fd_sc_hd__nand2_1 _16555_ (.A(net172),
    .B(net273),
    .Y(_08026_));
 sky130_fd_sc_hd__a22o_1 _16556_ (.A1(\mul1.b[3] ),
    .A2(net263),
    .B1(net268),
    .B2(net177),
    .X(_08027_));
 sky130_fd_sc_hd__and2b_1 _16557_ (.A_N(_08025_),
    .B(_08027_),
    .X(_08028_));
 sky130_fd_sc_hd__a31o_1 _16558_ (.A1(net172),
    .A2(net273),
    .A3(_08027_),
    .B1(_08025_),
    .X(_08029_));
 sky130_fd_sc_hd__a22o_1 _16559_ (.A1(net166),
    .A2(net273),
    .B1(net278),
    .B2(net160),
    .X(_08030_));
 sky130_fd_sc_hd__nand4_2 _16560_ (.A(net166),
    .B(net160),
    .C(net273),
    .D(net278),
    .Y(_08031_));
 sky130_fd_sc_hd__nand4_2 _16561_ (.A(\mul1.b[8] ),
    .B(net284),
    .C(_08030_),
    .D(_08031_),
    .Y(_08032_));
 sky130_fd_sc_hd__a22o_1 _16562_ (.A1(net155),
    .A2(net284),
    .B1(_08030_),
    .B2(_08031_),
    .X(_08033_));
 sky130_fd_sc_hd__nand3_1 _16563_ (.A(_08029_),
    .B(_08032_),
    .C(_08033_),
    .Y(_08034_));
 sky130_fd_sc_hd__nand2_1 _16564_ (.A(_07982_),
    .B(_07983_),
    .Y(_08035_));
 sky130_fd_sc_hd__a21o_1 _16565_ (.A1(_08032_),
    .A2(_08033_),
    .B1(_08029_),
    .X(_08036_));
 sky130_fd_sc_hd__and3_1 _16566_ (.A(_08034_),
    .B(_08035_),
    .C(_08036_),
    .X(_08037_));
 sky130_fd_sc_hd__a21bo_1 _16567_ (.A1(_08035_),
    .A2(_08036_),
    .B1_N(_08034_),
    .X(_08038_));
 sky130_fd_sc_hd__nand2_1 _16568_ (.A(net127),
    .B(net310),
    .Y(_08039_));
 sky130_fd_sc_hd__and4_1 _16569_ (.A(net300),
    .B(net136),
    .C(net131),
    .D(net305),
    .X(_08040_));
 sky130_fd_sc_hd__a22o_1 _16570_ (.A1(net300),
    .A2(net136),
    .B1(net131),
    .B2(net305),
    .X(_08041_));
 sky130_fd_sc_hd__and2b_1 _16571_ (.A_N(_08040_),
    .B(_08041_),
    .X(_08042_));
 sky130_fd_sc_hd__xnor2_1 _16572_ (.A(_08039_),
    .B(_08042_),
    .Y(_08043_));
 sky130_fd_sc_hd__nand4_1 _16573_ (.A(net284),
    .B(net292),
    .C(net150),
    .D(net145),
    .Y(_08044_));
 sky130_fd_sc_hd__a22o_1 _16574_ (.A1(net284),
    .A2(net151),
    .B1(net145),
    .B2(net292),
    .X(_08045_));
 sky130_fd_sc_hd__nand4_1 _16575_ (.A(net141),
    .B(net295),
    .C(_08044_),
    .D(_08045_),
    .Y(_08046_));
 sky130_fd_sc_hd__a22o_1 _16576_ (.A1(net141),
    .A2(net295),
    .B1(_08044_),
    .B2(_08045_),
    .X(_08047_));
 sky130_fd_sc_hd__a21bo_1 _16577_ (.A1(_07990_),
    .A2(_07991_),
    .B1_N(_07992_),
    .X(_08048_));
 sky130_fd_sc_hd__nand3_1 _16578_ (.A(_08046_),
    .B(_08047_),
    .C(_08048_),
    .Y(_08049_));
 sky130_fd_sc_hd__a21o_1 _16579_ (.A1(_08046_),
    .A2(_08047_),
    .B1(_08048_),
    .X(_08050_));
 sky130_fd_sc_hd__nand3_1 _16580_ (.A(_08043_),
    .B(_08049_),
    .C(_08050_),
    .Y(_08051_));
 sky130_fd_sc_hd__a21o_1 _16581_ (.A1(_08049_),
    .A2(_08050_),
    .B1(_08043_),
    .X(_08052_));
 sky130_fd_sc_hd__and3_1 _16582_ (.A(_08038_),
    .B(_08051_),
    .C(_08052_),
    .X(_08053_));
 sky130_fd_sc_hd__a21oi_2 _16583_ (.A1(_08051_),
    .A2(_08052_),
    .B1(_08038_),
    .Y(_08054_));
 sky130_fd_sc_hd__a211oi_4 _16584_ (.A1(_07996_),
    .A2(_08003_),
    .B1(_08053_),
    .C1(_08054_),
    .Y(_08055_));
 sky130_fd_sc_hd__o211a_1 _16585_ (.A1(_08053_),
    .A2(_08054_),
    .B1(_07996_),
    .C1(_08003_),
    .X(_08056_));
 sky130_fd_sc_hd__nand2_2 _16586_ (.A(_08031_),
    .B(_08032_),
    .Y(_08057_));
 sky130_fd_sc_hd__and4_1 _16587_ (.A(\mul1.b[3] ),
    .B(net177),
    .C(net258),
    .D(net263),
    .X(_08058_));
 sky130_fd_sc_hd__a22oi_1 _16588_ (.A1(\mul1.b[3] ),
    .A2(net258),
    .B1(net263),
    .B2(net177),
    .Y(_08059_));
 sky130_fd_sc_hd__and4bb_1 _16589_ (.A_N(_08058_),
    .B_N(_08059_),
    .C(net172),
    .D(net268),
    .X(_08060_));
 sky130_fd_sc_hd__nor2_1 _16590_ (.A(_08058_),
    .B(_08060_),
    .Y(_08061_));
 sky130_fd_sc_hd__nand2_1 _16591_ (.A(net155),
    .B(net279),
    .Y(_08062_));
 sky130_fd_sc_hd__and4_1 _16592_ (.A(net268),
    .B(net166),
    .C(net160),
    .D(net274),
    .X(_08063_));
 sky130_fd_sc_hd__a22o_1 _16593_ (.A1(net268),
    .A2(net166),
    .B1(net160),
    .B2(net274),
    .X(_08064_));
 sky130_fd_sc_hd__and2b_1 _16594_ (.A_N(_08063_),
    .B(_08064_),
    .X(_08065_));
 sky130_fd_sc_hd__xnor2_2 _16595_ (.A(_08062_),
    .B(_08065_),
    .Y(_08066_));
 sky130_fd_sc_hd__nand2b_1 _16596_ (.A_N(_08061_),
    .B(_08066_),
    .Y(_08067_));
 sky130_fd_sc_hd__xnor2_2 _16597_ (.A(_08061_),
    .B(_08066_),
    .Y(_08068_));
 sky130_fd_sc_hd__nand2_1 _16598_ (.A(_08057_),
    .B(_08068_),
    .Y(_08069_));
 sky130_fd_sc_hd__xor2_2 _16599_ (.A(_08057_),
    .B(_08068_),
    .X(_08070_));
 sky130_fd_sc_hd__nand2_1 _16600_ (.A(net175),
    .B(net263),
    .Y(_08071_));
 sky130_fd_sc_hd__a22oi_2 _16601_ (.A1(net257),
    .A2(net185),
    .B1(net180),
    .B2(net258),
    .Y(_08072_));
 sky130_fd_sc_hd__and4_1 _16602_ (.A(net257),
    .B(net185),
    .C(net180),
    .D(net258),
    .X(_08073_));
 sky130_fd_sc_hd__nor2_1 _16603_ (.A(_08072_),
    .B(_08073_),
    .Y(_08074_));
 sky130_fd_sc_hd__xnor2_2 _16604_ (.A(_08071_),
    .B(_08074_),
    .Y(_08075_));
 sky130_fd_sc_hd__and2_1 _16605_ (.A(net187),
    .B(net252),
    .X(_08076_));
 sky130_fd_sc_hd__nand4_1 _16606_ (.A(net625),
    .B(net247),
    .C(net192),
    .D(net630),
    .Y(_08077_));
 sky130_fd_sc_hd__a22o_1 _16607_ (.A1(net625),
    .A2(net247),
    .B1(net192),
    .B2(net630),
    .X(_08078_));
 sky130_fd_sc_hd__nand3_1 _16608_ (.A(_08076_),
    .B(_08077_),
    .C(_08078_),
    .Y(_08079_));
 sky130_fd_sc_hd__a21o_1 _16609_ (.A1(_08077_),
    .A2(_08078_),
    .B1(_08076_),
    .X(_08080_));
 sky130_fd_sc_hd__nand4_2 _16610_ (.A(\mul1.b[0] ),
    .B(\mul1.b[1] ),
    .C(net630),
    .D(net252),
    .Y(_08081_));
 sky130_fd_sc_hd__and2_1 _16611_ (.A(\mul1.b[2] ),
    .B(net257),
    .X(_08082_));
 sky130_fd_sc_hd__a22o_1 _16612_ (.A1(\mul1.b[0] ),
    .A2(net630),
    .B1(net252),
    .B2(\mul1.b[1] ),
    .X(_08083_));
 sky130_fd_sc_hd__nand3_1 _16613_ (.A(_08081_),
    .B(_08082_),
    .C(_08083_),
    .Y(_08084_));
 sky130_fd_sc_hd__a21bo_1 _16614_ (.A1(_08082_),
    .A2(_08083_),
    .B1_N(_08081_),
    .X(_08085_));
 sky130_fd_sc_hd__nand3_2 _16615_ (.A(_08079_),
    .B(_08080_),
    .C(_08085_),
    .Y(_08086_));
 sky130_fd_sc_hd__a21o_1 _16616_ (.A1(_08079_),
    .A2(_08080_),
    .B1(_08085_),
    .X(_08087_));
 sky130_fd_sc_hd__nand3_2 _16617_ (.A(_08075_),
    .B(_08086_),
    .C(_08087_),
    .Y(_08088_));
 sky130_fd_sc_hd__a21o_1 _16618_ (.A1(_08086_),
    .A2(_08087_),
    .B1(_08075_),
    .X(_08089_));
 sky130_fd_sc_hd__nand4_2 _16619_ (.A(net622),
    .B(net189),
    .C(net252),
    .D(net257),
    .Y(_08090_));
 sky130_fd_sc_hd__and2_1 _16620_ (.A(net186),
    .B(net258),
    .X(_08091_));
 sky130_fd_sc_hd__a22o_1 _16621_ (.A1(net622),
    .A2(net252),
    .B1(net257),
    .B2(net189),
    .X(_08092_));
 sky130_fd_sc_hd__nand3_1 _16622_ (.A(_08090_),
    .B(_08091_),
    .C(_08092_),
    .Y(_08093_));
 sky130_fd_sc_hd__a21bo_1 _16623_ (.A1(_08091_),
    .A2(_08092_),
    .B1_N(_08090_),
    .X(_08094_));
 sky130_fd_sc_hd__a21o_1 _16624_ (.A1(_08081_),
    .A2(_08083_),
    .B1(_08082_),
    .X(_08095_));
 sky130_fd_sc_hd__nand3_1 _16625_ (.A(_08084_),
    .B(_08094_),
    .C(_08095_),
    .Y(_08096_));
 sky130_fd_sc_hd__a21o_1 _16626_ (.A1(_08084_),
    .A2(_08095_),
    .B1(_08094_),
    .X(_08097_));
 sky130_fd_sc_hd__o2bb2a_1 _16627_ (.A1_N(net172),
    .A2_N(net268),
    .B1(_08058_),
    .B2(_08059_),
    .X(_08098_));
 sky130_fd_sc_hd__nor2_1 _16628_ (.A(_08060_),
    .B(_08098_),
    .Y(_08099_));
 sky130_fd_sc_hd__nand3_2 _16629_ (.A(_08096_),
    .B(_08097_),
    .C(_08099_),
    .Y(_08100_));
 sky130_fd_sc_hd__a21bo_1 _16630_ (.A1(_08097_),
    .A2(_08099_),
    .B1_N(_08096_),
    .X(_08101_));
 sky130_fd_sc_hd__nand3_4 _16631_ (.A(_08088_),
    .B(_08089_),
    .C(_08101_),
    .Y(_08102_));
 sky130_fd_sc_hd__a21o_1 _16632_ (.A1(_08088_),
    .A2(_08089_),
    .B1(_08101_),
    .X(_08103_));
 sky130_fd_sc_hd__and3_1 _16633_ (.A(_08070_),
    .B(_08102_),
    .C(_08103_),
    .X(_08104_));
 sky130_fd_sc_hd__nand3_2 _16634_ (.A(_08070_),
    .B(_08102_),
    .C(_08103_),
    .Y(_08105_));
 sky130_fd_sc_hd__a21oi_2 _16635_ (.A1(_08102_),
    .A2(_08103_),
    .B1(_08070_),
    .Y(_08106_));
 sky130_fd_sc_hd__nand4_1 _16636_ (.A(net622),
    .B(net189),
    .C(net257),
    .D(net258),
    .Y(_08107_));
 sky130_fd_sc_hd__and2_1 _16637_ (.A(net186),
    .B(net263),
    .X(_08108_));
 sky130_fd_sc_hd__a22o_1 _16638_ (.A1(net622),
    .A2(net257),
    .B1(net258),
    .B2(net189),
    .X(_08109_));
 sky130_fd_sc_hd__nand3_1 _16639_ (.A(_08107_),
    .B(_08108_),
    .C(_08109_),
    .Y(_08110_));
 sky130_fd_sc_hd__a21bo_1 _16640_ (.A1(_08108_),
    .A2(_08109_),
    .B1_N(_08107_),
    .X(_08111_));
 sky130_fd_sc_hd__a21o_1 _16641_ (.A1(_08090_),
    .A2(_08092_),
    .B1(_08091_),
    .X(_08112_));
 sky130_fd_sc_hd__nand3_1 _16642_ (.A(_08093_),
    .B(_08111_),
    .C(_08112_),
    .Y(_08113_));
 sky130_fd_sc_hd__a21o_1 _16643_ (.A1(_08093_),
    .A2(_08112_),
    .B1(_08111_),
    .X(_08114_));
 sky130_fd_sc_hd__xnor2_2 _16644_ (.A(_08026_),
    .B(_08028_),
    .Y(_08115_));
 sky130_fd_sc_hd__nand3_2 _16645_ (.A(_08113_),
    .B(_08114_),
    .C(_08115_),
    .Y(_08116_));
 sky130_fd_sc_hd__a21bo_1 _16646_ (.A1(_08114_),
    .A2(_08115_),
    .B1_N(_08113_),
    .X(_08117_));
 sky130_fd_sc_hd__a21o_1 _16647_ (.A1(_08096_),
    .A2(_08097_),
    .B1(_08099_),
    .X(_08118_));
 sky130_fd_sc_hd__nand3_4 _16648_ (.A(_08100_),
    .B(_08117_),
    .C(_08118_),
    .Y(_08119_));
 sky130_fd_sc_hd__a21o_1 _16649_ (.A1(_08100_),
    .A2(_08118_),
    .B1(_08117_),
    .X(_08120_));
 sky130_fd_sc_hd__a21oi_1 _16650_ (.A1(_08034_),
    .A2(_08036_),
    .B1(_08035_),
    .Y(_08121_));
 sky130_fd_sc_hd__nor2_1 _16651_ (.A(_08037_),
    .B(_08121_),
    .Y(_08122_));
 sky130_fd_sc_hd__and3_1 _16652_ (.A(_08119_),
    .B(_08120_),
    .C(_08122_),
    .X(_08123_));
 sky130_fd_sc_hd__nand3_2 _16653_ (.A(_08119_),
    .B(_08120_),
    .C(_08122_),
    .Y(_08124_));
 sky130_fd_sc_hd__a211oi_4 _16654_ (.A1(_08119_),
    .A2(_08124_),
    .B1(_08104_),
    .C1(_08106_),
    .Y(_08125_));
 sky130_fd_sc_hd__o211a_1 _16655_ (.A1(_08104_),
    .A2(_08106_),
    .B1(_08119_),
    .C1(_08124_),
    .X(_08126_));
 sky130_fd_sc_hd__nor4_2 _16656_ (.A(_08055_),
    .B(_08056_),
    .C(_08125_),
    .D(_08126_),
    .Y(_08127_));
 sky130_fd_sc_hd__or4_1 _16657_ (.A(_08055_),
    .B(_08056_),
    .C(_08125_),
    .D(_08126_),
    .X(_08128_));
 sky130_fd_sc_hd__o22ai_2 _16658_ (.A1(_08055_),
    .A2(_08056_),
    .B1(_08125_),
    .B2(_08126_),
    .Y(_08129_));
 sky130_fd_sc_hd__nand4_1 _16659_ (.A(net621),
    .B(net188),
    .C(net258),
    .D(net263),
    .Y(_08130_));
 sky130_fd_sc_hd__and2_1 _16660_ (.A(net186),
    .B(net268),
    .X(_08131_));
 sky130_fd_sc_hd__a22o_1 _16661_ (.A1(net621),
    .A2(net258),
    .B1(net263),
    .B2(net188),
    .X(_08132_));
 sky130_fd_sc_hd__nand3_1 _16662_ (.A(_08130_),
    .B(_08131_),
    .C(_08132_),
    .Y(_08133_));
 sky130_fd_sc_hd__a21bo_1 _16663_ (.A1(_08131_),
    .A2(_08132_),
    .B1_N(_08130_),
    .X(_08134_));
 sky130_fd_sc_hd__a21o_1 _16664_ (.A1(_08107_),
    .A2(_08109_),
    .B1(_08108_),
    .X(_08135_));
 sky130_fd_sc_hd__nand3_1 _16665_ (.A(_08110_),
    .B(_08134_),
    .C(_08135_),
    .Y(_08136_));
 sky130_fd_sc_hd__a21o_1 _16666_ (.A1(_08110_),
    .A2(_08135_),
    .B1(_08134_),
    .X(_08137_));
 sky130_fd_sc_hd__o2bb2a_1 _16667_ (.A1_N(net171),
    .A2_N(net278),
    .B1(_07978_),
    .B2(_07979_),
    .X(_08138_));
 sky130_fd_sc_hd__nor2_1 _16668_ (.A(_07980_),
    .B(_08138_),
    .Y(_08139_));
 sky130_fd_sc_hd__nand3_1 _16669_ (.A(_08136_),
    .B(_08137_),
    .C(_08139_),
    .Y(_08140_));
 sky130_fd_sc_hd__a21bo_1 _16670_ (.A1(_08137_),
    .A2(_08139_),
    .B1_N(_08136_),
    .X(_08141_));
 sky130_fd_sc_hd__a21o_1 _16671_ (.A1(_08113_),
    .A2(_08114_),
    .B1(_08115_),
    .X(_08142_));
 sky130_fd_sc_hd__nand3_4 _16672_ (.A(_08116_),
    .B(_08141_),
    .C(_08142_),
    .Y(_08143_));
 sky130_fd_sc_hd__a21o_1 _16673_ (.A1(_08116_),
    .A2(_08142_),
    .B1(_08141_),
    .X(_08144_));
 sky130_fd_sc_hd__xnor2_1 _16674_ (.A(_07986_),
    .B(_07988_),
    .Y(_08145_));
 sky130_fd_sc_hd__and3_1 _16675_ (.A(_08143_),
    .B(_08144_),
    .C(_08145_),
    .X(_08146_));
 sky130_fd_sc_hd__nand3_2 _16676_ (.A(_08143_),
    .B(_08144_),
    .C(_08145_),
    .Y(_08147_));
 sky130_fd_sc_hd__a21oi_2 _16677_ (.A1(_08119_),
    .A2(_08120_),
    .B1(_08122_),
    .Y(_08148_));
 sky130_fd_sc_hd__a211oi_4 _16678_ (.A1(_08143_),
    .A2(_08147_),
    .B1(_08148_),
    .C1(_08123_),
    .Y(_08149_));
 sky130_fd_sc_hd__o211a_1 _16679_ (.A1(_08123_),
    .A2(_08148_),
    .B1(_08147_),
    .C1(_08143_),
    .X(_08150_));
 sky130_fd_sc_hd__xnor2_1 _16680_ (.A(_08006_),
    .B(_08008_),
    .Y(_08151_));
 sky130_fd_sc_hd__nor3_1 _16681_ (.A(_08149_),
    .B(_08150_),
    .C(_08151_),
    .Y(_08152_));
 sky130_fd_sc_hd__or3_2 _16682_ (.A(_08149_),
    .B(_08150_),
    .C(_08151_),
    .X(_08153_));
 sky130_fd_sc_hd__o211ai_2 _16683_ (.A1(_08149_),
    .A2(_08152_),
    .B1(_08128_),
    .C1(_08129_),
    .Y(_08154_));
 sky130_fd_sc_hd__inv_2 _16684_ (.A(_08154_),
    .Y(_08155_));
 sky130_fd_sc_hd__a211o_1 _16685_ (.A1(_08128_),
    .A2(_08129_),
    .B1(_08149_),
    .C1(_08152_),
    .X(_08156_));
 sky130_fd_sc_hd__and3_2 _16686_ (.A(_08024_),
    .B(_08154_),
    .C(_08156_),
    .X(_08157_));
 sky130_fd_sc_hd__a21oi_1 _16687_ (.A1(_08154_),
    .A2(_08156_),
    .B1(_08024_),
    .Y(_08158_));
 sky130_fd_sc_hd__nand4_2 _16688_ (.A(net621),
    .B(net188),
    .C(net263),
    .D(net268),
    .Y(_08159_));
 sky130_fd_sc_hd__and2_1 _16689_ (.A(net186),
    .B(net273),
    .X(_08160_));
 sky130_fd_sc_hd__a22o_1 _16690_ (.A1(net621),
    .A2(net263),
    .B1(net268),
    .B2(net188),
    .X(_08161_));
 sky130_fd_sc_hd__nand3_1 _16691_ (.A(_08159_),
    .B(_08160_),
    .C(_08161_),
    .Y(_08162_));
 sky130_fd_sc_hd__a21bo_1 _16692_ (.A1(_08160_),
    .A2(_08161_),
    .B1_N(_08159_),
    .X(_08163_));
 sky130_fd_sc_hd__a21o_1 _16693_ (.A1(_08130_),
    .A2(_08132_),
    .B1(_08131_),
    .X(_08164_));
 sky130_fd_sc_hd__nand3_1 _16694_ (.A(_08133_),
    .B(_08163_),
    .C(_08164_),
    .Y(_08165_));
 sky130_fd_sc_hd__a21o_1 _16695_ (.A1(_08133_),
    .A2(_08164_),
    .B1(_08163_),
    .X(_08166_));
 sky130_fd_sc_hd__o2bb2a_1 _16696_ (.A1_N(net171),
    .A2_N(net283),
    .B1(_07912_),
    .B2(_07913_),
    .X(_08167_));
 sky130_fd_sc_hd__nor2_1 _16697_ (.A(_07914_),
    .B(_08167_),
    .Y(_08168_));
 sky130_fd_sc_hd__nand3_2 _16698_ (.A(_08165_),
    .B(_08166_),
    .C(_08168_),
    .Y(_08169_));
 sky130_fd_sc_hd__a21bo_1 _16699_ (.A1(_08166_),
    .A2(_08168_),
    .B1_N(_08165_),
    .X(_08170_));
 sky130_fd_sc_hd__a21o_1 _16700_ (.A1(_08136_),
    .A2(_08137_),
    .B1(_08139_),
    .X(_08171_));
 sky130_fd_sc_hd__nand3_2 _16701_ (.A(_08140_),
    .B(_08170_),
    .C(_08171_),
    .Y(_08172_));
 sky130_fd_sc_hd__a21o_1 _16702_ (.A1(_08140_),
    .A2(_08171_),
    .B1(_08170_),
    .X(_08173_));
 sky130_fd_sc_hd__xor2_2 _16703_ (.A(_07926_),
    .B(_07927_),
    .X(_08174_));
 sky130_fd_sc_hd__and3_1 _16704_ (.A(_08172_),
    .B(_08173_),
    .C(_08174_),
    .X(_08175_));
 sky130_fd_sc_hd__nand3_1 _16705_ (.A(_08172_),
    .B(_08173_),
    .C(_08174_),
    .Y(_08176_));
 sky130_fd_sc_hd__a21oi_1 _16706_ (.A1(_08143_),
    .A2(_08144_),
    .B1(_08145_),
    .Y(_08177_));
 sky130_fd_sc_hd__a211o_2 _16707_ (.A1(_08172_),
    .A2(_08176_),
    .B1(_08177_),
    .C1(_08146_),
    .X(_08178_));
 sky130_fd_sc_hd__inv_2 _16708_ (.A(_08178_),
    .Y(_08179_));
 sky130_fd_sc_hd__o211ai_2 _16709_ (.A1(_08146_),
    .A2(_08177_),
    .B1(_08176_),
    .C1(_08172_),
    .Y(_08180_));
 sky130_fd_sc_hd__a211o_1 _16710_ (.A1(_07948_),
    .A2(_07964_),
    .B1(_07963_),
    .C1(_07955_),
    .X(_08181_));
 sky130_fd_sc_hd__and4_1 _16711_ (.A(_07965_),
    .B(_08178_),
    .C(_08180_),
    .D(_08181_),
    .X(_08182_));
 sky130_fd_sc_hd__nand4_2 _16712_ (.A(_07965_),
    .B(_08178_),
    .C(_08180_),
    .D(_08181_),
    .Y(_08183_));
 sky130_fd_sc_hd__o21ai_2 _16713_ (.A1(_08149_),
    .A2(_08150_),
    .B1(_08151_),
    .Y(_08184_));
 sky130_fd_sc_hd__o211ai_4 _16714_ (.A1(_08179_),
    .A2(_08182_),
    .B1(_08184_),
    .C1(_08153_),
    .Y(_08185_));
 sky130_fd_sc_hd__and3_1 _16715_ (.A(_07948_),
    .B(_07965_),
    .C(_07976_),
    .X(_08186_));
 sky130_fd_sc_hd__nor2_1 _16716_ (.A(_07977_),
    .B(_08186_),
    .Y(_08187_));
 sky130_fd_sc_hd__a211o_1 _16717_ (.A1(_08153_),
    .A2(_08184_),
    .B1(_08182_),
    .C1(_08179_),
    .X(_08188_));
 sky130_fd_sc_hd__nand3_4 _16718_ (.A(_08185_),
    .B(_08187_),
    .C(_08188_),
    .Y(_08189_));
 sky130_fd_sc_hd__a211o_1 _16719_ (.A1(_08185_),
    .A2(_08189_),
    .B1(_08157_),
    .C1(_08158_),
    .X(_08190_));
 sky130_fd_sc_hd__o211ai_2 _16720_ (.A1(_08157_),
    .A2(_08158_),
    .B1(_08185_),
    .C1(_08189_),
    .Y(_08191_));
 sky130_fd_sc_hd__and3_1 _16721_ (.A(_07977_),
    .B(_08190_),
    .C(_08191_),
    .X(_08192_));
 sky130_fd_sc_hd__a21oi_1 _16722_ (.A1(_08190_),
    .A2(_08191_),
    .B1(_07977_),
    .Y(_08193_));
 sky130_fd_sc_hd__nor2_2 _16723_ (.A(_08192_),
    .B(_08193_),
    .Y(_08194_));
 sky130_fd_sc_hd__nand4_1 _16724_ (.A(net621),
    .B(net189),
    .C(net268),
    .D(net273),
    .Y(_08195_));
 sky130_fd_sc_hd__and2_1 _16725_ (.A(net186),
    .B(net278),
    .X(_08196_));
 sky130_fd_sc_hd__a22o_1 _16726_ (.A1(net622),
    .A2(net268),
    .B1(net273),
    .B2(net189),
    .X(_08197_));
 sky130_fd_sc_hd__nand3_1 _16727_ (.A(_08195_),
    .B(_08196_),
    .C(_08197_),
    .Y(_08198_));
 sky130_fd_sc_hd__a21bo_1 _16728_ (.A1(_08196_),
    .A2(_08197_),
    .B1_N(_08195_),
    .X(_08199_));
 sky130_fd_sc_hd__a21o_1 _16729_ (.A1(_08159_),
    .A2(_08161_),
    .B1(_08160_),
    .X(_08200_));
 sky130_fd_sc_hd__nand3_1 _16730_ (.A(_08162_),
    .B(_08199_),
    .C(_08200_),
    .Y(_08201_));
 sky130_fd_sc_hd__a21o_1 _16731_ (.A1(_08162_),
    .A2(_08200_),
    .B1(_08199_),
    .X(_08202_));
 sky130_fd_sc_hd__nand2_1 _16732_ (.A(net171),
    .B(net288),
    .Y(_08203_));
 sky130_fd_sc_hd__and3_1 _16733_ (.A(net182),
    .B(net176),
    .C(net283),
    .X(_08204_));
 sky130_fd_sc_hd__and4_1 _16734_ (.A(net182),
    .B(net177),
    .C(net278),
    .D(net283),
    .X(_08205_));
 sky130_fd_sc_hd__a22o_1 _16735_ (.A1(net182),
    .A2(net278),
    .B1(net283),
    .B2(net177),
    .X(_08206_));
 sky130_fd_sc_hd__and2b_1 _16736_ (.A_N(_08205_),
    .B(_08206_),
    .X(_08207_));
 sky130_fd_sc_hd__xnor2_1 _16737_ (.A(_08203_),
    .B(_08207_),
    .Y(_08208_));
 sky130_fd_sc_hd__nand3_1 _16738_ (.A(_08201_),
    .B(_08202_),
    .C(_08208_),
    .Y(_08209_));
 sky130_fd_sc_hd__a21bo_1 _16739_ (.A1(_08202_),
    .A2(_08208_),
    .B1_N(_08201_),
    .X(_08210_));
 sky130_fd_sc_hd__a21o_1 _16740_ (.A1(_08165_),
    .A2(_08166_),
    .B1(_08168_),
    .X(_08211_));
 sky130_fd_sc_hd__nand3_4 _16741_ (.A(_08169_),
    .B(_08210_),
    .C(_08211_),
    .Y(_08212_));
 sky130_fd_sc_hd__a21o_1 _16742_ (.A1(_08169_),
    .A2(_08211_),
    .B1(_08210_),
    .X(_08213_));
 sky130_fd_sc_hd__and4_1 _16743_ (.A(net166),
    .B(net160),
    .C(net294),
    .D(net298),
    .X(_08214_));
 sky130_fd_sc_hd__nand2_1 _16744_ (.A(\mul1.b[8] ),
    .B(net303),
    .Y(_08215_));
 sky130_fd_sc_hd__a22o_1 _16745_ (.A1(net166),
    .A2(net294),
    .B1(net298),
    .B2(net160),
    .X(_08216_));
 sky130_fd_sc_hd__and2b_1 _16746_ (.A_N(_08214_),
    .B(_08216_),
    .X(_08217_));
 sky130_fd_sc_hd__a31o_1 _16747_ (.A1(\mul1.b[8] ),
    .A2(net303),
    .A3(_08216_),
    .B1(_08214_),
    .X(_08218_));
 sky130_fd_sc_hd__a31o_1 _16748_ (.A1(net171),
    .A2(net288),
    .A3(_08206_),
    .B1(_08205_),
    .X(_08219_));
 sky130_fd_sc_hd__xnor2_2 _16749_ (.A(_07923_),
    .B(_07925_),
    .Y(_08220_));
 sky130_fd_sc_hd__nand2_1 _16750_ (.A(_08219_),
    .B(_08220_),
    .Y(_08221_));
 sky130_fd_sc_hd__xor2_2 _16751_ (.A(_08219_),
    .B(_08220_),
    .X(_08222_));
 sky130_fd_sc_hd__nand2_1 _16752_ (.A(_08218_),
    .B(_08222_),
    .Y(_08223_));
 sky130_fd_sc_hd__xor2_2 _16753_ (.A(_08218_),
    .B(_08222_),
    .X(_08224_));
 sky130_fd_sc_hd__nand3_4 _16754_ (.A(_08212_),
    .B(_08213_),
    .C(_08224_),
    .Y(_08225_));
 sky130_fd_sc_hd__a21oi_2 _16755_ (.A1(_08172_),
    .A2(_08173_),
    .B1(_08174_),
    .Y(_08226_));
 sky130_fd_sc_hd__a211oi_4 _16756_ (.A1(_08212_),
    .A2(_08225_),
    .B1(_08226_),
    .C1(_08175_),
    .Y(_08227_));
 sky130_fd_sc_hd__o211a_1 _16757_ (.A1(_08175_),
    .A2(_08226_),
    .B1(_08225_),
    .C1(_08212_),
    .X(_08228_));
 sky130_fd_sc_hd__xnor2_2 _16758_ (.A(_07951_),
    .B(_07953_),
    .Y(_08229_));
 sky130_fd_sc_hd__and4_1 _16759_ (.A(net150),
    .B(net145),
    .C(net309),
    .D(net315),
    .X(_08230_));
 sky130_fd_sc_hd__nand2_1 _16760_ (.A(net141),
    .B(net319),
    .Y(_08231_));
 sky130_fd_sc_hd__a22o_1 _16761_ (.A1(net150),
    .A2(net309),
    .B1(net315),
    .B2(net145),
    .X(_08232_));
 sky130_fd_sc_hd__and2b_1 _16762_ (.A_N(_08230_),
    .B(_08232_),
    .X(_08233_));
 sky130_fd_sc_hd__a31o_1 _16763_ (.A1(net141),
    .A2(net319),
    .A3(_08232_),
    .B1(_08230_),
    .X(_08234_));
 sky130_fd_sc_hd__and2_1 _16764_ (.A(_08229_),
    .B(_08234_),
    .X(_08235_));
 sky130_fd_sc_hd__xor2_2 _16765_ (.A(_08229_),
    .B(_08234_),
    .X(_08236_));
 sky130_fd_sc_hd__a22o_1 _16766_ (.A1(net136),
    .A2(net319),
    .B1(net323),
    .B2(net131),
    .X(_08237_));
 sky130_fd_sc_hd__inv_2 _16767_ (.A(_08237_),
    .Y(_08238_));
 sky130_fd_sc_hd__and4_1 _16768_ (.A(net136),
    .B(net131),
    .C(net319),
    .D(net323),
    .X(_08239_));
 sky130_fd_sc_hd__nor2_1 _16769_ (.A(_08238_),
    .B(_08239_),
    .Y(_08240_));
 sky130_fd_sc_hd__and2_1 _16770_ (.A(_08236_),
    .B(_08240_),
    .X(_08241_));
 sky130_fd_sc_hd__xnor2_1 _16771_ (.A(_07956_),
    .B(_07962_),
    .Y(_08242_));
 sky130_fd_sc_hd__a21o_1 _16772_ (.A1(_08221_),
    .A2(_08223_),
    .B1(_08242_),
    .X(_08243_));
 sky130_fd_sc_hd__nand3_1 _16773_ (.A(_08221_),
    .B(_08223_),
    .C(_08242_),
    .Y(_08244_));
 sky130_fd_sc_hd__o211ai_2 _16774_ (.A1(_08235_),
    .A2(_08241_),
    .B1(_08243_),
    .C1(_08244_),
    .Y(_08245_));
 sky130_fd_sc_hd__a211o_1 _16775_ (.A1(_08243_),
    .A2(_08244_),
    .B1(_08235_),
    .C1(_08241_),
    .X(_08246_));
 sky130_fd_sc_hd__and4bb_2 _16776_ (.A_N(_08227_),
    .B_N(_08228_),
    .C(_08245_),
    .D(_08246_),
    .X(_08247_));
 sky130_fd_sc_hd__a22o_1 _16777_ (.A1(_08178_),
    .A2(_08180_),
    .B1(_08181_),
    .B2(_07965_),
    .X(_08248_));
 sky130_fd_sc_hd__o211a_1 _16778_ (.A1(_08227_),
    .A2(_08247_),
    .B1(_08248_),
    .C1(_08183_),
    .X(_08249_));
 sky130_fd_sc_hd__o211ai_2 _16779_ (.A1(_08227_),
    .A2(_08247_),
    .B1(_08248_),
    .C1(_08183_),
    .Y(_08250_));
 sky130_fd_sc_hd__a211o_1 _16780_ (.A1(_08183_),
    .A2(_08248_),
    .B1(_08247_),
    .C1(_08227_),
    .X(_08251_));
 sky130_fd_sc_hd__xnor2_1 _16781_ (.A(_07966_),
    .B(_07967_),
    .Y(_08252_));
 sky130_fd_sc_hd__a21oi_2 _16782_ (.A1(_08243_),
    .A2(_08245_),
    .B1(_08252_),
    .Y(_08253_));
 sky130_fd_sc_hd__and3_1 _16783_ (.A(_08243_),
    .B(_08245_),
    .C(_08252_),
    .X(_08254_));
 sky130_fd_sc_hd__nor2_1 _16784_ (.A(_08253_),
    .B(_08254_),
    .Y(_08255_));
 sky130_fd_sc_hd__and3_2 _16785_ (.A(_08250_),
    .B(_08251_),
    .C(_08255_),
    .X(_08256_));
 sky130_fd_sc_hd__a21o_1 _16786_ (.A1(_08185_),
    .A2(_08188_),
    .B1(_08187_),
    .X(_08257_));
 sky130_fd_sc_hd__o211ai_4 _16787_ (.A1(_08249_),
    .A2(_08256_),
    .B1(_08257_),
    .C1(_08189_),
    .Y(_08258_));
 sky130_fd_sc_hd__a211o_1 _16788_ (.A1(_08189_),
    .A2(_08257_),
    .B1(_08256_),
    .C1(_08249_),
    .X(_08259_));
 sky130_fd_sc_hd__nand3_4 _16789_ (.A(_08253_),
    .B(_08258_),
    .C(_08259_),
    .Y(_08260_));
 sky130_fd_sc_hd__nand2_2 _16790_ (.A(_08258_),
    .B(_08260_),
    .Y(_08261_));
 sky130_fd_sc_hd__nand2_1 _16791_ (.A(_08194_),
    .B(_08261_),
    .Y(_08262_));
 sky130_fd_sc_hd__xnor2_4 _16792_ (.A(_08194_),
    .B(_08261_),
    .Y(_08263_));
 sky130_fd_sc_hd__a21o_1 _16793_ (.A1(_08258_),
    .A2(_08259_),
    .B1(_08253_),
    .X(_08264_));
 sky130_fd_sc_hd__nand4_2 _16794_ (.A(net621),
    .B(net188),
    .C(net273),
    .D(net278),
    .Y(_08265_));
 sky130_fd_sc_hd__and2_1 _16795_ (.A(net186),
    .B(net283),
    .X(_08266_));
 sky130_fd_sc_hd__a22o_1 _16796_ (.A1(net621),
    .A2(net273),
    .B1(net278),
    .B2(net188),
    .X(_08267_));
 sky130_fd_sc_hd__nand3_1 _16797_ (.A(_08265_),
    .B(_08266_),
    .C(_08267_),
    .Y(_08268_));
 sky130_fd_sc_hd__a21bo_1 _16798_ (.A1(_08266_),
    .A2(_08267_),
    .B1_N(_08265_),
    .X(_08269_));
 sky130_fd_sc_hd__a21o_1 _16799_ (.A1(_08195_),
    .A2(_08197_),
    .B1(_08196_),
    .X(_08270_));
 sky130_fd_sc_hd__nand3_1 _16800_ (.A(_08198_),
    .B(_08269_),
    .C(_08270_),
    .Y(_08271_));
 sky130_fd_sc_hd__a21o_1 _16801_ (.A1(_08198_),
    .A2(_08270_),
    .B1(_08269_),
    .X(_08272_));
 sky130_fd_sc_hd__nand2_1 _16802_ (.A(net172),
    .B(net293),
    .Y(_08273_));
 sky130_fd_sc_hd__a22o_1 _16803_ (.A1(net182),
    .A2(net283),
    .B1(net288),
    .B2(net177),
    .X(_08274_));
 sky130_fd_sc_hd__a21bo_1 _16804_ (.A1(net288),
    .A2(_08204_),
    .B1_N(_08274_),
    .X(_08275_));
 sky130_fd_sc_hd__xor2_1 _16805_ (.A(_08273_),
    .B(_08275_),
    .X(_08276_));
 sky130_fd_sc_hd__nand3_1 _16806_ (.A(_08271_),
    .B(_08272_),
    .C(_08276_),
    .Y(_08277_));
 sky130_fd_sc_hd__a21bo_1 _16807_ (.A1(_08272_),
    .A2(_08276_),
    .B1_N(_08271_),
    .X(_08278_));
 sky130_fd_sc_hd__a21o_1 _16808_ (.A1(_08201_),
    .A2(_08202_),
    .B1(_08208_),
    .X(_08279_));
 sky130_fd_sc_hd__and3_1 _16809_ (.A(_08209_),
    .B(_08278_),
    .C(_08279_),
    .X(_08280_));
 sky130_fd_sc_hd__nand3_1 _16810_ (.A(_08209_),
    .B(_08278_),
    .C(_08279_),
    .Y(_08281_));
 sky130_fd_sc_hd__a21o_1 _16811_ (.A1(_08209_),
    .A2(_08279_),
    .B1(_08278_),
    .X(_08282_));
 sky130_fd_sc_hd__and4_1 _16812_ (.A(net165),
    .B(net159),
    .C(net299),
    .D(net304),
    .X(_08283_));
 sky130_fd_sc_hd__nand4_1 _16813_ (.A(net166),
    .B(net159),
    .C(net299),
    .D(net304),
    .Y(_08284_));
 sky130_fd_sc_hd__a22o_1 _16814_ (.A1(net166),
    .A2(net299),
    .B1(net303),
    .B2(net159),
    .X(_08285_));
 sky130_fd_sc_hd__and4_1 _16815_ (.A(net155),
    .B(net309),
    .C(_08284_),
    .D(_08285_),
    .X(_08286_));
 sky130_fd_sc_hd__nor2_1 _16816_ (.A(_08283_),
    .B(_08286_),
    .Y(_08287_));
 sky130_fd_sc_hd__a32o_1 _16817_ (.A1(net171),
    .A2(net293),
    .A3(_08274_),
    .B1(_08204_),
    .B2(net288),
    .X(_08288_));
 sky130_fd_sc_hd__xnor2_1 _16818_ (.A(_08215_),
    .B(_08217_),
    .Y(_08289_));
 sky130_fd_sc_hd__nand2_1 _16819_ (.A(_08288_),
    .B(_08289_),
    .Y(_08290_));
 sky130_fd_sc_hd__xor2_1 _16820_ (.A(_08288_),
    .B(_08289_),
    .X(_08291_));
 sky130_fd_sc_hd__nand2b_1 _16821_ (.A_N(_08287_),
    .B(_08291_),
    .Y(_08292_));
 sky130_fd_sc_hd__xnor2_1 _16822_ (.A(_08287_),
    .B(_08291_),
    .Y(_08293_));
 sky130_fd_sc_hd__and3_1 _16823_ (.A(_08281_),
    .B(_08282_),
    .C(_08293_),
    .X(_08294_));
 sky130_fd_sc_hd__a21o_1 _16824_ (.A1(_08212_),
    .A2(_08213_),
    .B1(_08224_),
    .X(_08295_));
 sky130_fd_sc_hd__o211a_1 _16825_ (.A1(_08280_),
    .A2(_08294_),
    .B1(_08295_),
    .C1(_08225_),
    .X(_08296_));
 sky130_fd_sc_hd__inv_2 _16826_ (.A(_08296_),
    .Y(_08297_));
 sky130_fd_sc_hd__a211oi_2 _16827_ (.A1(_08225_),
    .A2(_08295_),
    .B1(_08294_),
    .C1(_08280_),
    .Y(_08298_));
 sky130_fd_sc_hd__xnor2_1 _16828_ (.A(_08231_),
    .B(_08233_),
    .Y(_08299_));
 sky130_fd_sc_hd__and4_1 _16829_ (.A(net150),
    .B(net145),
    .C(net314),
    .D(net320),
    .X(_08300_));
 sky130_fd_sc_hd__inv_2 _16830_ (.A(_08300_),
    .Y(_08301_));
 sky130_fd_sc_hd__a22o_1 _16831_ (.A1(net150),
    .A2(net314),
    .B1(net320),
    .B2(net145),
    .X(_08302_));
 sky130_fd_sc_hd__and4b_1 _16832_ (.A_N(_08300_),
    .B(_08302_),
    .C(net141),
    .D(net322),
    .X(_08303_));
 sky130_fd_sc_hd__or2_1 _16833_ (.A(_08300_),
    .B(_08303_),
    .X(_08304_));
 sky130_fd_sc_hd__nand2_1 _16834_ (.A(_08299_),
    .B(_08304_),
    .Y(_08305_));
 sky130_fd_sc_hd__nand2_1 _16835_ (.A(net136),
    .B(net323),
    .Y(_08306_));
 sky130_fd_sc_hd__xor2_1 _16836_ (.A(_08299_),
    .B(_08304_),
    .X(_08307_));
 sky130_fd_sc_hd__nand2b_1 _16837_ (.A_N(_08306_),
    .B(_08307_),
    .Y(_08308_));
 sky130_fd_sc_hd__xnor2_2 _16838_ (.A(_08236_),
    .B(_08240_),
    .Y(_08309_));
 sky130_fd_sc_hd__a21oi_4 _16839_ (.A1(_08290_),
    .A2(_08292_),
    .B1(_08309_),
    .Y(_08310_));
 sky130_fd_sc_hd__and3_1 _16840_ (.A(_08290_),
    .B(_08292_),
    .C(_08309_),
    .X(_08311_));
 sky130_fd_sc_hd__a211oi_4 _16841_ (.A1(_08305_),
    .A2(_08308_),
    .B1(_08310_),
    .C1(_08311_),
    .Y(_08312_));
 sky130_fd_sc_hd__o211a_1 _16842_ (.A1(_08310_),
    .A2(_08311_),
    .B1(_08305_),
    .C1(_08308_),
    .X(_08313_));
 sky130_fd_sc_hd__nor4_1 _16843_ (.A(_08296_),
    .B(_08298_),
    .C(_08312_),
    .D(_08313_),
    .Y(_08314_));
 sky130_fd_sc_hd__or4_1 _16844_ (.A(_08296_),
    .B(_08298_),
    .C(_08312_),
    .D(_08313_),
    .X(_08315_));
 sky130_fd_sc_hd__a2bb2oi_1 _16845_ (.A1_N(_08227_),
    .A2_N(_08228_),
    .B1(_08245_),
    .B2(_08246_),
    .Y(_08316_));
 sky130_fd_sc_hd__a211o_2 _16846_ (.A1(_08297_),
    .A2(_08315_),
    .B1(_08316_),
    .C1(_08247_),
    .X(_08317_));
 sky130_fd_sc_hd__o211ai_2 _16847_ (.A1(_08247_),
    .A2(_08316_),
    .B1(_08315_),
    .C1(_08297_),
    .Y(_08318_));
 sky130_fd_sc_hd__o21ai_2 _16848_ (.A1(_08310_),
    .A2(_08312_),
    .B1(_08239_),
    .Y(_08319_));
 sky130_fd_sc_hd__or3_1 _16849_ (.A(_08239_),
    .B(_08310_),
    .C(_08312_),
    .X(_08320_));
 sky130_fd_sc_hd__and2_1 _16850_ (.A(_08319_),
    .B(_08320_),
    .X(_08321_));
 sky130_fd_sc_hd__nand3_2 _16851_ (.A(_08317_),
    .B(_08318_),
    .C(_08321_),
    .Y(_08322_));
 sky130_fd_sc_hd__a21oi_2 _16852_ (.A1(_08250_),
    .A2(_08251_),
    .B1(_08255_),
    .Y(_08323_));
 sky130_fd_sc_hd__a211oi_4 _16853_ (.A1(_08317_),
    .A2(_08322_),
    .B1(_08323_),
    .C1(_08256_),
    .Y(_08324_));
 sky130_fd_sc_hd__o211a_1 _16854_ (.A1(_08256_),
    .A2(_08323_),
    .B1(_08322_),
    .C1(_08317_),
    .X(_08325_));
 sky130_fd_sc_hd__nor3_2 _16855_ (.A(_08319_),
    .B(_08324_),
    .C(_08325_),
    .Y(_08326_));
 sky130_fd_sc_hd__o211ai_4 _16856_ (.A1(_08324_),
    .A2(_08326_),
    .B1(_08260_),
    .C1(_08264_),
    .Y(_08327_));
 sky130_fd_sc_hd__o21a_1 _16857_ (.A1(_08324_),
    .A2(_08325_),
    .B1(_08319_),
    .X(_08328_));
 sky130_fd_sc_hd__a21o_1 _16858_ (.A1(_08317_),
    .A2(_08318_),
    .B1(_08321_),
    .X(_08329_));
 sky130_fd_sc_hd__and2_1 _16859_ (.A(_08322_),
    .B(_08329_),
    .X(_08330_));
 sky130_fd_sc_hd__nand4_1 _16860_ (.A(net621),
    .B(net188),
    .C(net278),
    .D(net283),
    .Y(_08331_));
 sky130_fd_sc_hd__and2_1 _16861_ (.A(net186),
    .B(net288),
    .X(_08332_));
 sky130_fd_sc_hd__a22o_1 _16862_ (.A1(net621),
    .A2(net278),
    .B1(net283),
    .B2(net188),
    .X(_08333_));
 sky130_fd_sc_hd__nand3_1 _16863_ (.A(_08331_),
    .B(_08332_),
    .C(_08333_),
    .Y(_08334_));
 sky130_fd_sc_hd__a21bo_1 _16864_ (.A1(_08332_),
    .A2(_08333_),
    .B1_N(_08331_),
    .X(_08335_));
 sky130_fd_sc_hd__a21o_1 _16865_ (.A1(_08265_),
    .A2(_08267_),
    .B1(_08266_),
    .X(_08336_));
 sky130_fd_sc_hd__nand3_1 _16866_ (.A(_08268_),
    .B(_08335_),
    .C(_08336_),
    .Y(_08337_));
 sky130_fd_sc_hd__a22o_1 _16867_ (.A1(net181),
    .A2(net288),
    .B1(net293),
    .B2(net176),
    .X(_08338_));
 sky130_fd_sc_hd__and3_1 _16868_ (.A(net182),
    .B(net176),
    .C(net288),
    .X(_08339_));
 sky130_fd_sc_hd__a21bo_1 _16869_ (.A1(net293),
    .A2(_08339_),
    .B1_N(_08338_),
    .X(_08340_));
 sky130_fd_sc_hd__nand2_1 _16870_ (.A(net172),
    .B(net298),
    .Y(_08341_));
 sky130_fd_sc_hd__xor2_2 _16871_ (.A(_08340_),
    .B(_08341_),
    .X(_08342_));
 sky130_fd_sc_hd__a21o_1 _16872_ (.A1(_08268_),
    .A2(_08336_),
    .B1(_08335_),
    .X(_08343_));
 sky130_fd_sc_hd__nand3_1 _16873_ (.A(_08337_),
    .B(_08342_),
    .C(_08343_),
    .Y(_08344_));
 sky130_fd_sc_hd__a21bo_1 _16874_ (.A1(_08342_),
    .A2(_08343_),
    .B1_N(_08337_),
    .X(_08345_));
 sky130_fd_sc_hd__a21o_1 _16875_ (.A1(_08271_),
    .A2(_08272_),
    .B1(_08276_),
    .X(_08346_));
 sky130_fd_sc_hd__nand3_2 _16876_ (.A(_08277_),
    .B(_08345_),
    .C(_08346_),
    .Y(_08347_));
 sky130_fd_sc_hd__a32o_1 _16877_ (.A1(net171),
    .A2(net298),
    .A3(_08338_),
    .B1(_08339_),
    .B2(net293),
    .X(_08348_));
 sky130_fd_sc_hd__a22o_1 _16878_ (.A1(net155),
    .A2(net309),
    .B1(_08284_),
    .B2(_08285_),
    .X(_08349_));
 sky130_fd_sc_hd__and2b_1 _16879_ (.A_N(_08286_),
    .B(_08349_),
    .X(_08350_));
 sky130_fd_sc_hd__and2_1 _16880_ (.A(_08348_),
    .B(_08350_),
    .X(_08351_));
 sky130_fd_sc_hd__xor2_1 _16881_ (.A(_08348_),
    .B(_08350_),
    .X(_08352_));
 sky130_fd_sc_hd__and3_1 _16882_ (.A(net165),
    .B(net159),
    .C(net303),
    .X(_08353_));
 sky130_fd_sc_hd__nand2_1 _16883_ (.A(net155),
    .B(net313),
    .Y(_08354_));
 sky130_fd_sc_hd__a22o_1 _16884_ (.A1(net165),
    .A2(net303),
    .B1(net308),
    .B2(net159),
    .X(_08355_));
 sky130_fd_sc_hd__a21bo_1 _16885_ (.A1(net308),
    .A2(_08353_),
    .B1_N(_08355_),
    .X(_08356_));
 sky130_fd_sc_hd__o2bb2a_1 _16886_ (.A1_N(net308),
    .A2_N(_08353_),
    .B1(_08354_),
    .B2(_08356_),
    .X(_08357_));
 sky130_fd_sc_hd__inv_2 _16887_ (.A(_08357_),
    .Y(_08358_));
 sky130_fd_sc_hd__xnor2_1 _16888_ (.A(_08352_),
    .B(_08357_),
    .Y(_08359_));
 sky130_fd_sc_hd__a21o_1 _16889_ (.A1(_08277_),
    .A2(_08346_),
    .B1(_08345_),
    .X(_08360_));
 sky130_fd_sc_hd__nand3_2 _16890_ (.A(_08347_),
    .B(_08359_),
    .C(_08360_),
    .Y(_08361_));
 sky130_fd_sc_hd__a21oi_1 _16891_ (.A1(_08281_),
    .A2(_08282_),
    .B1(_08293_),
    .Y(_08362_));
 sky130_fd_sc_hd__a211o_1 _16892_ (.A1(_08347_),
    .A2(_08361_),
    .B1(_08362_),
    .C1(_08294_),
    .X(_08363_));
 sky130_fd_sc_hd__a21oi_1 _16893_ (.A1(_08352_),
    .A2(_08358_),
    .B1(_08351_),
    .Y(_08364_));
 sky130_fd_sc_hd__xnor2_1 _16894_ (.A(_08306_),
    .B(_08307_),
    .Y(_08365_));
 sky130_fd_sc_hd__and2b_1 _16895_ (.A_N(_08364_),
    .B(_08365_),
    .X(_08366_));
 sky130_fd_sc_hd__xnor2_1 _16896_ (.A(_08364_),
    .B(_08365_),
    .Y(_08367_));
 sky130_fd_sc_hd__a22oi_1 _16897_ (.A1(net141),
    .A2(net325),
    .B1(_08301_),
    .B2(_08302_),
    .Y(_08368_));
 sky130_fd_sc_hd__nor2_1 _16898_ (.A(_08303_),
    .B(_08368_),
    .Y(_08369_));
 sky130_fd_sc_hd__and4_1 _16899_ (.A(net150),
    .B(net145),
    .C(net320),
    .D(net325),
    .X(_08370_));
 sky130_fd_sc_hd__and2_1 _16900_ (.A(_08369_),
    .B(_08370_),
    .X(_08371_));
 sky130_fd_sc_hd__xor2_1 _16901_ (.A(_08367_),
    .B(_08371_),
    .X(_08372_));
 sky130_fd_sc_hd__o211ai_1 _16902_ (.A1(_08294_),
    .A2(_08362_),
    .B1(_08361_),
    .C1(_08347_),
    .Y(_08373_));
 sky130_fd_sc_hd__nand3_1 _16903_ (.A(_08363_),
    .B(_08372_),
    .C(_08373_),
    .Y(_08374_));
 sky130_fd_sc_hd__o22a_1 _16904_ (.A1(_08296_),
    .A2(_08298_),
    .B1(_08312_),
    .B2(_08313_),
    .X(_08375_));
 sky130_fd_sc_hd__a211o_1 _16905_ (.A1(_08363_),
    .A2(_08374_),
    .B1(_08375_),
    .C1(_08314_),
    .X(_08376_));
 sky130_fd_sc_hd__a21o_1 _16906_ (.A1(_08367_),
    .A2(_08371_),
    .B1(_08366_),
    .X(_08377_));
 sky130_fd_sc_hd__o211ai_2 _16907_ (.A1(_08314_),
    .A2(_08375_),
    .B1(_08374_),
    .C1(_08363_),
    .Y(_08378_));
 sky130_fd_sc_hd__nand3_1 _16908_ (.A(_08376_),
    .B(_08377_),
    .C(_08378_),
    .Y(_08379_));
 sky130_fd_sc_hd__nand2_1 _16909_ (.A(_08376_),
    .B(_08379_),
    .Y(_08380_));
 sky130_fd_sc_hd__and4bb_1 _16910_ (.A_N(_08326_),
    .B_N(_08328_),
    .C(_08330_),
    .D(_08380_),
    .X(_08381_));
 sky130_fd_sc_hd__a211o_1 _16911_ (.A1(_08260_),
    .A2(_08264_),
    .B1(_08324_),
    .C1(_08326_),
    .X(_08382_));
 sky130_fd_sc_hd__nand2_1 _16912_ (.A(_08381_),
    .B(_08382_),
    .Y(_08383_));
 sky130_fd_sc_hd__a21bo_1 _16913_ (.A1(_08381_),
    .A2(_08382_),
    .B1_N(_08327_),
    .X(_08384_));
 sky130_fd_sc_hd__xor2_4 _16914_ (.A(_08263_),
    .B(_08384_),
    .X(_08385_));
 sky130_fd_sc_hd__a21o_1 _16915_ (.A1(_08376_),
    .A2(_08378_),
    .B1(_08377_),
    .X(_08386_));
 sky130_fd_sc_hd__nand2_1 _16916_ (.A(_08379_),
    .B(_08386_),
    .Y(_08387_));
 sky130_fd_sc_hd__nand4_2 _16917_ (.A(net621),
    .B(net188),
    .C(net283),
    .D(net288),
    .Y(_08388_));
 sky130_fd_sc_hd__and2_1 _16918_ (.A(net186),
    .B(net293),
    .X(_08389_));
 sky130_fd_sc_hd__a22o_1 _16919_ (.A1(net621),
    .A2(net283),
    .B1(net288),
    .B2(net188),
    .X(_08390_));
 sky130_fd_sc_hd__nand3_1 _16920_ (.A(_08388_),
    .B(_08389_),
    .C(_08390_),
    .Y(_08391_));
 sky130_fd_sc_hd__a21bo_1 _16921_ (.A1(_08389_),
    .A2(_08390_),
    .B1_N(_08388_),
    .X(_08392_));
 sky130_fd_sc_hd__a21o_1 _16922_ (.A1(_08331_),
    .A2(_08333_),
    .B1(_08332_),
    .X(_08393_));
 sky130_fd_sc_hd__nand3_1 _16923_ (.A(_08334_),
    .B(_08392_),
    .C(_08393_),
    .Y(_08394_));
 sky130_fd_sc_hd__a22oi_2 _16924_ (.A1(net181),
    .A2(net293),
    .B1(net298),
    .B2(net176),
    .Y(_08395_));
 sky130_fd_sc_hd__and4_1 _16925_ (.A(net181),
    .B(net176),
    .C(net293),
    .D(net298),
    .X(_08396_));
 sky130_fd_sc_hd__nor2_1 _16926_ (.A(_08395_),
    .B(_08396_),
    .Y(_08397_));
 sky130_fd_sc_hd__nand2_1 _16927_ (.A(net171),
    .B(net303),
    .Y(_08398_));
 sky130_fd_sc_hd__xnor2_1 _16928_ (.A(_08397_),
    .B(_08398_),
    .Y(_08399_));
 sky130_fd_sc_hd__a21o_1 _16929_ (.A1(_08334_),
    .A2(_08393_),
    .B1(_08392_),
    .X(_08400_));
 sky130_fd_sc_hd__nand3_1 _16930_ (.A(_08394_),
    .B(_08399_),
    .C(_08400_),
    .Y(_08401_));
 sky130_fd_sc_hd__a21bo_1 _16931_ (.A1(_08399_),
    .A2(_08400_),
    .B1_N(_08394_),
    .X(_08402_));
 sky130_fd_sc_hd__a21o_1 _16932_ (.A1(_08337_),
    .A2(_08343_),
    .B1(_08342_),
    .X(_08403_));
 sky130_fd_sc_hd__and3_2 _16933_ (.A(_08344_),
    .B(_08402_),
    .C(_08403_),
    .X(_08404_));
 sky130_fd_sc_hd__o21ba_1 _16934_ (.A1(_08395_),
    .A2(_08398_),
    .B1_N(_08396_),
    .X(_08405_));
 sky130_fd_sc_hd__xor2_2 _16935_ (.A(_08354_),
    .B(_08356_),
    .X(_08406_));
 sky130_fd_sc_hd__nand2b_1 _16936_ (.A_N(_08405_),
    .B(_08406_),
    .Y(_08407_));
 sky130_fd_sc_hd__xnor2_2 _16937_ (.A(_08405_),
    .B(_08406_),
    .Y(_08408_));
 sky130_fd_sc_hd__and4_1 _16938_ (.A(net165),
    .B(net159),
    .C(net308),
    .D(net313),
    .X(_08409_));
 sky130_fd_sc_hd__nand2_1 _16939_ (.A(net155),
    .B(net318),
    .Y(_08410_));
 sky130_fd_sc_hd__a22o_1 _16940_ (.A1(net165),
    .A2(net308),
    .B1(net313),
    .B2(net159),
    .X(_08411_));
 sky130_fd_sc_hd__and2b_1 _16941_ (.A_N(_08409_),
    .B(_08411_),
    .X(_08412_));
 sky130_fd_sc_hd__a31o_1 _16942_ (.A1(net155),
    .A2(net318),
    .A3(_08411_),
    .B1(_08409_),
    .X(_08413_));
 sky130_fd_sc_hd__xnor2_2 _16943_ (.A(_08408_),
    .B(_08413_),
    .Y(_08414_));
 sky130_fd_sc_hd__a21oi_1 _16944_ (.A1(_08344_),
    .A2(_08403_),
    .B1(_08402_),
    .Y(_08415_));
 sky130_fd_sc_hd__nor3_2 _16945_ (.A(_08404_),
    .B(_08414_),
    .C(_08415_),
    .Y(_08416_));
 sky130_fd_sc_hd__or3_1 _16946_ (.A(_08404_),
    .B(_08414_),
    .C(_08415_),
    .X(_08417_));
 sky130_fd_sc_hd__a21o_1 _16947_ (.A1(_08347_),
    .A2(_08360_),
    .B1(_08359_),
    .X(_08418_));
 sky130_fd_sc_hd__o211ai_4 _16948_ (.A1(_08404_),
    .A2(_08416_),
    .B1(_08418_),
    .C1(_08361_),
    .Y(_08419_));
 sky130_fd_sc_hd__inv_2 _16949_ (.A(_08419_),
    .Y(_08420_));
 sky130_fd_sc_hd__a21bo_1 _16950_ (.A1(_08408_),
    .A2(_08413_),
    .B1_N(_08407_),
    .X(_08421_));
 sky130_fd_sc_hd__nor2_1 _16951_ (.A(_08369_),
    .B(_08370_),
    .Y(_08422_));
 sky130_fd_sc_hd__or2_1 _16952_ (.A(_08371_),
    .B(_08422_),
    .X(_08423_));
 sky130_fd_sc_hd__and2b_1 _16953_ (.A_N(_08423_),
    .B(_08421_),
    .X(_08424_));
 sky130_fd_sc_hd__xnor2_1 _16954_ (.A(_08421_),
    .B(_08423_),
    .Y(_08425_));
 sky130_fd_sc_hd__a211o_1 _16955_ (.A1(_08361_),
    .A2(_08418_),
    .B1(_08416_),
    .C1(_08404_),
    .X(_08426_));
 sky130_fd_sc_hd__nand3_1 _16956_ (.A(_08419_),
    .B(_08425_),
    .C(_08426_),
    .Y(_08427_));
 sky130_fd_sc_hd__a21o_1 _16957_ (.A1(_08363_),
    .A2(_08373_),
    .B1(_08372_),
    .X(_08428_));
 sky130_fd_sc_hd__and2_1 _16958_ (.A(_08374_),
    .B(_08428_),
    .X(_08429_));
 sky130_fd_sc_hd__a21bo_1 _16959_ (.A1(_08419_),
    .A2(_08427_),
    .B1_N(_08429_),
    .X(_08430_));
 sky130_fd_sc_hd__a211o_1 _16960_ (.A1(_08425_),
    .A2(_08426_),
    .B1(_08429_),
    .C1(_08420_),
    .X(_08431_));
 sky130_fd_sc_hd__nand3_2 _16961_ (.A(_08424_),
    .B(_08430_),
    .C(_08431_),
    .Y(_08432_));
 sky130_fd_sc_hd__a21o_1 _16962_ (.A1(_08430_),
    .A2(_08432_),
    .B1(_08387_),
    .X(_08433_));
 sky130_fd_sc_hd__a21o_1 _16963_ (.A1(_08430_),
    .A2(_08431_),
    .B1(_08424_),
    .X(_08434_));
 sky130_fd_sc_hd__a21o_1 _16964_ (.A1(_08419_),
    .A2(_08426_),
    .B1(_08425_),
    .X(_08435_));
 sky130_fd_sc_hd__o21ai_1 _16965_ (.A1(_08404_),
    .A2(_08415_),
    .B1(_08414_),
    .Y(_08436_));
 sky130_fd_sc_hd__a21o_1 _16966_ (.A1(_08394_),
    .A2(_08400_),
    .B1(_08399_),
    .X(_08437_));
 sky130_fd_sc_hd__a21o_1 _16967_ (.A1(_08388_),
    .A2(_08390_),
    .B1(_08389_),
    .X(_08438_));
 sky130_fd_sc_hd__nand4_1 _16968_ (.A(net621),
    .B(net188),
    .C(net288),
    .D(net293),
    .Y(_08439_));
 sky130_fd_sc_hd__and2_1 _16969_ (.A(net186),
    .B(net298),
    .X(_08440_));
 sky130_fd_sc_hd__a22o_1 _16970_ (.A1(net621),
    .A2(net288),
    .B1(net293),
    .B2(net188),
    .X(_08441_));
 sky130_fd_sc_hd__nand3_1 _16971_ (.A(_08439_),
    .B(_08440_),
    .C(_08441_),
    .Y(_08442_));
 sky130_fd_sc_hd__a21bo_1 _16972_ (.A1(_08440_),
    .A2(_08441_),
    .B1_N(_08439_),
    .X(_08443_));
 sky130_fd_sc_hd__nand3_1 _16973_ (.A(_08391_),
    .B(_08438_),
    .C(_08443_),
    .Y(_08444_));
 sky130_fd_sc_hd__a22oi_1 _16974_ (.A1(net181),
    .A2(net298),
    .B1(net303),
    .B2(net176),
    .Y(_08445_));
 sky130_fd_sc_hd__and4_1 _16975_ (.A(net181),
    .B(net176),
    .C(net298),
    .D(net303),
    .X(_08446_));
 sky130_fd_sc_hd__o2bb2a_1 _16976_ (.A1_N(net171),
    .A2_N(net308),
    .B1(_08445_),
    .B2(_08446_),
    .X(_08447_));
 sky130_fd_sc_hd__and4bb_1 _16977_ (.A_N(_08445_),
    .B_N(_08446_),
    .C(net171),
    .D(net308),
    .X(_08448_));
 sky130_fd_sc_hd__nor2_1 _16978_ (.A(_08447_),
    .B(_08448_),
    .Y(_08449_));
 sky130_fd_sc_hd__a21o_1 _16979_ (.A1(_08391_),
    .A2(_08438_),
    .B1(_08443_),
    .X(_08450_));
 sky130_fd_sc_hd__nand3_1 _16980_ (.A(_08444_),
    .B(_08449_),
    .C(_08450_),
    .Y(_08451_));
 sky130_fd_sc_hd__a21bo_1 _16981_ (.A1(_08449_),
    .A2(_08450_),
    .B1_N(_08444_),
    .X(_08452_));
 sky130_fd_sc_hd__and3_2 _16982_ (.A(_08401_),
    .B(_08437_),
    .C(_08452_),
    .X(_08453_));
 sky130_fd_sc_hd__nor2_1 _16983_ (.A(_08446_),
    .B(_08448_),
    .Y(_08454_));
 sky130_fd_sc_hd__xnor2_1 _16984_ (.A(_08410_),
    .B(_08412_),
    .Y(_08455_));
 sky130_fd_sc_hd__and2b_1 _16985_ (.A_N(_08454_),
    .B(_08455_),
    .X(_08456_));
 sky130_fd_sc_hd__xnor2_1 _16986_ (.A(_08454_),
    .B(_08455_),
    .Y(_08457_));
 sky130_fd_sc_hd__and4_1 _16987_ (.A(net165),
    .B(net159),
    .C(net313),
    .D(net318),
    .X(_08458_));
 sky130_fd_sc_hd__a22oi_1 _16988_ (.A1(net165),
    .A2(net313),
    .B1(net318),
    .B2(net159),
    .Y(_08459_));
 sky130_fd_sc_hd__and4bb_1 _16989_ (.A_N(_08458_),
    .B_N(_08459_),
    .C(net155),
    .D(net322),
    .X(_08460_));
 sky130_fd_sc_hd__nor2_1 _16990_ (.A(_08458_),
    .B(_08460_),
    .Y(_08461_));
 sky130_fd_sc_hd__and2b_1 _16991_ (.A_N(_08461_),
    .B(_08457_),
    .X(_08462_));
 sky130_fd_sc_hd__xor2_1 _16992_ (.A(_08457_),
    .B(_08461_),
    .X(_08463_));
 sky130_fd_sc_hd__a21oi_1 _16993_ (.A1(_08401_),
    .A2(_08437_),
    .B1(_08452_),
    .Y(_08464_));
 sky130_fd_sc_hd__nor3_2 _16994_ (.A(_08453_),
    .B(_08463_),
    .C(_08464_),
    .Y(_08465_));
 sky130_fd_sc_hd__o211a_1 _16995_ (.A1(_08453_),
    .A2(_08465_),
    .B1(_08417_),
    .C1(_08436_),
    .X(_08466_));
 sky130_fd_sc_hd__a22oi_1 _16996_ (.A1(net150),
    .A2(net320),
    .B1(net325),
    .B2(net145),
    .Y(_08467_));
 sky130_fd_sc_hd__nor2_1 _16997_ (.A(_08370_),
    .B(_08467_),
    .Y(_08468_));
 sky130_fd_sc_hd__o21ai_1 _16998_ (.A1(_08456_),
    .A2(_08462_),
    .B1(_08468_),
    .Y(_08469_));
 sky130_fd_sc_hd__or3_1 _16999_ (.A(_08456_),
    .B(_08462_),
    .C(_08468_),
    .X(_08470_));
 sky130_fd_sc_hd__nand2_1 _17000_ (.A(_08469_),
    .B(_08470_),
    .Y(_08471_));
 sky130_fd_sc_hd__a211oi_2 _17001_ (.A1(_08417_),
    .A2(_08436_),
    .B1(_08453_),
    .C1(_08465_),
    .Y(_08472_));
 sky130_fd_sc_hd__nor3_2 _17002_ (.A(_08466_),
    .B(_08471_),
    .C(_08472_),
    .Y(_08473_));
 sky130_fd_sc_hd__o211a_1 _17003_ (.A1(_08466_),
    .A2(_08473_),
    .B1(_08427_),
    .C1(_08435_),
    .X(_08474_));
 sky130_fd_sc_hd__a211oi_1 _17004_ (.A1(_08427_),
    .A2(_08435_),
    .B1(_08466_),
    .C1(_08473_),
    .Y(_08475_));
 sky130_fd_sc_hd__nor3_1 _17005_ (.A(_08469_),
    .B(_08474_),
    .C(_08475_),
    .Y(_08476_));
 sky130_fd_sc_hd__o211ai_1 _17006_ (.A1(_08474_),
    .A2(_08476_),
    .B1(_08432_),
    .C1(_08434_),
    .Y(_08477_));
 sky130_fd_sc_hd__a211o_1 _17007_ (.A1(_08432_),
    .A2(_08434_),
    .B1(_08474_),
    .C1(_08476_),
    .X(_08478_));
 sky130_fd_sc_hd__o21a_1 _17008_ (.A1(_08474_),
    .A2(_08475_),
    .B1(_08469_),
    .X(_08479_));
 sky130_fd_sc_hd__o21a_1 _17009_ (.A1(_08466_),
    .A2(_08472_),
    .B1(_08471_),
    .X(_08480_));
 sky130_fd_sc_hd__o21a_1 _17010_ (.A1(_08453_),
    .A2(_08464_),
    .B1(_08463_),
    .X(_08481_));
 sky130_fd_sc_hd__a21o_1 _17011_ (.A1(_08444_),
    .A2(_08450_),
    .B1(_08449_),
    .X(_08482_));
 sky130_fd_sc_hd__a21o_1 _17012_ (.A1(_08439_),
    .A2(_08441_),
    .B1(_08440_),
    .X(_08483_));
 sky130_fd_sc_hd__nand4_2 _17013_ (.A(net622),
    .B(net188),
    .C(net293),
    .D(net298),
    .Y(_08484_));
 sky130_fd_sc_hd__and2_1 _17014_ (.A(net186),
    .B(net303),
    .X(_08485_));
 sky130_fd_sc_hd__a22o_1 _17015_ (.A1(net621),
    .A2(net293),
    .B1(net298),
    .B2(net188),
    .X(_08486_));
 sky130_fd_sc_hd__nand3_1 _17016_ (.A(_08484_),
    .B(_08485_),
    .C(_08486_),
    .Y(_08487_));
 sky130_fd_sc_hd__a21bo_1 _17017_ (.A1(_08485_),
    .A2(_08486_),
    .B1_N(_08484_),
    .X(_08488_));
 sky130_fd_sc_hd__nand3_1 _17018_ (.A(_08442_),
    .B(_08483_),
    .C(_08488_),
    .Y(_08489_));
 sky130_fd_sc_hd__and4_1 _17019_ (.A(net181),
    .B(net176),
    .C(net303),
    .D(net308),
    .X(_08490_));
 sky130_fd_sc_hd__a22o_1 _17020_ (.A1(net181),
    .A2(net303),
    .B1(net308),
    .B2(net176),
    .X(_08491_));
 sky130_fd_sc_hd__and2b_1 _17021_ (.A_N(_08490_),
    .B(_08491_),
    .X(_08492_));
 sky130_fd_sc_hd__nand2_1 _17022_ (.A(net171),
    .B(net313),
    .Y(_08493_));
 sky130_fd_sc_hd__xnor2_1 _17023_ (.A(_08492_),
    .B(_08493_),
    .Y(_08494_));
 sky130_fd_sc_hd__a21o_1 _17024_ (.A1(_08442_),
    .A2(_08483_),
    .B1(_08488_),
    .X(_08495_));
 sky130_fd_sc_hd__nand3_1 _17025_ (.A(_08489_),
    .B(_08494_),
    .C(_08495_),
    .Y(_08496_));
 sky130_fd_sc_hd__a21bo_1 _17026_ (.A1(_08494_),
    .A2(_08495_),
    .B1_N(_08489_),
    .X(_08497_));
 sky130_fd_sc_hd__and3_1 _17027_ (.A(_08451_),
    .B(_08482_),
    .C(_08497_),
    .X(_08498_));
 sky130_fd_sc_hd__nand3_1 _17028_ (.A(_08451_),
    .B(_08482_),
    .C(_08497_),
    .Y(_08499_));
 sky130_fd_sc_hd__and4_1 _17029_ (.A(net165),
    .B(net159),
    .C(net318),
    .D(net322),
    .X(_08500_));
 sky130_fd_sc_hd__inv_2 _17030_ (.A(_08500_),
    .Y(_08501_));
 sky130_fd_sc_hd__a31o_1 _17031_ (.A1(net171),
    .A2(net313),
    .A3(_08491_),
    .B1(_08490_),
    .X(_08502_));
 sky130_fd_sc_hd__o2bb2a_1 _17032_ (.A1_N(net155),
    .A2_N(net322),
    .B1(_08458_),
    .B2(_08459_),
    .X(_08503_));
 sky130_fd_sc_hd__nor2_1 _17033_ (.A(_08460_),
    .B(_08503_),
    .Y(_08504_));
 sky130_fd_sc_hd__nand2_1 _17034_ (.A(_08502_),
    .B(_08504_),
    .Y(_08505_));
 sky130_fd_sc_hd__xnor2_1 _17035_ (.A(_08502_),
    .B(_08504_),
    .Y(_08506_));
 sky130_fd_sc_hd__xnor2_1 _17036_ (.A(_08501_),
    .B(_08506_),
    .Y(_08507_));
 sky130_fd_sc_hd__a21oi_1 _17037_ (.A1(_08451_),
    .A2(_08482_),
    .B1(_08497_),
    .Y(_08508_));
 sky130_fd_sc_hd__or3_2 _17038_ (.A(_08498_),
    .B(_08507_),
    .C(_08508_),
    .X(_08509_));
 sky130_fd_sc_hd__a211oi_1 _17039_ (.A1(_08499_),
    .A2(_08509_),
    .B1(_08465_),
    .C1(_08481_),
    .Y(_08510_));
 sky130_fd_sc_hd__a211o_1 _17040_ (.A1(_08499_),
    .A2(_08509_),
    .B1(_08465_),
    .C1(_08481_),
    .X(_08511_));
 sky130_fd_sc_hd__nand2_1 _17041_ (.A(net150),
    .B(net322),
    .Y(_08512_));
 sky130_fd_sc_hd__o21a_1 _17042_ (.A1(_08501_),
    .A2(_08506_),
    .B1(_08505_),
    .X(_08513_));
 sky130_fd_sc_hd__nor2_1 _17043_ (.A(_08512_),
    .B(_08513_),
    .Y(_08514_));
 sky130_fd_sc_hd__xnor2_1 _17044_ (.A(_08512_),
    .B(_08513_),
    .Y(_08515_));
 sky130_fd_sc_hd__o211a_1 _17045_ (.A1(_08465_),
    .A2(_08481_),
    .B1(_08499_),
    .C1(_08509_),
    .X(_08516_));
 sky130_fd_sc_hd__or3_2 _17046_ (.A(_08510_),
    .B(_08515_),
    .C(_08516_),
    .X(_08517_));
 sky130_fd_sc_hd__a211o_1 _17047_ (.A1(_08511_),
    .A2(_08517_),
    .B1(_08473_),
    .C1(_08480_),
    .X(_08518_));
 sky130_fd_sc_hd__o211ai_2 _17048_ (.A1(_08473_),
    .A2(_08480_),
    .B1(_08511_),
    .C1(_08517_),
    .Y(_08519_));
 sky130_fd_sc_hd__nand3_2 _17049_ (.A(_08514_),
    .B(_08518_),
    .C(_08519_),
    .Y(_08520_));
 sky130_fd_sc_hd__a211o_1 _17050_ (.A1(_08518_),
    .A2(_08520_),
    .B1(_08476_),
    .C1(_08479_),
    .X(_08521_));
 sky130_fd_sc_hd__a21o_1 _17051_ (.A1(_08518_),
    .A2(_08519_),
    .B1(_08514_),
    .X(_08522_));
 sky130_fd_sc_hd__and4_1 _17052_ (.A(net181),
    .B(net176),
    .C(net308),
    .D(net313),
    .X(_08523_));
 sky130_fd_sc_hd__a22o_1 _17053_ (.A1(net181),
    .A2(net308),
    .B1(net313),
    .B2(net176),
    .X(_08524_));
 sky130_fd_sc_hd__and2b_1 _17054_ (.A_N(_08523_),
    .B(_08524_),
    .X(_08525_));
 sky130_fd_sc_hd__nand2_1 _17055_ (.A(net171),
    .B(net318),
    .Y(_08526_));
 sky130_fd_sc_hd__a31o_1 _17056_ (.A1(net171),
    .A2(net318),
    .A3(_08524_),
    .B1(_08523_),
    .X(_08527_));
 sky130_fd_sc_hd__a22o_1 _17057_ (.A1(net165),
    .A2(net318),
    .B1(net322),
    .B2(net159),
    .X(_08528_));
 sky130_fd_sc_hd__and2_1 _17058_ (.A(_08501_),
    .B(_08528_),
    .X(_08529_));
 sky130_fd_sc_hd__nand2_1 _17059_ (.A(_08527_),
    .B(_08529_),
    .Y(_08530_));
 sky130_fd_sc_hd__o21ai_1 _17060_ (.A1(_08498_),
    .A2(_08508_),
    .B1(_08507_),
    .Y(_08531_));
 sky130_fd_sc_hd__a21o_1 _17061_ (.A1(_08489_),
    .A2(_08495_),
    .B1(_08494_),
    .X(_08532_));
 sky130_fd_sc_hd__a21o_1 _17062_ (.A1(_08484_),
    .A2(_08486_),
    .B1(_08485_),
    .X(_08533_));
 sky130_fd_sc_hd__nand4_2 _17063_ (.A(net622),
    .B(net189),
    .C(net299),
    .D(net304),
    .Y(_08534_));
 sky130_fd_sc_hd__and2_1 _17064_ (.A(net186),
    .B(net309),
    .X(_08535_));
 sky130_fd_sc_hd__a22o_1 _17065_ (.A1(net622),
    .A2(net299),
    .B1(net304),
    .B2(net189),
    .X(_08536_));
 sky130_fd_sc_hd__nand3_1 _17066_ (.A(_08534_),
    .B(_08535_),
    .C(_08536_),
    .Y(_08537_));
 sky130_fd_sc_hd__a21bo_1 _17067_ (.A1(_08535_),
    .A2(_08536_),
    .B1_N(_08534_),
    .X(_08538_));
 sky130_fd_sc_hd__nand3_1 _17068_ (.A(_08487_),
    .B(_08533_),
    .C(_08538_),
    .Y(_08539_));
 sky130_fd_sc_hd__xnor2_1 _17069_ (.A(_08525_),
    .B(_08526_),
    .Y(_08540_));
 sky130_fd_sc_hd__a21o_1 _17070_ (.A1(_08487_),
    .A2(_08533_),
    .B1(_08538_),
    .X(_08541_));
 sky130_fd_sc_hd__nand3_1 _17071_ (.A(_08539_),
    .B(_08540_),
    .C(_08541_),
    .Y(_08542_));
 sky130_fd_sc_hd__a21bo_1 _17072_ (.A1(_08540_),
    .A2(_08541_),
    .B1_N(_08539_),
    .X(_08543_));
 sky130_fd_sc_hd__and3_1 _17073_ (.A(_08496_),
    .B(_08532_),
    .C(_08543_),
    .X(_08544_));
 sky130_fd_sc_hd__or2_1 _17074_ (.A(_08527_),
    .B(_08529_),
    .X(_08545_));
 sky130_fd_sc_hd__nand2_1 _17075_ (.A(_08530_),
    .B(_08545_),
    .Y(_08546_));
 sky130_fd_sc_hd__a21oi_1 _17076_ (.A1(_08496_),
    .A2(_08532_),
    .B1(_08543_),
    .Y(_08547_));
 sky130_fd_sc_hd__nor3_1 _17077_ (.A(_08544_),
    .B(_08546_),
    .C(_08547_),
    .Y(_08548_));
 sky130_fd_sc_hd__or3_1 _17078_ (.A(_08544_),
    .B(_08546_),
    .C(_08547_),
    .X(_08549_));
 sky130_fd_sc_hd__o211a_1 _17079_ (.A1(_08544_),
    .A2(_08548_),
    .B1(_08509_),
    .C1(_08531_),
    .X(_08550_));
 sky130_fd_sc_hd__a211oi_1 _17080_ (.A1(_08509_),
    .A2(_08531_),
    .B1(_08544_),
    .C1(_08548_),
    .Y(_08551_));
 sky130_fd_sc_hd__or3_1 _17081_ (.A(_08530_),
    .B(_08550_),
    .C(_08551_),
    .X(_08552_));
 sky130_fd_sc_hd__o21ai_1 _17082_ (.A1(_08550_),
    .A2(_08551_),
    .B1(_08530_),
    .Y(_08553_));
 sky130_fd_sc_hd__o21ai_1 _17083_ (.A1(_08544_),
    .A2(_08547_),
    .B1(_08546_),
    .Y(_08554_));
 sky130_fd_sc_hd__a21o_1 _17084_ (.A1(_08539_),
    .A2(_08541_),
    .B1(_08540_),
    .X(_08555_));
 sky130_fd_sc_hd__a21o_1 _17085_ (.A1(_08534_),
    .A2(_08536_),
    .B1(_08535_),
    .X(_08556_));
 sky130_fd_sc_hd__and4_1 _17086_ (.A(net622),
    .B(net189),
    .C(net304),
    .D(net309),
    .X(_08557_));
 sky130_fd_sc_hd__nand2_1 _17087_ (.A(net186),
    .B(net313),
    .Y(_08558_));
 sky130_fd_sc_hd__a22oi_2 _17088_ (.A1(net622),
    .A2(net304),
    .B1(net309),
    .B2(net189),
    .Y(_08559_));
 sky130_fd_sc_hd__or3_1 _17089_ (.A(_08557_),
    .B(_08558_),
    .C(_08559_),
    .X(_08560_));
 sky130_fd_sc_hd__o21bai_1 _17090_ (.A1(_08558_),
    .A2(_08559_),
    .B1_N(_08557_),
    .Y(_08561_));
 sky130_fd_sc_hd__nand3_1 _17091_ (.A(_08537_),
    .B(_08556_),
    .C(_08561_),
    .Y(_08562_));
 sky130_fd_sc_hd__a22oi_1 _17092_ (.A1(net181),
    .A2(net313),
    .B1(net318),
    .B2(net176),
    .Y(_08563_));
 sky130_fd_sc_hd__and4_1 _17093_ (.A(net181),
    .B(net176),
    .C(net313),
    .D(net318),
    .X(_08564_));
 sky130_fd_sc_hd__nor2_1 _17094_ (.A(_08563_),
    .B(_08564_),
    .Y(_08565_));
 sky130_fd_sc_hd__nand2_1 _17095_ (.A(net171),
    .B(net322),
    .Y(_08566_));
 sky130_fd_sc_hd__and3_1 _17096_ (.A(net171),
    .B(net322),
    .C(_08565_),
    .X(_08567_));
 sky130_fd_sc_hd__xnor2_1 _17097_ (.A(_08565_),
    .B(_08566_),
    .Y(_08568_));
 sky130_fd_sc_hd__a21o_1 _17098_ (.A1(_08537_),
    .A2(_08556_),
    .B1(_08561_),
    .X(_08569_));
 sky130_fd_sc_hd__nand3_1 _17099_ (.A(_08562_),
    .B(_08568_),
    .C(_08569_),
    .Y(_08570_));
 sky130_fd_sc_hd__a21bo_1 _17100_ (.A1(_08568_),
    .A2(_08569_),
    .B1_N(_08562_),
    .X(_08571_));
 sky130_fd_sc_hd__and3_1 _17101_ (.A(_08542_),
    .B(_08555_),
    .C(_08571_),
    .X(_08572_));
 sky130_fd_sc_hd__o211a_1 _17102_ (.A1(_08564_),
    .A2(_08567_),
    .B1(net165),
    .C1(net322),
    .X(_08573_));
 sky130_fd_sc_hd__a211oi_1 _17103_ (.A1(net165),
    .A2(net322),
    .B1(_08564_),
    .C1(_08567_),
    .Y(_08574_));
 sky130_fd_sc_hd__or2_1 _17104_ (.A(_08573_),
    .B(_08574_),
    .X(_08575_));
 sky130_fd_sc_hd__a21oi_1 _17105_ (.A1(_08542_),
    .A2(_08555_),
    .B1(_08571_),
    .Y(_08576_));
 sky130_fd_sc_hd__nor3_1 _17106_ (.A(_08572_),
    .B(_08575_),
    .C(_08576_),
    .Y(_08577_));
 sky130_fd_sc_hd__o211a_1 _17107_ (.A1(_08572_),
    .A2(_08577_),
    .B1(_08549_),
    .C1(_08554_),
    .X(_08578_));
 sky130_fd_sc_hd__o211ai_1 _17108_ (.A1(_08572_),
    .A2(_08577_),
    .B1(_08549_),
    .C1(_08554_),
    .Y(_08579_));
 sky130_fd_sc_hd__a211o_1 _17109_ (.A1(_08549_),
    .A2(_08554_),
    .B1(_08572_),
    .C1(_08577_),
    .X(_08580_));
 sky130_fd_sc_hd__and3_1 _17110_ (.A(_08573_),
    .B(_08579_),
    .C(_08580_),
    .X(_08581_));
 sky130_fd_sc_hd__o211a_1 _17111_ (.A1(_08578_),
    .A2(_08581_),
    .B1(_08552_),
    .C1(_08553_),
    .X(_08582_));
 sky130_fd_sc_hd__o21ai_1 _17112_ (.A1(_08510_),
    .A2(_08516_),
    .B1(_08515_),
    .Y(_08583_));
 sky130_fd_sc_hd__o21bai_1 _17113_ (.A1(_08530_),
    .A2(_08551_),
    .B1_N(_08550_),
    .Y(_08584_));
 sky130_fd_sc_hd__and3_1 _17114_ (.A(_08517_),
    .B(_08583_),
    .C(_08584_),
    .X(_08585_));
 sky130_fd_sc_hd__a21o_1 _17115_ (.A1(_08517_),
    .A2(_08583_),
    .B1(_08584_),
    .X(_08586_));
 sky130_fd_sc_hd__o21a_1 _17116_ (.A1(_08582_),
    .A2(_08585_),
    .B1(_08586_),
    .X(_08587_));
 sky130_fd_sc_hd__nand3_1 _17117_ (.A(_08520_),
    .B(_08522_),
    .C(_08587_),
    .Y(_08588_));
 sky130_fd_sc_hd__a21oi_1 _17118_ (.A1(_08579_),
    .A2(_08580_),
    .B1(_08573_),
    .Y(_08589_));
 sky130_fd_sc_hd__o21a_1 _17119_ (.A1(_08572_),
    .A2(_08576_),
    .B1(_08575_),
    .X(_08590_));
 sky130_fd_sc_hd__or2_1 _17120_ (.A(_08577_),
    .B(_08590_),
    .X(_08591_));
 sky130_fd_sc_hd__a21o_1 _17121_ (.A1(_08562_),
    .A2(_08569_),
    .B1(_08568_),
    .X(_08592_));
 sky130_fd_sc_hd__o21ai_1 _17122_ (.A1(_08557_),
    .A2(_08559_),
    .B1(_08558_),
    .Y(_08593_));
 sky130_fd_sc_hd__and4_1 _17123_ (.A(net622),
    .B(net189),
    .C(net309),
    .D(net313),
    .X(_08594_));
 sky130_fd_sc_hd__nand4_1 _17124_ (.A(net622),
    .B(net189),
    .C(net308),
    .D(net314),
    .Y(_08595_));
 sky130_fd_sc_hd__a22o_1 _17125_ (.A1(net622),
    .A2(net309),
    .B1(net314),
    .B2(net189),
    .X(_08596_));
 sky130_fd_sc_hd__and4_1 _17126_ (.A(net186),
    .B(net320),
    .C(_08595_),
    .D(_08596_),
    .X(_08597_));
 sky130_fd_sc_hd__o211ai_2 _17127_ (.A1(_08594_),
    .A2(_08597_),
    .B1(_08560_),
    .C1(_08593_),
    .Y(_08598_));
 sky130_fd_sc_hd__a22oi_1 _17128_ (.A1(net181),
    .A2(net318),
    .B1(net322),
    .B2(net176),
    .Y(_08599_));
 sky130_fd_sc_hd__and4_1 _17129_ (.A(net181),
    .B(net176),
    .C(net318),
    .D(net322),
    .X(_08600_));
 sky130_fd_sc_hd__nor2_1 _17130_ (.A(_08599_),
    .B(_08600_),
    .Y(_08601_));
 sky130_fd_sc_hd__a211o_1 _17131_ (.A1(_08560_),
    .A2(_08593_),
    .B1(_08594_),
    .C1(_08597_),
    .X(_08602_));
 sky130_fd_sc_hd__nand3_1 _17132_ (.A(_08598_),
    .B(_08601_),
    .C(_08602_),
    .Y(_08603_));
 sky130_fd_sc_hd__nand2_1 _17133_ (.A(_08598_),
    .B(_08603_),
    .Y(_08604_));
 sky130_fd_sc_hd__nand3_1 _17134_ (.A(_08570_),
    .B(_08592_),
    .C(_08604_),
    .Y(_08605_));
 sky130_fd_sc_hd__a21o_1 _17135_ (.A1(_08570_),
    .A2(_08592_),
    .B1(_08604_),
    .X(_08606_));
 sky130_fd_sc_hd__a21boi_1 _17136_ (.A1(_08600_),
    .A2(_08606_),
    .B1_N(_08605_),
    .Y(_08607_));
 sky130_fd_sc_hd__a21oi_1 _17137_ (.A1(_08605_),
    .A2(_08606_),
    .B1(_08600_),
    .Y(_08608_));
 sky130_fd_sc_hd__a21o_1 _17138_ (.A1(_08598_),
    .A2(_08602_),
    .B1(_08601_),
    .X(_08609_));
 sky130_fd_sc_hd__a22oi_1 _17139_ (.A1(net186),
    .A2(net318),
    .B1(_08595_),
    .B2(_08596_),
    .Y(_08610_));
 sky130_fd_sc_hd__nor2_1 _17140_ (.A(_08597_),
    .B(_08610_),
    .Y(_08611_));
 sky130_fd_sc_hd__and4_1 _17141_ (.A(net621),
    .B(net188),
    .C(net314),
    .D(net320),
    .X(_08612_));
 sky130_fd_sc_hd__a22o_1 _17142_ (.A1(net621),
    .A2(net313),
    .B1(net318),
    .B2(net188),
    .X(_08613_));
 sky130_fd_sc_hd__a31o_1 _17143_ (.A1(net186),
    .A2(net322),
    .A3(_08613_),
    .B1(_08612_),
    .X(_08614_));
 sky130_fd_sc_hd__nand2_1 _17144_ (.A(net181),
    .B(net322),
    .Y(_08615_));
 sky130_fd_sc_hd__or2_1 _17145_ (.A(net186),
    .B(net313),
    .X(_08616_));
 sky130_fd_sc_hd__and4_1 _17146_ (.A(net622),
    .B(net189),
    .C(net318),
    .D(net322),
    .X(_08617_));
 sky130_fd_sc_hd__a21bo_1 _17147_ (.A1(_08558_),
    .A2(_08616_),
    .B1_N(_08617_),
    .X(_08618_));
 sky130_fd_sc_hd__o2bb2a_1 _17148_ (.A1_N(_08615_),
    .A2_N(_08618_),
    .B1(_08611_),
    .B2(_08614_),
    .X(_08619_));
 sky130_fd_sc_hd__and2_1 _17149_ (.A(_08611_),
    .B(_08614_),
    .X(_08620_));
 sky130_fd_sc_hd__nor2_1 _17150_ (.A(_08615_),
    .B(_08618_),
    .Y(_08621_));
 sky130_fd_sc_hd__o311a_1 _17151_ (.A1(_08619_),
    .A2(_08620_),
    .A3(_08621_),
    .B1(_08609_),
    .C1(_08603_),
    .X(_08622_));
 sky130_fd_sc_hd__a21oi_1 _17152_ (.A1(_08620_),
    .A2(_08621_),
    .B1(_08622_),
    .Y(_08623_));
 sky130_fd_sc_hd__a31o_1 _17153_ (.A1(_08600_),
    .A2(_08605_),
    .A3(_08606_),
    .B1(_08623_),
    .X(_08624_));
 sky130_fd_sc_hd__o22a_1 _17154_ (.A1(_08591_),
    .A2(_08607_),
    .B1(_08608_),
    .B2(_08624_),
    .X(_08625_));
 sky130_fd_sc_hd__a2111o_1 _17155_ (.A1(_08591_),
    .A2(_08607_),
    .B1(_08625_),
    .C1(_08589_),
    .D1(_08581_),
    .X(_08626_));
 sky130_fd_sc_hd__and3_1 _17156_ (.A(_08552_),
    .B(_08553_),
    .C(_08578_),
    .X(_08627_));
 sky130_fd_sc_hd__a21o_1 _17157_ (.A1(_08552_),
    .A2(_08553_),
    .B1(_08578_),
    .X(_08628_));
 sky130_fd_sc_hd__nand2_1 _17158_ (.A(_08586_),
    .B(_08628_),
    .Y(_08629_));
 sky130_fd_sc_hd__or4_1 _17159_ (.A(_08585_),
    .B(_08626_),
    .C(_08627_),
    .D(_08629_),
    .X(_08630_));
 sky130_fd_sc_hd__a21oi_1 _17160_ (.A1(_08520_),
    .A2(_08522_),
    .B1(_08587_),
    .Y(_08631_));
 sky130_fd_sc_hd__o211a_1 _17161_ (.A1(_08476_),
    .A2(_08479_),
    .B1(_08518_),
    .C1(_08520_),
    .X(_08632_));
 sky130_fd_sc_hd__a211o_1 _17162_ (.A1(_08588_),
    .A2(_08630_),
    .B1(_08631_),
    .C1(_08632_),
    .X(_08633_));
 sky130_fd_sc_hd__a21bo_1 _17163_ (.A1(_08521_),
    .A2(_08633_),
    .B1_N(_08478_),
    .X(_08634_));
 sky130_fd_sc_hd__a32o_1 _17164_ (.A1(_08387_),
    .A2(_08430_),
    .A3(_08432_),
    .B1(_08477_),
    .B2(_08634_),
    .X(_08635_));
 sky130_fd_sc_hd__and3_1 _17165_ (.A(_08260_),
    .B(_08264_),
    .C(_08324_),
    .X(_08636_));
 sky130_fd_sc_hd__a21oi_1 _17166_ (.A1(_08260_),
    .A2(_08264_),
    .B1(_08324_),
    .Y(_08637_));
 sky130_fd_sc_hd__xnor2_1 _17167_ (.A(_08330_),
    .B(_08380_),
    .Y(_08638_));
 sky130_fd_sc_hd__or3_1 _17168_ (.A(_08326_),
    .B(_08328_),
    .C(_08638_),
    .X(_08639_));
 sky130_fd_sc_hd__or3_1 _17169_ (.A(_08636_),
    .B(_08637_),
    .C(_08639_),
    .X(_08640_));
 sky130_fd_sc_hd__a21o_2 _17170_ (.A1(_08433_),
    .A2(_08635_),
    .B1(_08640_),
    .X(_08641_));
 sky130_fd_sc_hd__xnor2_4 _17171_ (.A(_08385_),
    .B(_08641_),
    .Y(_08642_));
 sky130_fd_sc_hd__nor2_1 _17172_ (.A(_03049_),
    .B(_08642_),
    .Y(_08643_));
 sky130_fd_sc_hd__nor2_1 _17173_ (.A(net43),
    .B(_03792_),
    .Y(_08644_));
 sky130_fd_sc_hd__a21o_1 _17174_ (.A1(net802),
    .A2(net7),
    .B1(_03056_),
    .X(_08645_));
 sky130_fd_sc_hd__o32a_1 _17175_ (.A1(_08643_),
    .A2(_08644_),
    .A3(_08645_),
    .B1(net3),
    .B2(net840),
    .X(_00299_));
 sky130_fd_sc_hd__a21bo_2 _17176_ (.A1(_07977_),
    .A2(_08191_),
    .B1_N(_08190_),
    .X(_08646_));
 sky130_fd_sc_hd__o21a_2 _17177_ (.A1(_07974_),
    .A2(_08023_),
    .B1(_08022_),
    .X(_08647_));
 sky130_fd_sc_hd__nor2_1 _17178_ (.A(_08053_),
    .B(_08055_),
    .Y(_08648_));
 sky130_fd_sc_hd__a31o_1 _17179_ (.A1(net114),
    .A2(net323),
    .A3(_08013_),
    .B1(_08012_),
    .X(_08649_));
 sky130_fd_sc_hd__a31oi_2 _17180_ (.A1(net127),
    .A2(net310),
    .A3(_08041_),
    .B1(_08040_),
    .Y(_08650_));
 sky130_fd_sc_hd__nand4_1 _17181_ (.A(net310),
    .B(net315),
    .C(net122),
    .D(net117),
    .Y(_08651_));
 sky130_fd_sc_hd__a22o_1 _17182_ (.A1(net310),
    .A2(net122),
    .B1(net117),
    .B2(net315),
    .X(_08652_));
 sky130_fd_sc_hd__and4_1 _17183_ (.A(net319),
    .B(net114),
    .C(_08651_),
    .D(_08652_),
    .X(_08653_));
 sky130_fd_sc_hd__a22o_1 _17184_ (.A1(net319),
    .A2(net114),
    .B1(_08651_),
    .B2(_08652_),
    .X(_08654_));
 sky130_fd_sc_hd__and2b_1 _17185_ (.A_N(_08653_),
    .B(_08654_),
    .X(_08655_));
 sky130_fd_sc_hd__or3b_1 _17186_ (.A(_08650_),
    .B(_08653_),
    .C_N(_08654_),
    .X(_08656_));
 sky130_fd_sc_hd__xnor2_2 _17187_ (.A(_08650_),
    .B(_08655_),
    .Y(_08657_));
 sky130_fd_sc_hd__xnor2_2 _17188_ (.A(_08649_),
    .B(_08657_),
    .Y(_08658_));
 sky130_fd_sc_hd__o21ai_2 _17189_ (.A1(_07970_),
    .A2(_08018_),
    .B1(_08016_),
    .Y(_08659_));
 sky130_fd_sc_hd__nor2_1 _17190_ (.A(_08658_),
    .B(_08659_),
    .Y(_08660_));
 sky130_fd_sc_hd__xor2_2 _17191_ (.A(_08658_),
    .B(_08659_),
    .X(_08661_));
 sky130_fd_sc_hd__nand2_1 _17192_ (.A(net323),
    .B(net107),
    .Y(_08662_));
 sky130_fd_sc_hd__and3_1 _17193_ (.A(net323),
    .B(net107),
    .C(_08661_),
    .X(_08663_));
 sky130_fd_sc_hd__xnor2_2 _17194_ (.A(_08661_),
    .B(_08662_),
    .Y(_08664_));
 sky130_fd_sc_hd__and2b_1 _17195_ (.A_N(_08648_),
    .B(_08664_),
    .X(_08665_));
 sky130_fd_sc_hd__xnor2_2 _17196_ (.A(_08648_),
    .B(_08664_),
    .Y(_08666_));
 sky130_fd_sc_hd__nand2_1 _17197_ (.A(_07972_),
    .B(_08019_),
    .Y(_08667_));
 sky130_fd_sc_hd__xnor2_1 _17198_ (.A(_08666_),
    .B(_08667_),
    .Y(_08668_));
 sky130_fd_sc_hd__nand2_1 _17199_ (.A(_08049_),
    .B(_08051_),
    .Y(_08669_));
 sky130_fd_sc_hd__and4_1 _17200_ (.A(net295),
    .B(net300),
    .C(net136),
    .D(net131),
    .X(_08670_));
 sky130_fd_sc_hd__inv_2 _17201_ (.A(_08670_),
    .Y(_08671_));
 sky130_fd_sc_hd__a22o_1 _17202_ (.A1(net295),
    .A2(net136),
    .B1(net131),
    .B2(net300),
    .X(_08672_));
 sky130_fd_sc_hd__and4b_1 _17203_ (.A_N(_08670_),
    .B(_08672_),
    .C(net305),
    .D(net127),
    .X(_08673_));
 sky130_fd_sc_hd__a22oi_1 _17204_ (.A1(net305),
    .A2(net127),
    .B1(_08671_),
    .B2(_08672_),
    .Y(_08674_));
 sky130_fd_sc_hd__nor2_1 _17205_ (.A(_08673_),
    .B(_08674_),
    .Y(_08675_));
 sky130_fd_sc_hd__nand2_1 _17206_ (.A(net289),
    .B(net141),
    .Y(_08676_));
 sky130_fd_sc_hd__and4_1 _17207_ (.A(net279),
    .B(net284),
    .C(net151),
    .D(net146),
    .X(_08677_));
 sky130_fd_sc_hd__a22o_1 _17208_ (.A1(net279),
    .A2(net151),
    .B1(net146),
    .B2(net284),
    .X(_08678_));
 sky130_fd_sc_hd__and2b_1 _17209_ (.A_N(_08677_),
    .B(_08678_),
    .X(_08679_));
 sky130_fd_sc_hd__xnor2_1 _17210_ (.A(_08676_),
    .B(_08679_),
    .Y(_08680_));
 sky130_fd_sc_hd__and2_1 _17211_ (.A(_08044_),
    .B(_08046_),
    .X(_08681_));
 sky130_fd_sc_hd__and2b_1 _17212_ (.A_N(_08681_),
    .B(_08680_),
    .X(_08682_));
 sky130_fd_sc_hd__xnor2_1 _17213_ (.A(_08680_),
    .B(_08681_),
    .Y(_08683_));
 sky130_fd_sc_hd__and2_1 _17214_ (.A(_08675_),
    .B(_08683_),
    .X(_08684_));
 sky130_fd_sc_hd__xnor2_1 _17215_ (.A(_08675_),
    .B(_08683_),
    .Y(_08685_));
 sky130_fd_sc_hd__a21o_1 _17216_ (.A1(_08067_),
    .A2(_08069_),
    .B1(_08685_),
    .X(_08686_));
 sky130_fd_sc_hd__nand3_1 _17217_ (.A(_08067_),
    .B(_08069_),
    .C(_08685_),
    .Y(_08687_));
 sky130_fd_sc_hd__and3_1 _17218_ (.A(_08669_),
    .B(_08686_),
    .C(_08687_),
    .X(_08688_));
 sky130_fd_sc_hd__nand3_1 _17219_ (.A(_08669_),
    .B(_08686_),
    .C(_08687_),
    .Y(_08689_));
 sky130_fd_sc_hd__a21oi_2 _17220_ (.A1(_08686_),
    .A2(_08687_),
    .B1(_08669_),
    .Y(_08690_));
 sky130_fd_sc_hd__a31o_1 _17221_ (.A1(net155),
    .A2(net279),
    .A3(_08064_),
    .B1(_08063_),
    .X(_08691_));
 sky130_fd_sc_hd__o21ba_1 _17222_ (.A1(_08071_),
    .A2(_08072_),
    .B1_N(_08073_),
    .X(_08692_));
 sky130_fd_sc_hd__nand2_1 _17223_ (.A(net273),
    .B(net156),
    .Y(_08693_));
 sky130_fd_sc_hd__and4_1 _17224_ (.A(net263),
    .B(net272),
    .C(net167),
    .D(net164),
    .X(_08694_));
 sky130_fd_sc_hd__a22o_1 _17225_ (.A1(net263),
    .A2(net168),
    .B1(net164),
    .B2(net272),
    .X(_08695_));
 sky130_fd_sc_hd__and2b_1 _17226_ (.A_N(_08694_),
    .B(_08695_),
    .X(_08696_));
 sky130_fd_sc_hd__xnor2_2 _17227_ (.A(_08693_),
    .B(_08696_),
    .Y(_08697_));
 sky130_fd_sc_hd__nand2b_1 _17228_ (.A_N(_08692_),
    .B(_08697_),
    .Y(_08698_));
 sky130_fd_sc_hd__xnor2_2 _17229_ (.A(_08692_),
    .B(_08697_),
    .Y(_08699_));
 sky130_fd_sc_hd__nand2_1 _17230_ (.A(_08691_),
    .B(_08699_),
    .Y(_08700_));
 sky130_fd_sc_hd__xor2_2 _17231_ (.A(_08691_),
    .B(_08699_),
    .X(_08701_));
 sky130_fd_sc_hd__nand2_1 _17232_ (.A(net258),
    .B(net175),
    .Y(_08702_));
 sky130_fd_sc_hd__a22oi_2 _17233_ (.A1(net252),
    .A2(net185),
    .B1(net180),
    .B2(net257),
    .Y(_08703_));
 sky130_fd_sc_hd__and4_1 _17234_ (.A(net252),
    .B(net257),
    .C(net185),
    .D(net180),
    .X(_08704_));
 sky130_fd_sc_hd__nor2_1 _17235_ (.A(_08703_),
    .B(_08704_),
    .Y(_08705_));
 sky130_fd_sc_hd__xnor2_2 _17236_ (.A(_08702_),
    .B(_08705_),
    .Y(_08706_));
 sky130_fd_sc_hd__and2_1 _17237_ (.A(net630),
    .B(net187),
    .X(_08707_));
 sky130_fd_sc_hd__nand4_1 _17238_ (.A(net625),
    .B(net247),
    .C(net192),
    .D(net240),
    .Y(_08708_));
 sky130_fd_sc_hd__a22o_1 _17239_ (.A1(net247),
    .A2(net192),
    .B1(net240),
    .B2(net625),
    .X(_08709_));
 sky130_fd_sc_hd__nand3_1 _17240_ (.A(_08707_),
    .B(_08708_),
    .C(_08709_),
    .Y(_08710_));
 sky130_fd_sc_hd__a21o_1 _17241_ (.A1(_08708_),
    .A2(_08709_),
    .B1(_08707_),
    .X(_08711_));
 sky130_fd_sc_hd__a21bo_1 _17242_ (.A1(_08076_),
    .A2(_08078_),
    .B1_N(_08077_),
    .X(_08712_));
 sky130_fd_sc_hd__nand3_1 _17243_ (.A(_08710_),
    .B(_08711_),
    .C(_08712_),
    .Y(_08713_));
 sky130_fd_sc_hd__a21o_1 _17244_ (.A1(_08710_),
    .A2(_08711_),
    .B1(_08712_),
    .X(_08714_));
 sky130_fd_sc_hd__nand3_2 _17245_ (.A(_08706_),
    .B(_08713_),
    .C(_08714_),
    .Y(_08715_));
 sky130_fd_sc_hd__a21o_1 _17246_ (.A1(_08713_),
    .A2(_08714_),
    .B1(_08706_),
    .X(_08716_));
 sky130_fd_sc_hd__a21bo_1 _17247_ (.A1(_08075_),
    .A2(_08087_),
    .B1_N(_08086_),
    .X(_08717_));
 sky130_fd_sc_hd__nand3_4 _17248_ (.A(_08715_),
    .B(_08716_),
    .C(_08717_),
    .Y(_08718_));
 sky130_fd_sc_hd__a21o_1 _17249_ (.A1(_08715_),
    .A2(_08716_),
    .B1(_08717_),
    .X(_08719_));
 sky130_fd_sc_hd__and3_1 _17250_ (.A(_08701_),
    .B(_08718_),
    .C(_08719_),
    .X(_08720_));
 sky130_fd_sc_hd__nand3_2 _17251_ (.A(_08701_),
    .B(_08718_),
    .C(_08719_),
    .Y(_08721_));
 sky130_fd_sc_hd__a21oi_2 _17252_ (.A1(_08718_),
    .A2(_08719_),
    .B1(_08701_),
    .Y(_08722_));
 sky130_fd_sc_hd__a211oi_4 _17253_ (.A1(_08102_),
    .A2(_08105_),
    .B1(_08720_),
    .C1(_08722_),
    .Y(_08723_));
 sky130_fd_sc_hd__o211a_1 _17254_ (.A1(_08720_),
    .A2(_08722_),
    .B1(_08102_),
    .C1(_08105_),
    .X(_08724_));
 sky130_fd_sc_hd__nor4_1 _17255_ (.A(_08688_),
    .B(_08690_),
    .C(_08723_),
    .D(_08724_),
    .Y(_08725_));
 sky130_fd_sc_hd__or4_2 _17256_ (.A(_08688_),
    .B(_08690_),
    .C(_08723_),
    .D(_08724_),
    .X(_08726_));
 sky130_fd_sc_hd__o22ai_4 _17257_ (.A1(_08688_),
    .A2(_08690_),
    .B1(_08723_),
    .B2(_08724_),
    .Y(_08727_));
 sky130_fd_sc_hd__o211ai_4 _17258_ (.A1(_08125_),
    .A2(_08127_),
    .B1(_08726_),
    .C1(_08727_),
    .Y(_08728_));
 sky130_fd_sc_hd__a211o_1 _17259_ (.A1(_08726_),
    .A2(_08727_),
    .B1(_08125_),
    .C1(_08127_),
    .X(_08729_));
 sky130_fd_sc_hd__nand3_2 _17260_ (.A(_08668_),
    .B(_08728_),
    .C(_08729_),
    .Y(_08730_));
 sky130_fd_sc_hd__a21o_1 _17261_ (.A1(_08728_),
    .A2(_08729_),
    .B1(_08668_),
    .X(_08731_));
 sky130_fd_sc_hd__o211a_1 _17262_ (.A1(_08155_),
    .A2(_08157_),
    .B1(_08730_),
    .C1(_08731_),
    .X(_08732_));
 sky130_fd_sc_hd__a211oi_2 _17263_ (.A1(_08730_),
    .A2(_08731_),
    .B1(_08155_),
    .C1(_08157_),
    .Y(_08733_));
 sky130_fd_sc_hd__nor2_2 _17264_ (.A(_08732_),
    .B(_08733_),
    .Y(_08734_));
 sky130_fd_sc_hd__xnor2_4 _17265_ (.A(_08647_),
    .B(_08734_),
    .Y(_08735_));
 sky130_fd_sc_hd__nand2_1 _17266_ (.A(_08646_),
    .B(_08735_),
    .Y(_08736_));
 sky130_fd_sc_hd__xnor2_4 _17267_ (.A(_08646_),
    .B(_08735_),
    .Y(_08737_));
 sky130_fd_sc_hd__o21a_1 _17268_ (.A1(_08263_),
    .A2(_08327_),
    .B1(_08262_),
    .X(_08738_));
 sky130_fd_sc_hd__xnor2_4 _17269_ (.A(_08737_),
    .B(_08738_),
    .Y(_08739_));
 sky130_fd_sc_hd__o22a_4 _17270_ (.A1(_08263_),
    .A2(_08383_),
    .B1(_08385_),
    .B2(_08641_),
    .X(_08740_));
 sky130_fd_sc_hd__xnor2_4 _17271_ (.A(_08739_),
    .B(_08740_),
    .Y(_08741_));
 sky130_fd_sc_hd__o22a_1 _17272_ (.A1(net43),
    .A2(_03893_),
    .B1(_08741_),
    .B2(_03049_),
    .X(_08742_));
 sky130_fd_sc_hd__a21bo_1 _17273_ (.A1(net778),
    .A2(net7),
    .B1_N(_08742_),
    .X(_08743_));
 sky130_fd_sc_hd__mux2_1 _17274_ (.A0(net869),
    .A1(_08743_),
    .S(net3),
    .X(_00300_));
 sky130_fd_sc_hd__a31oi_4 _17275_ (.A1(_07972_),
    .A2(_08019_),
    .A3(_08666_),
    .B1(_08665_),
    .Y(_08744_));
 sky130_fd_sc_hd__a22o_1 _17276_ (.A1(net319),
    .A2(net107),
    .B1(net102),
    .B2(net323),
    .X(_08745_));
 sky130_fd_sc_hd__and4_1 _17277_ (.A(net319),
    .B(net323),
    .C(net107),
    .D(net102),
    .X(_08746_));
 sky130_fd_sc_hd__inv_2 _17278_ (.A(_08746_),
    .Y(_08747_));
 sky130_fd_sc_hd__and2_1 _17279_ (.A(_08745_),
    .B(_08747_),
    .X(_08748_));
 sky130_fd_sc_hd__a41o_1 _17280_ (.A1(net310),
    .A2(net315),
    .A3(net122),
    .A4(net117),
    .B1(_08653_),
    .X(_08749_));
 sky130_fd_sc_hd__or2_1 _17281_ (.A(_08670_),
    .B(_08673_),
    .X(_08750_));
 sky130_fd_sc_hd__nand2_1 _17282_ (.A(net315),
    .B(net114),
    .Y(_08751_));
 sky130_fd_sc_hd__and4_1 _17283_ (.A(net305),
    .B(net310),
    .C(net122),
    .D(net117),
    .X(_08752_));
 sky130_fd_sc_hd__a22o_1 _17284_ (.A1(net305),
    .A2(net122),
    .B1(net117),
    .B2(net310),
    .X(_08753_));
 sky130_fd_sc_hd__and2b_1 _17285_ (.A_N(_08752_),
    .B(_08753_),
    .X(_08754_));
 sky130_fd_sc_hd__xnor2_1 _17286_ (.A(_08751_),
    .B(_08754_),
    .Y(_08755_));
 sky130_fd_sc_hd__nand2_1 _17287_ (.A(_08750_),
    .B(_08755_),
    .Y(_08756_));
 sky130_fd_sc_hd__xor2_1 _17288_ (.A(_08750_),
    .B(_08755_),
    .X(_08757_));
 sky130_fd_sc_hd__nand2_1 _17289_ (.A(_08749_),
    .B(_08757_),
    .Y(_08758_));
 sky130_fd_sc_hd__xnor2_1 _17290_ (.A(_08749_),
    .B(_08757_),
    .Y(_08759_));
 sky130_fd_sc_hd__a21bo_1 _17291_ (.A1(_08649_),
    .A2(_08657_),
    .B1_N(_08656_),
    .X(_08760_));
 sky130_fd_sc_hd__and2b_1 _17292_ (.A_N(_08759_),
    .B(_08760_),
    .X(_08761_));
 sky130_fd_sc_hd__xnor2_1 _17293_ (.A(_08759_),
    .B(_08760_),
    .Y(_08762_));
 sky130_fd_sc_hd__xnor2_1 _17294_ (.A(_08748_),
    .B(_08762_),
    .Y(_08763_));
 sky130_fd_sc_hd__a21o_1 _17295_ (.A1(_08686_),
    .A2(_08689_),
    .B1(_08763_),
    .X(_08764_));
 sky130_fd_sc_hd__inv_2 _17296_ (.A(_08764_),
    .Y(_08765_));
 sky130_fd_sc_hd__nand3_1 _17297_ (.A(_08686_),
    .B(_08689_),
    .C(_08763_),
    .Y(_08766_));
 sky130_fd_sc_hd__o211a_1 _17298_ (.A1(_08660_),
    .A2(_08663_),
    .B1(_08764_),
    .C1(_08766_),
    .X(_08767_));
 sky130_fd_sc_hd__a211oi_2 _17299_ (.A1(_08764_),
    .A2(_08766_),
    .B1(_08660_),
    .C1(_08663_),
    .Y(_08768_));
 sky130_fd_sc_hd__and4_1 _17300_ (.A(net289),
    .B(net295),
    .C(net136),
    .D(net131),
    .X(_08769_));
 sky130_fd_sc_hd__inv_2 _17301_ (.A(_08769_),
    .Y(_08770_));
 sky130_fd_sc_hd__a22o_1 _17302_ (.A1(net289),
    .A2(net136),
    .B1(net131),
    .B2(net295),
    .X(_08771_));
 sky130_fd_sc_hd__and4b_1 _17303_ (.A_N(_08769_),
    .B(_08771_),
    .C(net300),
    .D(net127),
    .X(_08772_));
 sky130_fd_sc_hd__a22oi_1 _17304_ (.A1(net300),
    .A2(net127),
    .B1(_08770_),
    .B2(_08771_),
    .Y(_08773_));
 sky130_fd_sc_hd__nor2_1 _17305_ (.A(_08772_),
    .B(_08773_),
    .Y(_08774_));
 sky130_fd_sc_hd__nand2_1 _17306_ (.A(net284),
    .B(net142),
    .Y(_08775_));
 sky130_fd_sc_hd__and4_1 _17307_ (.A(net274),
    .B(net279),
    .C(net151),
    .D(net146),
    .X(_08776_));
 sky130_fd_sc_hd__a22o_1 _17308_ (.A1(net274),
    .A2(net151),
    .B1(net146),
    .B2(net279),
    .X(_08777_));
 sky130_fd_sc_hd__and2b_1 _17309_ (.A_N(_08776_),
    .B(_08777_),
    .X(_08778_));
 sky130_fd_sc_hd__xnor2_1 _17310_ (.A(_08775_),
    .B(_08778_),
    .Y(_08779_));
 sky130_fd_sc_hd__a31o_1 _17311_ (.A1(net289),
    .A2(net141),
    .A3(_08678_),
    .B1(_08677_),
    .X(_08780_));
 sky130_fd_sc_hd__and2_2 _17312_ (.A(_08779_),
    .B(_08780_),
    .X(_08781_));
 sky130_fd_sc_hd__xor2_1 _17313_ (.A(_08779_),
    .B(_08780_),
    .X(_08782_));
 sky130_fd_sc_hd__and2_2 _17314_ (.A(_08774_),
    .B(_08782_),
    .X(_08783_));
 sky130_fd_sc_hd__xnor2_1 _17315_ (.A(_08774_),
    .B(_08782_),
    .Y(_08784_));
 sky130_fd_sc_hd__a21o_2 _17316_ (.A1(_08698_),
    .A2(_08700_),
    .B1(_08784_),
    .X(_08785_));
 sky130_fd_sc_hd__nand3_2 _17317_ (.A(_08698_),
    .B(_08700_),
    .C(_08784_),
    .Y(_08786_));
 sky130_fd_sc_hd__o211a_1 _17318_ (.A1(_08682_),
    .A2(_08684_),
    .B1(_08785_),
    .C1(_08786_),
    .X(_08787_));
 sky130_fd_sc_hd__o211ai_2 _17319_ (.A1(_08682_),
    .A2(_08684_),
    .B1(_08785_),
    .C1(_08786_),
    .Y(_08788_));
 sky130_fd_sc_hd__a211oi_2 _17320_ (.A1(_08785_),
    .A2(_08786_),
    .B1(_08682_),
    .C1(_08684_),
    .Y(_08789_));
 sky130_fd_sc_hd__a31o_1 _17321_ (.A1(net273),
    .A2(net158),
    .A3(_08695_),
    .B1(_08694_),
    .X(_08790_));
 sky130_fd_sc_hd__o21ba_1 _17322_ (.A1(_08702_),
    .A2(_08703_),
    .B1_N(_08704_),
    .X(_08791_));
 sky130_fd_sc_hd__nand2_1 _17323_ (.A(net272),
    .B(net156),
    .Y(_08792_));
 sky130_fd_sc_hd__and4_1 _17324_ (.A(net258),
    .B(net263),
    .C(net168),
    .D(net164),
    .X(_08793_));
 sky130_fd_sc_hd__a22o_1 _17325_ (.A1(net258),
    .A2(net168),
    .B1(net164),
    .B2(net263),
    .X(_08794_));
 sky130_fd_sc_hd__and2b_1 _17326_ (.A_N(_08793_),
    .B(_08794_),
    .X(_08795_));
 sky130_fd_sc_hd__xnor2_2 _17327_ (.A(_08792_),
    .B(_08795_),
    .Y(_08796_));
 sky130_fd_sc_hd__nand2b_2 _17328_ (.A_N(_08791_),
    .B(_08796_),
    .Y(_08797_));
 sky130_fd_sc_hd__xnor2_2 _17329_ (.A(_08791_),
    .B(_08796_),
    .Y(_08798_));
 sky130_fd_sc_hd__nand2_2 _17330_ (.A(_08790_),
    .B(_08798_),
    .Y(_08799_));
 sky130_fd_sc_hd__xor2_2 _17331_ (.A(_08790_),
    .B(_08798_),
    .X(_08800_));
 sky130_fd_sc_hd__nand2_1 _17332_ (.A(net257),
    .B(net175),
    .Y(_08801_));
 sky130_fd_sc_hd__a22oi_2 _17333_ (.A1(net630),
    .A2(net185),
    .B1(net180),
    .B2(net252),
    .Y(_08802_));
 sky130_fd_sc_hd__and4_1 _17334_ (.A(net630),
    .B(net252),
    .C(net185),
    .D(net180),
    .X(_08803_));
 sky130_fd_sc_hd__nor2_1 _17335_ (.A(_08802_),
    .B(_08803_),
    .Y(_08804_));
 sky130_fd_sc_hd__xnor2_2 _17336_ (.A(_08801_),
    .B(_08804_),
    .Y(_08805_));
 sky130_fd_sc_hd__and2_1 _17337_ (.A(net247),
    .B(net187),
    .X(_08806_));
 sky130_fd_sc_hd__nand4_1 _17338_ (.A(net625),
    .B(net192),
    .C(net240),
    .D(net235),
    .Y(_08807_));
 sky130_fd_sc_hd__a22o_1 _17339_ (.A1(net192),
    .A2(net240),
    .B1(net235),
    .B2(net625),
    .X(_08808_));
 sky130_fd_sc_hd__nand3_1 _17340_ (.A(_08806_),
    .B(_08807_),
    .C(_08808_),
    .Y(_08809_));
 sky130_fd_sc_hd__a21o_1 _17341_ (.A1(_08807_),
    .A2(_08808_),
    .B1(_08806_),
    .X(_08810_));
 sky130_fd_sc_hd__a21bo_1 _17342_ (.A1(_08707_),
    .A2(_08709_),
    .B1_N(_08708_),
    .X(_08811_));
 sky130_fd_sc_hd__nand3_1 _17343_ (.A(_08809_),
    .B(_08810_),
    .C(_08811_),
    .Y(_08812_));
 sky130_fd_sc_hd__a21o_1 _17344_ (.A1(_08809_),
    .A2(_08810_),
    .B1(_08811_),
    .X(_08813_));
 sky130_fd_sc_hd__nand3_2 _17345_ (.A(_08805_),
    .B(_08812_),
    .C(_08813_),
    .Y(_08814_));
 sky130_fd_sc_hd__a21o_1 _17346_ (.A1(_08812_),
    .A2(_08813_),
    .B1(_08805_),
    .X(_08815_));
 sky130_fd_sc_hd__a21bo_1 _17347_ (.A1(_08706_),
    .A2(_08714_),
    .B1_N(_08713_),
    .X(_08816_));
 sky130_fd_sc_hd__nand3_4 _17348_ (.A(_08814_),
    .B(_08815_),
    .C(_08816_),
    .Y(_08817_));
 sky130_fd_sc_hd__a21o_1 _17349_ (.A1(_08814_),
    .A2(_08815_),
    .B1(_08816_),
    .X(_08818_));
 sky130_fd_sc_hd__and3_1 _17350_ (.A(_08800_),
    .B(_08817_),
    .C(_08818_),
    .X(_08819_));
 sky130_fd_sc_hd__nand3_2 _17351_ (.A(_08800_),
    .B(_08817_),
    .C(_08818_),
    .Y(_08820_));
 sky130_fd_sc_hd__a21oi_2 _17352_ (.A1(_08817_),
    .A2(_08818_),
    .B1(_08800_),
    .Y(_08821_));
 sky130_fd_sc_hd__a211oi_4 _17353_ (.A1(_08718_),
    .A2(_08721_),
    .B1(_08819_),
    .C1(_08821_),
    .Y(_08822_));
 sky130_fd_sc_hd__o211a_1 _17354_ (.A1(_08819_),
    .A2(_08821_),
    .B1(_08718_),
    .C1(_08721_),
    .X(_08823_));
 sky130_fd_sc_hd__nor4_2 _17355_ (.A(_08787_),
    .B(_08789_),
    .C(_08822_),
    .D(_08823_),
    .Y(_08824_));
 sky130_fd_sc_hd__or4_1 _17356_ (.A(_08787_),
    .B(_08789_),
    .C(_08822_),
    .D(_08823_),
    .X(_08825_));
 sky130_fd_sc_hd__o22ai_1 _17357_ (.A1(_08787_),
    .A2(_08789_),
    .B1(_08822_),
    .B2(_08823_),
    .Y(_08826_));
 sky130_fd_sc_hd__o211a_1 _17358_ (.A1(_08723_),
    .A2(_08725_),
    .B1(_08825_),
    .C1(_08826_),
    .X(_08827_));
 sky130_fd_sc_hd__a211oi_1 _17359_ (.A1(_08825_),
    .A2(_08826_),
    .B1(_08723_),
    .C1(_08725_),
    .Y(_08828_));
 sky130_fd_sc_hd__nor4_2 _17360_ (.A(_08767_),
    .B(_08768_),
    .C(_08827_),
    .D(_08828_),
    .Y(_08829_));
 sky130_fd_sc_hd__o22a_1 _17361_ (.A1(_08767_),
    .A2(_08768_),
    .B1(_08827_),
    .B2(_08828_),
    .X(_08830_));
 sky130_fd_sc_hd__nor2_2 _17362_ (.A(_08829_),
    .B(_08830_),
    .Y(_08831_));
 sky130_fd_sc_hd__nand2_2 _17363_ (.A(_08728_),
    .B(_08730_),
    .Y(_08832_));
 sky130_fd_sc_hd__nand2_1 _17364_ (.A(_08831_),
    .B(_08832_),
    .Y(_08833_));
 sky130_fd_sc_hd__xnor2_4 _17365_ (.A(_08831_),
    .B(_08832_),
    .Y(_08834_));
 sky130_fd_sc_hd__xor2_4 _17366_ (.A(_08744_),
    .B(_08834_),
    .X(_08835_));
 sky130_fd_sc_hd__o21bai_4 _17367_ (.A1(_08647_),
    .A2(_08733_),
    .B1_N(_08732_),
    .Y(_08836_));
 sky130_fd_sc_hd__and2_1 _17368_ (.A(_08835_),
    .B(_08836_),
    .X(_08837_));
 sky130_fd_sc_hd__xnor2_4 _17369_ (.A(_08835_),
    .B(_08836_),
    .Y(_08838_));
 sky130_fd_sc_hd__o21a_1 _17370_ (.A1(_08262_),
    .A2(_08737_),
    .B1(_08736_),
    .X(_08839_));
 sky130_fd_sc_hd__xnor2_4 _17371_ (.A(_08838_),
    .B(_08839_),
    .Y(_08840_));
 sky130_fd_sc_hd__or3_1 _17372_ (.A(_08263_),
    .B(_08327_),
    .C(_08737_),
    .X(_08841_));
 sky130_fd_sc_hd__o21ai_2 _17373_ (.A1(_08739_),
    .A2(_08740_),
    .B1(_08841_),
    .Y(_08842_));
 sky130_fd_sc_hd__xor2_4 _17374_ (.A(_08840_),
    .B(_08842_),
    .X(_08843_));
 sky130_fd_sc_hd__o22a_1 _17375_ (.A1(net43),
    .A2(_03993_),
    .B1(_08843_),
    .B2(_03049_),
    .X(_08844_));
 sky130_fd_sc_hd__a21bo_1 _17376_ (.A1(\temp[2] ),
    .A2(net7),
    .B1_N(_08844_),
    .X(_08845_));
 sky130_fd_sc_hd__mux2_1 _17377_ (.A0(net780),
    .A1(_08845_),
    .S(net3),
    .X(_00301_));
 sky130_fd_sc_hd__nor2_1 _17378_ (.A(net43),
    .B(_04100_),
    .Y(_08846_));
 sky130_fd_sc_hd__or3_1 _17379_ (.A(_08262_),
    .B(_08737_),
    .C(_08838_),
    .X(_08847_));
 sky130_fd_sc_hd__or2_1 _17380_ (.A(_08840_),
    .B(_08841_),
    .X(_08848_));
 sky130_fd_sc_hd__or3_1 _17381_ (.A(_08739_),
    .B(_08740_),
    .C(_08840_),
    .X(_08849_));
 sky130_fd_sc_hd__nor2_2 _17382_ (.A(_08765_),
    .B(_08767_),
    .Y(_08850_));
 sky130_fd_sc_hd__a21oi_1 _17383_ (.A1(_08748_),
    .A2(_08762_),
    .B1(_08761_),
    .Y(_08851_));
 sky130_fd_sc_hd__nand4_1 _17384_ (.A(\mul1.a[2] ),
    .B(net320),
    .C(net107),
    .D(net102),
    .Y(_08852_));
 sky130_fd_sc_hd__a22o_1 _17385_ (.A1(net315),
    .A2(net107),
    .B1(net102),
    .B2(net319),
    .X(_08853_));
 sky130_fd_sc_hd__nand2_1 _17386_ (.A(_08852_),
    .B(_08853_),
    .Y(_08854_));
 sky130_fd_sc_hd__nand2_1 _17387_ (.A(net323),
    .B(net98),
    .Y(_08855_));
 sky130_fd_sc_hd__xnor2_1 _17388_ (.A(_08854_),
    .B(_08855_),
    .Y(_08856_));
 sky130_fd_sc_hd__nor2_1 _17389_ (.A(_08747_),
    .B(_08856_),
    .Y(_08857_));
 sky130_fd_sc_hd__and2_1 _17390_ (.A(_08747_),
    .B(_08856_),
    .X(_08858_));
 sky130_fd_sc_hd__or2_1 _17391_ (.A(_08857_),
    .B(_08858_),
    .X(_08859_));
 sky130_fd_sc_hd__a31o_1 _17392_ (.A1(net315),
    .A2(net114),
    .A3(_08753_),
    .B1(_08752_),
    .X(_08860_));
 sky130_fd_sc_hd__or2_1 _17393_ (.A(_08769_),
    .B(_08772_),
    .X(_08861_));
 sky130_fd_sc_hd__nand2_1 _17394_ (.A(net310),
    .B(net114),
    .Y(_08862_));
 sky130_fd_sc_hd__and4_1 _17395_ (.A(net300),
    .B(net305),
    .C(net122),
    .D(net117),
    .X(_08863_));
 sky130_fd_sc_hd__a22o_1 _17396_ (.A1(net300),
    .A2(net122),
    .B1(net117),
    .B2(net305),
    .X(_08864_));
 sky130_fd_sc_hd__and2b_1 _17397_ (.A_N(_08863_),
    .B(_08864_),
    .X(_08865_));
 sky130_fd_sc_hd__xnor2_2 _17398_ (.A(_08862_),
    .B(_08865_),
    .Y(_08866_));
 sky130_fd_sc_hd__nand2_1 _17399_ (.A(_08861_),
    .B(_08866_),
    .Y(_08867_));
 sky130_fd_sc_hd__xor2_2 _17400_ (.A(_08861_),
    .B(_08866_),
    .X(_08868_));
 sky130_fd_sc_hd__nand2_1 _17401_ (.A(_08860_),
    .B(_08868_),
    .Y(_08869_));
 sky130_fd_sc_hd__xnor2_2 _17402_ (.A(_08860_),
    .B(_08868_),
    .Y(_08870_));
 sky130_fd_sc_hd__a21oi_4 _17403_ (.A1(_08756_),
    .A2(_08758_),
    .B1(_08870_),
    .Y(_08871_));
 sky130_fd_sc_hd__and3_1 _17404_ (.A(_08756_),
    .B(_08758_),
    .C(_08870_),
    .X(_08872_));
 sky130_fd_sc_hd__nor3_2 _17405_ (.A(_08859_),
    .B(_08871_),
    .C(_08872_),
    .Y(_08873_));
 sky130_fd_sc_hd__o21a_1 _17406_ (.A1(_08871_),
    .A2(_08872_),
    .B1(_08859_),
    .X(_08874_));
 sky130_fd_sc_hd__a211oi_2 _17407_ (.A1(_08785_),
    .A2(_08788_),
    .B1(_08873_),
    .C1(_08874_),
    .Y(_08875_));
 sky130_fd_sc_hd__o211a_1 _17408_ (.A1(_08873_),
    .A2(_08874_),
    .B1(_08785_),
    .C1(_08788_),
    .X(_08876_));
 sky130_fd_sc_hd__nor3_1 _17409_ (.A(_08851_),
    .B(_08875_),
    .C(_08876_),
    .Y(_08877_));
 sky130_fd_sc_hd__o21a_1 _17410_ (.A1(_08875_),
    .A2(_08876_),
    .B1(_08851_),
    .X(_08878_));
 sky130_fd_sc_hd__nand4_2 _17411_ (.A(net284),
    .B(net289),
    .C(net137),
    .D(net132),
    .Y(_08879_));
 sky130_fd_sc_hd__a22o_1 _17412_ (.A1(net284),
    .A2(net137),
    .B1(net132),
    .B2(net289),
    .X(_08880_));
 sky130_fd_sc_hd__nand4_1 _17413_ (.A(net295),
    .B(net128),
    .C(_08879_),
    .D(_08880_),
    .Y(_08881_));
 sky130_fd_sc_hd__a22o_1 _17414_ (.A1(net295),
    .A2(net127),
    .B1(_08879_),
    .B2(_08880_),
    .X(_08882_));
 sky130_fd_sc_hd__and2_1 _17415_ (.A(_08881_),
    .B(_08882_),
    .X(_08883_));
 sky130_fd_sc_hd__nand2_1 _17416_ (.A(net279),
    .B(net142),
    .Y(_08884_));
 sky130_fd_sc_hd__and4_1 _17417_ (.A(net272),
    .B(net274),
    .C(net151),
    .D(net146),
    .X(_08885_));
 sky130_fd_sc_hd__a22o_1 _17418_ (.A1(net272),
    .A2(net151),
    .B1(net146),
    .B2(net274),
    .X(_08886_));
 sky130_fd_sc_hd__and2b_1 _17419_ (.A_N(_08885_),
    .B(_08886_),
    .X(_08887_));
 sky130_fd_sc_hd__xnor2_2 _17420_ (.A(_08884_),
    .B(_08887_),
    .Y(_08888_));
 sky130_fd_sc_hd__a31o_1 _17421_ (.A1(net284),
    .A2(net142),
    .A3(_08777_),
    .B1(_08776_),
    .X(_08889_));
 sky130_fd_sc_hd__and2_2 _17422_ (.A(_08888_),
    .B(_08889_),
    .X(_08890_));
 sky130_fd_sc_hd__xor2_2 _17423_ (.A(_08888_),
    .B(_08889_),
    .X(_08891_));
 sky130_fd_sc_hd__and2_2 _17424_ (.A(_08883_),
    .B(_08891_),
    .X(_08892_));
 sky130_fd_sc_hd__xnor2_2 _17425_ (.A(_08883_),
    .B(_08891_),
    .Y(_08893_));
 sky130_fd_sc_hd__a21o_2 _17426_ (.A1(_08797_),
    .A2(_08799_),
    .B1(_08893_),
    .X(_08894_));
 sky130_fd_sc_hd__nand3_4 _17427_ (.A(_08797_),
    .B(_08799_),
    .C(_08893_),
    .Y(_08895_));
 sky130_fd_sc_hd__o211a_2 _17428_ (.A1(_08781_),
    .A2(_08783_),
    .B1(_08894_),
    .C1(_08895_),
    .X(_08896_));
 sky130_fd_sc_hd__o211ai_4 _17429_ (.A1(_08781_),
    .A2(_08783_),
    .B1(_08894_),
    .C1(_08895_),
    .Y(_08897_));
 sky130_fd_sc_hd__a211oi_4 _17430_ (.A1(_08894_),
    .A2(_08895_),
    .B1(_08781_),
    .C1(_08783_),
    .Y(_08898_));
 sky130_fd_sc_hd__a31o_1 _17431_ (.A1(net272),
    .A2(net156),
    .A3(_08794_),
    .B1(_08793_),
    .X(_08899_));
 sky130_fd_sc_hd__o21ba_1 _17432_ (.A1(_08801_),
    .A2(_08802_),
    .B1_N(_08803_),
    .X(_08900_));
 sky130_fd_sc_hd__nand2_1 _17433_ (.A(net263),
    .B(net156),
    .Y(_08901_));
 sky130_fd_sc_hd__and4_1 _17434_ (.A(net256),
    .B(net258),
    .C(net167),
    .D(net161),
    .X(_08902_));
 sky130_fd_sc_hd__a22o_1 _17435_ (.A1(net256),
    .A2(net167),
    .B1(net161),
    .B2(net258),
    .X(_08903_));
 sky130_fd_sc_hd__and2b_1 _17436_ (.A_N(_08902_),
    .B(_08903_),
    .X(_08904_));
 sky130_fd_sc_hd__xnor2_2 _17437_ (.A(_08901_),
    .B(_08904_),
    .Y(_08905_));
 sky130_fd_sc_hd__nand2b_2 _17438_ (.A_N(_08900_),
    .B(_08905_),
    .Y(_08906_));
 sky130_fd_sc_hd__xnor2_2 _17439_ (.A(_08900_),
    .B(_08905_),
    .Y(_08907_));
 sky130_fd_sc_hd__nand2_2 _17440_ (.A(_08899_),
    .B(_08907_),
    .Y(_08908_));
 sky130_fd_sc_hd__xor2_2 _17441_ (.A(_08899_),
    .B(_08907_),
    .X(_08909_));
 sky130_fd_sc_hd__nand2_1 _17442_ (.A(net251),
    .B(net175),
    .Y(_08910_));
 sky130_fd_sc_hd__and4_1 _17443_ (.A(net247),
    .B(net630),
    .C(net185),
    .D(net180),
    .X(_08911_));
 sky130_fd_sc_hd__a22oi_1 _17444_ (.A1(net247),
    .A2(net183),
    .B1(net180),
    .B2(net630),
    .Y(_08912_));
 sky130_fd_sc_hd__nor2_1 _17445_ (.A(_08911_),
    .B(_08912_),
    .Y(_08913_));
 sky130_fd_sc_hd__xnor2_2 _17446_ (.A(_08910_),
    .B(_08913_),
    .Y(_08914_));
 sky130_fd_sc_hd__and2_1 _17447_ (.A(net187),
    .B(net240),
    .X(_08915_));
 sky130_fd_sc_hd__nand4_1 _17448_ (.A(net625),
    .B(net192),
    .C(net235),
    .D(net232),
    .Y(_08916_));
 sky130_fd_sc_hd__a22o_1 _17449_ (.A1(net192),
    .A2(net235),
    .B1(net232),
    .B2(net625),
    .X(_08917_));
 sky130_fd_sc_hd__nand3_1 _17450_ (.A(_08915_),
    .B(_08916_),
    .C(_08917_),
    .Y(_08918_));
 sky130_fd_sc_hd__a21o_1 _17451_ (.A1(_08916_),
    .A2(_08917_),
    .B1(_08915_),
    .X(_08919_));
 sky130_fd_sc_hd__a21bo_1 _17452_ (.A1(_08806_),
    .A2(_08808_),
    .B1_N(_08807_),
    .X(_08920_));
 sky130_fd_sc_hd__nand3_2 _17453_ (.A(_08918_),
    .B(_08919_),
    .C(_08920_),
    .Y(_08921_));
 sky130_fd_sc_hd__a21o_1 _17454_ (.A1(_08918_),
    .A2(_08919_),
    .B1(_08920_),
    .X(_08922_));
 sky130_fd_sc_hd__nand3_2 _17455_ (.A(_08914_),
    .B(_08921_),
    .C(_08922_),
    .Y(_08923_));
 sky130_fd_sc_hd__a21o_1 _17456_ (.A1(_08921_),
    .A2(_08922_),
    .B1(_08914_),
    .X(_08924_));
 sky130_fd_sc_hd__a21bo_1 _17457_ (.A1(_08805_),
    .A2(_08813_),
    .B1_N(_08812_),
    .X(_08925_));
 sky130_fd_sc_hd__nand3_4 _17458_ (.A(_08923_),
    .B(_08924_),
    .C(_08925_),
    .Y(_08926_));
 sky130_fd_sc_hd__a21o_1 _17459_ (.A1(_08923_),
    .A2(_08924_),
    .B1(_08925_),
    .X(_08927_));
 sky130_fd_sc_hd__and3_1 _17460_ (.A(_08909_),
    .B(_08926_),
    .C(_08927_),
    .X(_08928_));
 sky130_fd_sc_hd__nand3_2 _17461_ (.A(_08909_),
    .B(_08926_),
    .C(_08927_),
    .Y(_08929_));
 sky130_fd_sc_hd__a21oi_2 _17462_ (.A1(_08926_),
    .A2(_08927_),
    .B1(_08909_),
    .Y(_08930_));
 sky130_fd_sc_hd__a211oi_4 _17463_ (.A1(_08817_),
    .A2(_08820_),
    .B1(_08928_),
    .C1(_08930_),
    .Y(_08931_));
 sky130_fd_sc_hd__o211a_1 _17464_ (.A1(_08928_),
    .A2(_08930_),
    .B1(_08817_),
    .C1(_08820_),
    .X(_08932_));
 sky130_fd_sc_hd__nor4_2 _17465_ (.A(_08896_),
    .B(_08898_),
    .C(_08931_),
    .D(_08932_),
    .Y(_08933_));
 sky130_fd_sc_hd__or4_2 _17466_ (.A(_08896_),
    .B(_08898_),
    .C(_08931_),
    .D(_08932_),
    .X(_08934_));
 sky130_fd_sc_hd__o22ai_4 _17467_ (.A1(_08896_),
    .A2(_08898_),
    .B1(_08931_),
    .B2(_08932_),
    .Y(_08935_));
 sky130_fd_sc_hd__o211ai_4 _17468_ (.A1(_08822_),
    .A2(_08824_),
    .B1(_08934_),
    .C1(_08935_),
    .Y(_08936_));
 sky130_fd_sc_hd__a211o_1 _17469_ (.A1(_08934_),
    .A2(_08935_),
    .B1(_08822_),
    .C1(_08824_),
    .X(_08937_));
 sky130_fd_sc_hd__or4bb_4 _17470_ (.A(_08877_),
    .B(_08878_),
    .C_N(_08936_),
    .D_N(_08937_),
    .X(_08938_));
 sky130_fd_sc_hd__a2bb2o_1 _17471_ (.A1_N(_08877_),
    .A2_N(_08878_),
    .B1(_08936_),
    .B2(_08937_),
    .X(_08939_));
 sky130_fd_sc_hd__o211a_1 _17472_ (.A1(_08827_),
    .A2(_08829_),
    .B1(_08938_),
    .C1(_08939_),
    .X(_08940_));
 sky130_fd_sc_hd__a211oi_2 _17473_ (.A1(_08938_),
    .A2(_08939_),
    .B1(_08827_),
    .C1(_08829_),
    .Y(_08941_));
 sky130_fd_sc_hd__nor2_1 _17474_ (.A(_08940_),
    .B(_08941_),
    .Y(_08942_));
 sky130_fd_sc_hd__xnor2_2 _17475_ (.A(_08850_),
    .B(_08942_),
    .Y(_08943_));
 sky130_fd_sc_hd__o21ai_2 _17476_ (.A1(_08744_),
    .A2(_08834_),
    .B1(_08833_),
    .Y(_08944_));
 sky130_fd_sc_hd__nand2_1 _17477_ (.A(_08943_),
    .B(_08944_),
    .Y(_08945_));
 sky130_fd_sc_hd__xor2_2 _17478_ (.A(_08943_),
    .B(_08944_),
    .X(_08946_));
 sky130_fd_sc_hd__nor2_1 _17479_ (.A(_08736_),
    .B(_08838_),
    .Y(_08947_));
 sky130_fd_sc_hd__nor2_1 _17480_ (.A(_08837_),
    .B(_08947_),
    .Y(_08948_));
 sky130_fd_sc_hd__xor2_1 _17481_ (.A(_08946_),
    .B(_08948_),
    .X(_08949_));
 sky130_fd_sc_hd__a31o_2 _17482_ (.A1(_08847_),
    .A2(_08848_),
    .A3(_08849_),
    .B1(_08949_),
    .X(_08950_));
 sky130_fd_sc_hd__nand4_1 _17483_ (.A(_08847_),
    .B(_08848_),
    .C(_08849_),
    .D(_08949_),
    .Y(_08951_));
 sky130_fd_sc_hd__and2_4 _17484_ (.A(_08950_),
    .B(_08951_),
    .X(_08952_));
 sky130_fd_sc_hd__a221o_1 _17485_ (.A1(\temp[3] ),
    .A2(net7),
    .B1(_08952_),
    .B2(net10),
    .C1(_08846_),
    .X(_08953_));
 sky130_fd_sc_hd__mux2_1 _17486_ (.A0(net736),
    .A1(_08953_),
    .S(net3),
    .X(_00302_));
 sky130_fd_sc_hd__nor2_1 _17487_ (.A(_08875_),
    .B(_08877_),
    .Y(_08954_));
 sky130_fd_sc_hd__or3_4 _17488_ (.A(_08747_),
    .B(_08856_),
    .C(_08954_),
    .X(_08955_));
 sky130_fd_sc_hd__xnor2_2 _17489_ (.A(_08857_),
    .B(_08954_),
    .Y(_08956_));
 sky130_fd_sc_hd__and4_1 _17490_ (.A(net310),
    .B(\mul1.a[2] ),
    .C(net107),
    .D(net102),
    .X(_08957_));
 sky130_fd_sc_hd__inv_2 _17491_ (.A(_08957_),
    .Y(_08958_));
 sky130_fd_sc_hd__a22o_1 _17492_ (.A1(net310),
    .A2(net107),
    .B1(net102),
    .B2(\mul1.a[2] ),
    .X(_08959_));
 sky130_fd_sc_hd__and4_1 _17493_ (.A(net320),
    .B(net98),
    .C(_08958_),
    .D(_08959_),
    .X(_08960_));
 sky130_fd_sc_hd__a22oi_1 _17494_ (.A1(net320),
    .A2(net98),
    .B1(_08958_),
    .B2(_08959_),
    .Y(_08961_));
 sky130_fd_sc_hd__or2_1 _17495_ (.A(_08960_),
    .B(_08961_),
    .X(_08962_));
 sky130_fd_sc_hd__o21ai_1 _17496_ (.A1(_08854_),
    .A2(_08855_),
    .B1(_08852_),
    .Y(_08963_));
 sky130_fd_sc_hd__and2b_1 _17497_ (.A_N(_08962_),
    .B(_08963_),
    .X(_08964_));
 sky130_fd_sc_hd__xnor2_1 _17498_ (.A(_08962_),
    .B(_08963_),
    .Y(_08965_));
 sky130_fd_sc_hd__nand2_1 _17499_ (.A(net325),
    .B(net97),
    .Y(_08966_));
 sky130_fd_sc_hd__xnor2_1 _17500_ (.A(_08965_),
    .B(_08966_),
    .Y(_08967_));
 sky130_fd_sc_hd__a31o_1 _17501_ (.A1(net310),
    .A2(net114),
    .A3(_08864_),
    .B1(_08863_),
    .X(_08968_));
 sky130_fd_sc_hd__and4_1 _17502_ (.A(net295),
    .B(net300),
    .C(net123),
    .D(net118),
    .X(_08969_));
 sky130_fd_sc_hd__a22oi_1 _17503_ (.A1(net295),
    .A2(net123),
    .B1(net118),
    .B2(net300),
    .Y(_08970_));
 sky130_fd_sc_hd__and4bb_1 _17504_ (.A_N(_08969_),
    .B_N(_08970_),
    .C(net305),
    .D(net114),
    .X(_08971_));
 sky130_fd_sc_hd__o2bb2a_1 _17505_ (.A1_N(net305),
    .A2_N(net114),
    .B1(_08969_),
    .B2(_08970_),
    .X(_08972_));
 sky130_fd_sc_hd__a211o_1 _17506_ (.A1(_08879_),
    .A2(_08881_),
    .B1(_08971_),
    .C1(_08972_),
    .X(_08973_));
 sky130_fd_sc_hd__o211ai_1 _17507_ (.A1(_08971_),
    .A2(_08972_),
    .B1(_08879_),
    .C1(_08881_),
    .Y(_08974_));
 sky130_fd_sc_hd__and2_1 _17508_ (.A(_08973_),
    .B(_08974_),
    .X(_08975_));
 sky130_fd_sc_hd__nand2_1 _17509_ (.A(_08968_),
    .B(_08975_),
    .Y(_08976_));
 sky130_fd_sc_hd__xnor2_1 _17510_ (.A(_08968_),
    .B(_08975_),
    .Y(_08977_));
 sky130_fd_sc_hd__a21o_2 _17511_ (.A1(_08867_),
    .A2(_08869_),
    .B1(_08977_),
    .X(_08978_));
 sky130_fd_sc_hd__nand3_1 _17512_ (.A(_08867_),
    .B(_08869_),
    .C(_08977_),
    .Y(_08979_));
 sky130_fd_sc_hd__and3_2 _17513_ (.A(_08967_),
    .B(_08978_),
    .C(_08979_),
    .X(_08980_));
 sky130_fd_sc_hd__inv_2 _17514_ (.A(_08980_),
    .Y(_08981_));
 sky130_fd_sc_hd__a21oi_2 _17515_ (.A1(_08978_),
    .A2(_08979_),
    .B1(_08967_),
    .Y(_08982_));
 sky130_fd_sc_hd__a211o_2 _17516_ (.A1(_08894_),
    .A2(_08897_),
    .B1(_08980_),
    .C1(_08982_),
    .X(_08983_));
 sky130_fd_sc_hd__o211ai_4 _17517_ (.A1(_08980_),
    .A2(_08982_),
    .B1(_08894_),
    .C1(_08897_),
    .Y(_08984_));
 sky130_fd_sc_hd__o211ai_4 _17518_ (.A1(_08871_),
    .A2(_08873_),
    .B1(_08983_),
    .C1(_08984_),
    .Y(_08985_));
 sky130_fd_sc_hd__a211o_1 _17519_ (.A1(_08983_),
    .A2(_08984_),
    .B1(_08871_),
    .C1(_08873_),
    .X(_08986_));
 sky130_fd_sc_hd__nand4_2 _17520_ (.A(net279),
    .B(net284),
    .C(net137),
    .D(net131),
    .Y(_08987_));
 sky130_fd_sc_hd__a22o_1 _17521_ (.A1(net279),
    .A2(net136),
    .B1(net131),
    .B2(net284),
    .X(_08988_));
 sky130_fd_sc_hd__nand4_1 _17522_ (.A(net289),
    .B(net127),
    .C(_08987_),
    .D(_08988_),
    .Y(_08989_));
 sky130_fd_sc_hd__a22o_1 _17523_ (.A1(net289),
    .A2(net127),
    .B1(_08987_),
    .B2(_08988_),
    .X(_08990_));
 sky130_fd_sc_hd__and2_1 _17524_ (.A(_08989_),
    .B(_08990_),
    .X(_08991_));
 sky130_fd_sc_hd__nand2_1 _17525_ (.A(net274),
    .B(net142),
    .Y(_08992_));
 sky130_fd_sc_hd__and4_1 _17526_ (.A(\mul1.a[12] ),
    .B(net268),
    .C(net152),
    .D(net147),
    .X(_08993_));
 sky130_fd_sc_hd__a22o_1 _17527_ (.A1(\mul1.a[12] ),
    .A2(net151),
    .B1(net146),
    .B2(net268),
    .X(_08994_));
 sky130_fd_sc_hd__and2b_1 _17528_ (.A_N(_08993_),
    .B(_08994_),
    .X(_08995_));
 sky130_fd_sc_hd__xnor2_2 _17529_ (.A(_08992_),
    .B(_08995_),
    .Y(_08996_));
 sky130_fd_sc_hd__a31o_1 _17530_ (.A1(net279),
    .A2(net141),
    .A3(_08886_),
    .B1(_08885_),
    .X(_08997_));
 sky130_fd_sc_hd__and2_2 _17531_ (.A(_08996_),
    .B(_08997_),
    .X(_08998_));
 sky130_fd_sc_hd__xor2_2 _17532_ (.A(_08996_),
    .B(_08997_),
    .X(_08999_));
 sky130_fd_sc_hd__and2_2 _17533_ (.A(_08991_),
    .B(_08999_),
    .X(_09000_));
 sky130_fd_sc_hd__xnor2_2 _17534_ (.A(_08991_),
    .B(_08999_),
    .Y(_09001_));
 sky130_fd_sc_hd__a21o_2 _17535_ (.A1(_08906_),
    .A2(_08908_),
    .B1(_09001_),
    .X(_09002_));
 sky130_fd_sc_hd__nand3_4 _17536_ (.A(_08906_),
    .B(_08908_),
    .C(_09001_),
    .Y(_09003_));
 sky130_fd_sc_hd__o211a_1 _17537_ (.A1(_08890_),
    .A2(_08892_),
    .B1(_09002_),
    .C1(_09003_),
    .X(_09004_));
 sky130_fd_sc_hd__o211ai_4 _17538_ (.A1(_08890_),
    .A2(_08892_),
    .B1(_09002_),
    .C1(_09003_),
    .Y(_09005_));
 sky130_fd_sc_hd__a211oi_4 _17539_ (.A1(_09002_),
    .A2(_09003_),
    .B1(_08890_),
    .C1(_08892_),
    .Y(_09006_));
 sky130_fd_sc_hd__a31o_1 _17540_ (.A1(\mul1.a[12] ),
    .A2(net156),
    .A3(_08903_),
    .B1(_08902_),
    .X(_09007_));
 sky130_fd_sc_hd__o21ba_1 _17541_ (.A1(_08910_),
    .A2(_08912_),
    .B1_N(_08911_),
    .X(_09008_));
 sky130_fd_sc_hd__nand2_1 _17542_ (.A(\mul1.a[13] ),
    .B(net156),
    .Y(_09009_));
 sky130_fd_sc_hd__and3_1 _17543_ (.A(net251),
    .B(net256),
    .C(net161),
    .X(_09010_));
 sky130_fd_sc_hd__a22o_1 _17544_ (.A1(net251),
    .A2(net167),
    .B1(net161),
    .B2(net256),
    .X(_09011_));
 sky130_fd_sc_hd__a21bo_1 _17545_ (.A1(net167),
    .A2(_09010_),
    .B1_N(_09011_),
    .X(_09012_));
 sky130_fd_sc_hd__xor2_2 _17546_ (.A(_09009_),
    .B(_09012_),
    .X(_09013_));
 sky130_fd_sc_hd__nand2b_2 _17547_ (.A_N(_09008_),
    .B(_09013_),
    .Y(_09014_));
 sky130_fd_sc_hd__xnor2_2 _17548_ (.A(_09008_),
    .B(_09013_),
    .Y(_09015_));
 sky130_fd_sc_hd__nand2_2 _17549_ (.A(_09007_),
    .B(_09015_),
    .Y(_09016_));
 sky130_fd_sc_hd__xor2_2 _17550_ (.A(_09007_),
    .B(_09015_),
    .X(_09017_));
 sky130_fd_sc_hd__a22oi_1 _17551_ (.A1(net247),
    .A2(net178),
    .B1(net240),
    .B2(net183),
    .Y(_09018_));
 sky130_fd_sc_hd__and4_1 _17552_ (.A(net247),
    .B(net183),
    .C(net178),
    .D(net240),
    .X(_09019_));
 sky130_fd_sc_hd__and4bb_1 _17553_ (.A_N(_09018_),
    .B_N(_09019_),
    .C(net630),
    .D(net173),
    .X(_09020_));
 sky130_fd_sc_hd__o2bb2a_1 _17554_ (.A1_N(net630),
    .A2_N(net173),
    .B1(_09018_),
    .B2(_09019_),
    .X(_09021_));
 sky130_fd_sc_hd__nor2_1 _17555_ (.A(_09020_),
    .B(_09021_),
    .Y(_09022_));
 sky130_fd_sc_hd__and2_1 _17556_ (.A(net187),
    .B(net235),
    .X(_09023_));
 sky130_fd_sc_hd__nand4_2 _17557_ (.A(net625),
    .B(net192),
    .C(net232),
    .D(net227),
    .Y(_09024_));
 sky130_fd_sc_hd__a22o_1 _17558_ (.A1(net190),
    .A2(net232),
    .B1(net227),
    .B2(net623),
    .X(_09025_));
 sky130_fd_sc_hd__nand3_1 _17559_ (.A(_09023_),
    .B(_09024_),
    .C(_09025_),
    .Y(_09026_));
 sky130_fd_sc_hd__a21o_1 _17560_ (.A1(_09024_),
    .A2(_09025_),
    .B1(_09023_),
    .X(_09027_));
 sky130_fd_sc_hd__a21bo_1 _17561_ (.A1(_08915_),
    .A2(_08917_),
    .B1_N(_08916_),
    .X(_09028_));
 sky130_fd_sc_hd__nand3_1 _17562_ (.A(_09026_),
    .B(_09027_),
    .C(_09028_),
    .Y(_09029_));
 sky130_fd_sc_hd__a21o_1 _17563_ (.A1(_09026_),
    .A2(_09027_),
    .B1(_09028_),
    .X(_09030_));
 sky130_fd_sc_hd__nand3_2 _17564_ (.A(_09022_),
    .B(_09029_),
    .C(_09030_),
    .Y(_09031_));
 sky130_fd_sc_hd__a21o_1 _17565_ (.A1(_09029_),
    .A2(_09030_),
    .B1(_09022_),
    .X(_09032_));
 sky130_fd_sc_hd__a21bo_1 _17566_ (.A1(_08914_),
    .A2(_08922_),
    .B1_N(_08921_),
    .X(_09033_));
 sky130_fd_sc_hd__nand3_4 _17567_ (.A(_09031_),
    .B(_09032_),
    .C(_09033_),
    .Y(_09034_));
 sky130_fd_sc_hd__a21o_1 _17568_ (.A1(_09031_),
    .A2(_09032_),
    .B1(_09033_),
    .X(_09035_));
 sky130_fd_sc_hd__and3_1 _17569_ (.A(_09017_),
    .B(_09034_),
    .C(_09035_),
    .X(_09036_));
 sky130_fd_sc_hd__nand3_2 _17570_ (.A(_09017_),
    .B(_09034_),
    .C(_09035_),
    .Y(_09037_));
 sky130_fd_sc_hd__a21oi_2 _17571_ (.A1(_09034_),
    .A2(_09035_),
    .B1(_09017_),
    .Y(_09038_));
 sky130_fd_sc_hd__a211oi_4 _17572_ (.A1(_08926_),
    .A2(_08929_),
    .B1(_09036_),
    .C1(_09038_),
    .Y(_09039_));
 sky130_fd_sc_hd__o211a_1 _17573_ (.A1(_09036_),
    .A2(_09038_),
    .B1(_08926_),
    .C1(_08929_),
    .X(_09040_));
 sky130_fd_sc_hd__nor4_2 _17574_ (.A(_09004_),
    .B(_09006_),
    .C(_09039_),
    .D(_09040_),
    .Y(_09041_));
 sky130_fd_sc_hd__or4_2 _17575_ (.A(_09004_),
    .B(_09006_),
    .C(_09039_),
    .D(_09040_),
    .X(_09042_));
 sky130_fd_sc_hd__o22ai_4 _17576_ (.A1(_09004_),
    .A2(_09006_),
    .B1(_09039_),
    .B2(_09040_),
    .Y(_09043_));
 sky130_fd_sc_hd__o211ai_4 _17577_ (.A1(_08931_),
    .A2(_08933_),
    .B1(_09042_),
    .C1(_09043_),
    .Y(_09044_));
 sky130_fd_sc_hd__a211o_1 _17578_ (.A1(_09042_),
    .A2(_09043_),
    .B1(_08931_),
    .C1(_08933_),
    .X(_09045_));
 sky130_fd_sc_hd__and4_1 _17579_ (.A(_08985_),
    .B(_08986_),
    .C(_09044_),
    .D(_09045_),
    .X(_09046_));
 sky130_fd_sc_hd__nand4_1 _17580_ (.A(_08985_),
    .B(_08986_),
    .C(_09044_),
    .D(_09045_),
    .Y(_09047_));
 sky130_fd_sc_hd__a22oi_4 _17581_ (.A1(_08985_),
    .A2(_08986_),
    .B1(_09044_),
    .B2(_09045_),
    .Y(_09048_));
 sky130_fd_sc_hd__a211o_1 _17582_ (.A1(_08936_),
    .A2(_08938_),
    .B1(_09046_),
    .C1(_09048_),
    .X(_09049_));
 sky130_fd_sc_hd__o211ai_4 _17583_ (.A1(_09046_),
    .A2(_09048_),
    .B1(_08936_),
    .C1(_08938_),
    .Y(_09050_));
 sky130_fd_sc_hd__and3_1 _17584_ (.A(_08956_),
    .B(_09049_),
    .C(_09050_),
    .X(_09051_));
 sky130_fd_sc_hd__a21oi_1 _17585_ (.A1(_09049_),
    .A2(_09050_),
    .B1(_08956_),
    .Y(_09052_));
 sky130_fd_sc_hd__nor2_2 _17586_ (.A(_09051_),
    .B(_09052_),
    .Y(_09053_));
 sky130_fd_sc_hd__o21bai_4 _17587_ (.A1(_08850_),
    .A2(_08941_),
    .B1_N(_08940_),
    .Y(_09054_));
 sky130_fd_sc_hd__nand2_1 _17588_ (.A(_09053_),
    .B(_09054_),
    .Y(_09055_));
 sky130_fd_sc_hd__xnor2_4 _17589_ (.A(_09053_),
    .B(_09054_),
    .Y(_09056_));
 sky130_fd_sc_hd__nand2_1 _17590_ (.A(_08837_),
    .B(_08946_),
    .Y(_09057_));
 sky130_fd_sc_hd__a21boi_2 _17591_ (.A1(_08837_),
    .A2(_08946_),
    .B1_N(_08945_),
    .Y(_09058_));
 sky130_fd_sc_hd__xnor2_4 _17592_ (.A(_09056_),
    .B(_09058_),
    .Y(_09059_));
 sky130_fd_sc_hd__nand2_1 _17593_ (.A(_08946_),
    .B(_08947_),
    .Y(_09060_));
 sky130_fd_sc_hd__nand2_2 _17594_ (.A(_08950_),
    .B(_09060_),
    .Y(_09061_));
 sky130_fd_sc_hd__xnor2_4 _17595_ (.A(_09059_),
    .B(_09061_),
    .Y(_09062_));
 sky130_fd_sc_hd__nor2_1 _17596_ (.A(net43),
    .B(_04209_),
    .Y(_09063_));
 sky130_fd_sc_hd__a221o_1 _17597_ (.A1(net706),
    .A2(net7),
    .B1(_09062_),
    .B2(net10),
    .C1(_03056_),
    .X(_09064_));
 sky130_fd_sc_hd__o22a_1 _17598_ (.A1(net861),
    .A2(net3),
    .B1(_09063_),
    .B2(_09064_),
    .X(_00303_));
 sky130_fd_sc_hd__nor2_1 _17599_ (.A(net44),
    .B(_04325_),
    .Y(_09065_));
 sky130_fd_sc_hd__a31oi_2 _17600_ (.A1(net325),
    .A2(net97),
    .A3(_08965_),
    .B1(_08964_),
    .Y(_09066_));
 sky130_fd_sc_hd__a21oi_2 _17601_ (.A1(_08983_),
    .A2(_08985_),
    .B1(_09066_),
    .Y(_09067_));
 sky130_fd_sc_hd__and3_1 _17602_ (.A(_08983_),
    .B(_08985_),
    .C(_09066_),
    .X(_09068_));
 sky130_fd_sc_hd__or2_1 _17603_ (.A(_09067_),
    .B(_09068_),
    .X(_09069_));
 sky130_fd_sc_hd__a22o_1 _17604_ (.A1(net320),
    .A2(net97),
    .B1(net90),
    .B2(net324),
    .X(_09070_));
 sky130_fd_sc_hd__inv_2 _17605_ (.A(_09070_),
    .Y(_09071_));
 sky130_fd_sc_hd__and4_2 _17606_ (.A(net321),
    .B(net324),
    .C(net97),
    .D(net90),
    .X(_09072_));
 sky130_fd_sc_hd__nor2_1 _17607_ (.A(_09071_),
    .B(_09072_),
    .Y(_09073_));
 sky130_fd_sc_hd__and4_1 _17608_ (.A(net307),
    .B(net312),
    .C(net107),
    .D(net102),
    .X(_09074_));
 sky130_fd_sc_hd__inv_2 _17609_ (.A(_09074_),
    .Y(_09075_));
 sky130_fd_sc_hd__a22o_1 _17610_ (.A1(net307),
    .A2(net107),
    .B1(net102),
    .B2(net312),
    .X(_09076_));
 sky130_fd_sc_hd__and4_1 _17611_ (.A(net317),
    .B(net98),
    .C(_09075_),
    .D(_09076_),
    .X(_09077_));
 sky130_fd_sc_hd__a22oi_1 _17612_ (.A1(net317),
    .A2(net98),
    .B1(_09075_),
    .B2(_09076_),
    .Y(_09078_));
 sky130_fd_sc_hd__or2_2 _17613_ (.A(_09077_),
    .B(_09078_),
    .X(_09079_));
 sky130_fd_sc_hd__or2_2 _17614_ (.A(_08957_),
    .B(_08960_),
    .X(_09080_));
 sky130_fd_sc_hd__and2b_1 _17615_ (.A_N(_09079_),
    .B(_09080_),
    .X(_09081_));
 sky130_fd_sc_hd__xor2_4 _17616_ (.A(_09079_),
    .B(_09080_),
    .X(_09082_));
 sky130_fd_sc_hd__xor2_2 _17617_ (.A(_09073_),
    .B(_09082_),
    .X(_09083_));
 sky130_fd_sc_hd__or2_1 _17618_ (.A(_08969_),
    .B(_08971_),
    .X(_09084_));
 sky130_fd_sc_hd__and4_1 _17619_ (.A(net289),
    .B(net295),
    .C(net122),
    .D(net117),
    .X(_09085_));
 sky130_fd_sc_hd__a22oi_1 _17620_ (.A1(net289),
    .A2(net123),
    .B1(net117),
    .B2(net295),
    .Y(_09086_));
 sky130_fd_sc_hd__and4bb_1 _17621_ (.A_N(_09085_),
    .B_N(_09086_),
    .C(net300),
    .D(net114),
    .X(_09087_));
 sky130_fd_sc_hd__o2bb2a_1 _17622_ (.A1_N(net300),
    .A2_N(net114),
    .B1(_09085_),
    .B2(_09086_),
    .X(_09088_));
 sky130_fd_sc_hd__a211o_1 _17623_ (.A1(_08987_),
    .A2(_08989_),
    .B1(_09087_),
    .C1(_09088_),
    .X(_09089_));
 sky130_fd_sc_hd__o211ai_1 _17624_ (.A1(_09087_),
    .A2(_09088_),
    .B1(_08987_),
    .C1(_08989_),
    .Y(_09090_));
 sky130_fd_sc_hd__and2_1 _17625_ (.A(_09089_),
    .B(_09090_),
    .X(_09091_));
 sky130_fd_sc_hd__nand2_1 _17626_ (.A(_09084_),
    .B(_09091_),
    .Y(_09092_));
 sky130_fd_sc_hd__xnor2_2 _17627_ (.A(_09084_),
    .B(_09091_),
    .Y(_09093_));
 sky130_fd_sc_hd__a21oi_4 _17628_ (.A1(_08973_),
    .A2(_08976_),
    .B1(_09093_),
    .Y(_09094_));
 sky130_fd_sc_hd__and3_1 _17629_ (.A(_08973_),
    .B(_08976_),
    .C(_09093_),
    .X(_09095_));
 sky130_fd_sc_hd__nor3_4 _17630_ (.A(_09083_),
    .B(_09094_),
    .C(_09095_),
    .Y(_09096_));
 sky130_fd_sc_hd__o21a_1 _17631_ (.A1(_09094_),
    .A2(_09095_),
    .B1(_09083_),
    .X(_09097_));
 sky130_fd_sc_hd__a211oi_4 _17632_ (.A1(_09002_),
    .A2(_09005_),
    .B1(_09096_),
    .C1(_09097_),
    .Y(_09098_));
 sky130_fd_sc_hd__o211a_1 _17633_ (.A1(_09096_),
    .A2(_09097_),
    .B1(_09002_),
    .C1(_09005_),
    .X(_09099_));
 sky130_fd_sc_hd__a211oi_4 _17634_ (.A1(_08978_),
    .A2(_08981_),
    .B1(_09098_),
    .C1(_09099_),
    .Y(_09100_));
 sky130_fd_sc_hd__o211a_1 _17635_ (.A1(_09098_),
    .A2(_09099_),
    .B1(_08978_),
    .C1(_08981_),
    .X(_09101_));
 sky130_fd_sc_hd__nand2_1 _17636_ (.A(net287),
    .B(net127),
    .Y(_09102_));
 sky130_fd_sc_hd__and3_1 _17637_ (.A(net277),
    .B(net282),
    .C(net133),
    .X(_09103_));
 sky130_fd_sc_hd__a22o_1 _17638_ (.A1(net277),
    .A2(net138),
    .B1(net133),
    .B2(net282),
    .X(_09104_));
 sky130_fd_sc_hd__a21bo_1 _17639_ (.A1(net138),
    .A2(_09103_),
    .B1_N(_09104_),
    .X(_09105_));
 sky130_fd_sc_hd__xor2_2 _17640_ (.A(_09102_),
    .B(_09105_),
    .X(_09106_));
 sky130_fd_sc_hd__nand2_1 _17641_ (.A(net271),
    .B(net144),
    .Y(_09107_));
 sky130_fd_sc_hd__and3_1 _17642_ (.A(net262),
    .B(net267),
    .C(net147),
    .X(_09108_));
 sky130_fd_sc_hd__a22o_1 _17643_ (.A1(net262),
    .A2(net152),
    .B1(net147),
    .B2(net267),
    .X(_09109_));
 sky130_fd_sc_hd__a21bo_1 _17644_ (.A1(net152),
    .A2(_09108_),
    .B1_N(_09109_),
    .X(_09110_));
 sky130_fd_sc_hd__xor2_2 _17645_ (.A(_09107_),
    .B(_09110_),
    .X(_09111_));
 sky130_fd_sc_hd__a31o_1 _17646_ (.A1(net274),
    .A2(net144),
    .A3(_08994_),
    .B1(_08993_),
    .X(_09112_));
 sky130_fd_sc_hd__and2_1 _17647_ (.A(_09111_),
    .B(_09112_),
    .X(_09113_));
 sky130_fd_sc_hd__xor2_2 _17648_ (.A(_09111_),
    .B(_09112_),
    .X(_09114_));
 sky130_fd_sc_hd__and2_1 _17649_ (.A(_09106_),
    .B(_09114_),
    .X(_09115_));
 sky130_fd_sc_hd__xnor2_2 _17650_ (.A(_09106_),
    .B(_09114_),
    .Y(_09116_));
 sky130_fd_sc_hd__a21o_4 _17651_ (.A1(_09014_),
    .A2(_09016_),
    .B1(_09116_),
    .X(_09117_));
 sky130_fd_sc_hd__nand3_4 _17652_ (.A(_09014_),
    .B(_09016_),
    .C(_09116_),
    .Y(_09118_));
 sky130_fd_sc_hd__o211a_1 _17653_ (.A1(_08998_),
    .A2(_09000_),
    .B1(_09117_),
    .C1(_09118_),
    .X(_09119_));
 sky130_fd_sc_hd__o211ai_4 _17654_ (.A1(_08998_),
    .A2(_09000_),
    .B1(_09117_),
    .C1(_09118_),
    .Y(_09120_));
 sky130_fd_sc_hd__a211oi_4 _17655_ (.A1(_09117_),
    .A2(_09118_),
    .B1(_08998_),
    .C1(_09000_),
    .Y(_09121_));
 sky130_fd_sc_hd__a32o_1 _17656_ (.A1(net258),
    .A2(net156),
    .A3(_09011_),
    .B1(_09010_),
    .B2(net167),
    .X(_09122_));
 sky130_fd_sc_hd__nand4_2 _17657_ (.A(net630),
    .B(net251),
    .C(net167),
    .D(net161),
    .Y(_09123_));
 sky130_fd_sc_hd__a22o_1 _17658_ (.A1(net630),
    .A2(net167),
    .B1(net161),
    .B2(net251),
    .X(_09124_));
 sky130_fd_sc_hd__nand4_2 _17659_ (.A(net256),
    .B(net156),
    .C(_09123_),
    .D(_09124_),
    .Y(_09125_));
 sky130_fd_sc_hd__a22o_1 _17660_ (.A1(net256),
    .A2(net156),
    .B1(_09123_),
    .B2(_09124_),
    .X(_09126_));
 sky130_fd_sc_hd__o211a_1 _17661_ (.A1(_09019_),
    .A2(_09020_),
    .B1(_09125_),
    .C1(_09126_),
    .X(_09127_));
 sky130_fd_sc_hd__a211o_1 _17662_ (.A1(_09125_),
    .A2(_09126_),
    .B1(_09019_),
    .C1(_09020_),
    .X(_09128_));
 sky130_fd_sc_hd__nand2b_1 _17663_ (.A_N(_09127_),
    .B(_09128_),
    .Y(_09129_));
 sky130_fd_sc_hd__xnor2_2 _17664_ (.A(_09122_),
    .B(_09129_),
    .Y(_09130_));
 sky130_fd_sc_hd__a22oi_1 _17665_ (.A1(net178),
    .A2(net240),
    .B1(net235),
    .B2(net183),
    .Y(_09131_));
 sky130_fd_sc_hd__and4_1 _17666_ (.A(net185),
    .B(net178),
    .C(net240),
    .D(net235),
    .X(_09132_));
 sky130_fd_sc_hd__and4bb_1 _17667_ (.A_N(_09131_),
    .B_N(_09132_),
    .C(net247),
    .D(net173),
    .X(_09133_));
 sky130_fd_sc_hd__o2bb2a_1 _17668_ (.A1_N(net247),
    .A2_N(net173),
    .B1(_09131_),
    .B2(_09132_),
    .X(_09134_));
 sky130_fd_sc_hd__nor2_1 _17669_ (.A(_09133_),
    .B(_09134_),
    .Y(_09135_));
 sky130_fd_sc_hd__and2_1 _17670_ (.A(\mul1.b[2] ),
    .B(net232),
    .X(_09136_));
 sky130_fd_sc_hd__nand4_1 _17671_ (.A(net623),
    .B(net190),
    .C(net227),
    .D(net221),
    .Y(_09137_));
 sky130_fd_sc_hd__a22o_1 _17672_ (.A1(net190),
    .A2(net227),
    .B1(net221),
    .B2(net623),
    .X(_09138_));
 sky130_fd_sc_hd__nand3_1 _17673_ (.A(_09136_),
    .B(_09137_),
    .C(_09138_),
    .Y(_09139_));
 sky130_fd_sc_hd__a21o_1 _17674_ (.A1(_09137_),
    .A2(_09138_),
    .B1(_09136_),
    .X(_09140_));
 sky130_fd_sc_hd__a21bo_1 _17675_ (.A1(_09023_),
    .A2(_09025_),
    .B1_N(_09024_),
    .X(_09141_));
 sky130_fd_sc_hd__nand3_2 _17676_ (.A(_09139_),
    .B(_09140_),
    .C(_09141_),
    .Y(_09142_));
 sky130_fd_sc_hd__a21o_1 _17677_ (.A1(_09139_),
    .A2(_09140_),
    .B1(_09141_),
    .X(_09143_));
 sky130_fd_sc_hd__nand3_2 _17678_ (.A(_09135_),
    .B(_09142_),
    .C(_09143_),
    .Y(_09144_));
 sky130_fd_sc_hd__a21o_1 _17679_ (.A1(_09142_),
    .A2(_09143_),
    .B1(_09135_),
    .X(_09145_));
 sky130_fd_sc_hd__a21bo_1 _17680_ (.A1(_09022_),
    .A2(_09030_),
    .B1_N(_09029_),
    .X(_09146_));
 sky130_fd_sc_hd__nand3_4 _17681_ (.A(_09144_),
    .B(_09145_),
    .C(_09146_),
    .Y(_09147_));
 sky130_fd_sc_hd__a21o_1 _17682_ (.A1(_09144_),
    .A2(_09145_),
    .B1(_09146_),
    .X(_09148_));
 sky130_fd_sc_hd__and3_1 _17683_ (.A(_09130_),
    .B(_09147_),
    .C(_09148_),
    .X(_09149_));
 sky130_fd_sc_hd__nand3_2 _17684_ (.A(_09130_),
    .B(_09147_),
    .C(_09148_),
    .Y(_09150_));
 sky130_fd_sc_hd__a21oi_2 _17685_ (.A1(_09147_),
    .A2(_09148_),
    .B1(_09130_),
    .Y(_09151_));
 sky130_fd_sc_hd__a211oi_4 _17686_ (.A1(_09034_),
    .A2(_09037_),
    .B1(_09149_),
    .C1(_09151_),
    .Y(_09152_));
 sky130_fd_sc_hd__o211a_1 _17687_ (.A1(_09149_),
    .A2(_09151_),
    .B1(_09034_),
    .C1(_09037_),
    .X(_09153_));
 sky130_fd_sc_hd__nor4_2 _17688_ (.A(_09119_),
    .B(_09121_),
    .C(_09152_),
    .D(_09153_),
    .Y(_09154_));
 sky130_fd_sc_hd__or4_2 _17689_ (.A(_09119_),
    .B(_09121_),
    .C(_09152_),
    .D(_09153_),
    .X(_09155_));
 sky130_fd_sc_hd__o22ai_4 _17690_ (.A1(_09119_),
    .A2(_09121_),
    .B1(_09152_),
    .B2(_09153_),
    .Y(_09156_));
 sky130_fd_sc_hd__o211ai_4 _17691_ (.A1(_09039_),
    .A2(_09041_),
    .B1(_09155_),
    .C1(_09156_),
    .Y(_09157_));
 sky130_fd_sc_hd__a211o_1 _17692_ (.A1(_09155_),
    .A2(_09156_),
    .B1(_09039_),
    .C1(_09041_),
    .X(_09158_));
 sky130_fd_sc_hd__and4bb_1 _17693_ (.A_N(_09100_),
    .B_N(_09101_),
    .C(_09157_),
    .D(_09158_),
    .X(_09159_));
 sky130_fd_sc_hd__or4bb_1 _17694_ (.A(_09100_),
    .B(_09101_),
    .C_N(_09157_),
    .D_N(_09158_),
    .X(_09160_));
 sky130_fd_sc_hd__a2bb2oi_1 _17695_ (.A1_N(_09100_),
    .A2_N(_09101_),
    .B1(_09157_),
    .B2(_09158_),
    .Y(_09161_));
 sky130_fd_sc_hd__a211oi_1 _17696_ (.A1(_09044_),
    .A2(_09047_),
    .B1(_09159_),
    .C1(_09161_),
    .Y(_09162_));
 sky130_fd_sc_hd__o211a_1 _17697_ (.A1(_09159_),
    .A2(_09161_),
    .B1(_09044_),
    .C1(_09047_),
    .X(_09163_));
 sky130_fd_sc_hd__or3_1 _17698_ (.A(_09069_),
    .B(_09162_),
    .C(_09163_),
    .X(_09164_));
 sky130_fd_sc_hd__o21ai_1 _17699_ (.A1(_09162_),
    .A2(_09163_),
    .B1(_09069_),
    .Y(_09165_));
 sky130_fd_sc_hd__nand2_2 _17700_ (.A(_09164_),
    .B(_09165_),
    .Y(_09166_));
 sky130_fd_sc_hd__a21boi_4 _17701_ (.A1(_08956_),
    .A2(_09050_),
    .B1_N(_09049_),
    .Y(_09167_));
 sky130_fd_sc_hd__or2_1 _17702_ (.A(_09166_),
    .B(_09167_),
    .X(_09168_));
 sky130_fd_sc_hd__xnor2_4 _17703_ (.A(_09166_),
    .B(_09167_),
    .Y(_09169_));
 sky130_fd_sc_hd__xnor2_4 _17704_ (.A(_08955_),
    .B(_09169_),
    .Y(_09170_));
 sky130_fd_sc_hd__or2_1 _17705_ (.A(_08945_),
    .B(_09056_),
    .X(_09171_));
 sky130_fd_sc_hd__o21a_1 _17706_ (.A1(_08945_),
    .A2(_09056_),
    .B1(_09055_),
    .X(_09172_));
 sky130_fd_sc_hd__xnor2_4 _17707_ (.A(_09170_),
    .B(_09172_),
    .Y(_09173_));
 sky130_fd_sc_hd__o22a_1 _17708_ (.A1(_09056_),
    .A2(_09057_),
    .B1(_09059_),
    .B2(_09060_),
    .X(_09174_));
 sky130_fd_sc_hd__o21a_2 _17709_ (.A1(_08950_),
    .A2(_09059_),
    .B1(_09174_),
    .X(_09175_));
 sky130_fd_sc_hd__xor2_4 _17710_ (.A(_09173_),
    .B(_09175_),
    .X(_09176_));
 sky130_fd_sc_hd__a221o_1 _17711_ (.A1(net809),
    .A2(net7),
    .B1(_09176_),
    .B2(_03050_),
    .C1(_09065_),
    .X(_09177_));
 sky130_fd_sc_hd__mux2_1 _17712_ (.A0(net875),
    .A1(_09177_),
    .S(net3),
    .X(_00304_));
 sky130_fd_sc_hd__o22a_2 _17713_ (.A1(_09170_),
    .A2(_09171_),
    .B1(_09173_),
    .B2(_09175_),
    .X(_09178_));
 sky130_fd_sc_hd__and2_2 _17714_ (.A(_09072_),
    .B(_09081_),
    .X(_09179_));
 sky130_fd_sc_hd__nor2_1 _17715_ (.A(_09072_),
    .B(_09081_),
    .Y(_09180_));
 sky130_fd_sc_hd__o32ai_4 _17716_ (.A1(_09071_),
    .A2(_09072_),
    .A3(_09082_),
    .B1(_09179_),
    .B2(_09180_),
    .Y(_09181_));
 sky130_fd_sc_hd__o21ai_2 _17717_ (.A1(_09098_),
    .A2(_09100_),
    .B1(_09181_),
    .Y(_09182_));
 sky130_fd_sc_hd__or3_1 _17718_ (.A(_09098_),
    .B(_09100_),
    .C(_09181_),
    .X(_09183_));
 sky130_fd_sc_hd__and2_1 _17719_ (.A(_09182_),
    .B(_09183_),
    .X(_09184_));
 sky130_fd_sc_hd__and4_1 _17720_ (.A(net317),
    .B(net321),
    .C(net94),
    .D(net90),
    .X(_09185_));
 sky130_fd_sc_hd__a22o_1 _17721_ (.A1(net317),
    .A2(net94),
    .B1(net90),
    .B2(net321),
    .X(_09186_));
 sky130_fd_sc_hd__inv_2 _17722_ (.A(_09186_),
    .Y(_09187_));
 sky130_fd_sc_hd__and4b_1 _17723_ (.A_N(_09185_),
    .B(_09186_),
    .C(net324),
    .D(net88),
    .X(_09188_));
 sky130_fd_sc_hd__o2bb2a_1 _17724_ (.A1_N(net324),
    .A2_N(net88),
    .B1(_09185_),
    .B2(_09187_),
    .X(_09189_));
 sky130_fd_sc_hd__or2_1 _17725_ (.A(_09188_),
    .B(_09189_),
    .X(_09190_));
 sky130_fd_sc_hd__and4_1 _17726_ (.A(\mul1.a[5] ),
    .B(net307),
    .C(net111),
    .D(net106),
    .X(_09191_));
 sky130_fd_sc_hd__a22o_1 _17727_ (.A1(\mul1.a[5] ),
    .A2(net111),
    .B1(net106),
    .B2(net307),
    .X(_09192_));
 sky130_fd_sc_hd__inv_2 _17728_ (.A(_09192_),
    .Y(_09193_));
 sky130_fd_sc_hd__and4b_1 _17729_ (.A_N(_09191_),
    .B(_09192_),
    .C(net312),
    .D(net100),
    .X(_09194_));
 sky130_fd_sc_hd__o2bb2a_1 _17730_ (.A1_N(net312),
    .A2_N(net100),
    .B1(_09191_),
    .B2(_09193_),
    .X(_09195_));
 sky130_fd_sc_hd__or2_1 _17731_ (.A(_09194_),
    .B(_09195_),
    .X(_09196_));
 sky130_fd_sc_hd__or2_2 _17732_ (.A(_09074_),
    .B(_09077_),
    .X(_09197_));
 sky130_fd_sc_hd__nand2b_1 _17733_ (.A_N(_09196_),
    .B(_09197_),
    .Y(_09198_));
 sky130_fd_sc_hd__xor2_2 _17734_ (.A(_09196_),
    .B(_09197_),
    .X(_09199_));
 sky130_fd_sc_hd__or2_1 _17735_ (.A(_09190_),
    .B(_09199_),
    .X(_09200_));
 sky130_fd_sc_hd__xor2_2 _17736_ (.A(_09190_),
    .B(_09199_),
    .X(_09201_));
 sky130_fd_sc_hd__or2_1 _17737_ (.A(_09085_),
    .B(_09087_),
    .X(_09202_));
 sky130_fd_sc_hd__a32o_1 _17738_ (.A1(net287),
    .A2(net129),
    .A3(_09104_),
    .B1(_09103_),
    .B2(net138),
    .X(_09203_));
 sky130_fd_sc_hd__nand4_2 _17739_ (.A(net287),
    .B(net292),
    .C(net122),
    .D(net117),
    .Y(_09204_));
 sky130_fd_sc_hd__a22o_1 _17740_ (.A1(net287),
    .A2(net122),
    .B1(net117),
    .B2(net292),
    .X(_09205_));
 sky130_fd_sc_hd__nand4_2 _17741_ (.A(\mul1.a[6] ),
    .B(net114),
    .C(_09204_),
    .D(_09205_),
    .Y(_09206_));
 sky130_fd_sc_hd__a22o_1 _17742_ (.A1(\mul1.a[6] ),
    .A2(net114),
    .B1(_09204_),
    .B2(_09205_),
    .X(_09207_));
 sky130_fd_sc_hd__and3_1 _17743_ (.A(_09203_),
    .B(_09206_),
    .C(_09207_),
    .X(_09208_));
 sky130_fd_sc_hd__a21o_1 _17744_ (.A1(_09206_),
    .A2(_09207_),
    .B1(_09203_),
    .X(_09209_));
 sky130_fd_sc_hd__and2b_1 _17745_ (.A_N(_09208_),
    .B(_09209_),
    .X(_09210_));
 sky130_fd_sc_hd__xnor2_1 _17746_ (.A(_09202_),
    .B(_09210_),
    .Y(_09211_));
 sky130_fd_sc_hd__a21oi_1 _17747_ (.A1(_09089_),
    .A2(_09092_),
    .B1(_09211_),
    .Y(_09212_));
 sky130_fd_sc_hd__a21o_1 _17748_ (.A1(_09089_),
    .A2(_09092_),
    .B1(_09211_),
    .X(_09213_));
 sky130_fd_sc_hd__nand3_1 _17749_ (.A(_09089_),
    .B(_09092_),
    .C(_09211_),
    .Y(_09214_));
 sky130_fd_sc_hd__and3_2 _17750_ (.A(_09201_),
    .B(_09213_),
    .C(_09214_),
    .X(_09215_));
 sky130_fd_sc_hd__a21oi_2 _17751_ (.A1(_09213_),
    .A2(_09214_),
    .B1(_09201_),
    .Y(_09216_));
 sky130_fd_sc_hd__a211o_2 _17752_ (.A1(_09117_),
    .A2(_09120_),
    .B1(_09215_),
    .C1(_09216_),
    .X(_09217_));
 sky130_fd_sc_hd__o211ai_4 _17753_ (.A1(_09215_),
    .A2(_09216_),
    .B1(_09117_),
    .C1(_09120_),
    .Y(_09218_));
 sky130_fd_sc_hd__o211ai_4 _17754_ (.A1(_09094_),
    .A2(_09096_),
    .B1(_09217_),
    .C1(_09218_),
    .Y(_09219_));
 sky130_fd_sc_hd__a211o_1 _17755_ (.A1(_09217_),
    .A2(_09218_),
    .B1(_09094_),
    .C1(_09096_),
    .X(_09220_));
 sky130_fd_sc_hd__a21o_1 _17756_ (.A1(_09122_),
    .A2(_09128_),
    .B1(_09127_),
    .X(_09221_));
 sky130_fd_sc_hd__nand2_1 _17757_ (.A(net282),
    .B(net129),
    .Y(_09222_));
 sky130_fd_sc_hd__and3_1 _17758_ (.A(net271),
    .B(net277),
    .C(net133),
    .X(_09223_));
 sky130_fd_sc_hd__a22o_1 _17759_ (.A1(net271),
    .A2(net138),
    .B1(net133),
    .B2(net277),
    .X(_09224_));
 sky130_fd_sc_hd__a21bo_1 _17760_ (.A1(net138),
    .A2(_09223_),
    .B1_N(_09224_),
    .X(_09225_));
 sky130_fd_sc_hd__xor2_1 _17761_ (.A(_09222_),
    .B(_09225_),
    .X(_09226_));
 sky130_fd_sc_hd__and2_1 _17762_ (.A(net267),
    .B(net144),
    .X(_09227_));
 sky130_fd_sc_hd__nand4_2 _17763_ (.A(net256),
    .B(net262),
    .C(net152),
    .D(net147),
    .Y(_09228_));
 sky130_fd_sc_hd__a22o_1 _17764_ (.A1(net256),
    .A2(net152),
    .B1(net147),
    .B2(net262),
    .X(_09229_));
 sky130_fd_sc_hd__nand3_1 _17765_ (.A(_09227_),
    .B(_09228_),
    .C(_09229_),
    .Y(_09230_));
 sky130_fd_sc_hd__a21o_1 _17766_ (.A1(_09228_),
    .A2(_09229_),
    .B1(_09227_),
    .X(_09231_));
 sky130_fd_sc_hd__a32o_1 _17767_ (.A1(net271),
    .A2(net144),
    .A3(_09109_),
    .B1(_09108_),
    .B2(net152),
    .X(_09232_));
 sky130_fd_sc_hd__nand3_1 _17768_ (.A(_09230_),
    .B(_09231_),
    .C(_09232_),
    .Y(_09233_));
 sky130_fd_sc_hd__a21o_1 _17769_ (.A1(_09230_),
    .A2(_09231_),
    .B1(_09232_),
    .X(_09234_));
 sky130_fd_sc_hd__nand3_2 _17770_ (.A(_09226_),
    .B(_09233_),
    .C(_09234_),
    .Y(_09235_));
 sky130_fd_sc_hd__a21o_1 _17771_ (.A1(_09233_),
    .A2(_09234_),
    .B1(_09226_),
    .X(_09236_));
 sky130_fd_sc_hd__nand3_4 _17772_ (.A(_09221_),
    .B(_09235_),
    .C(_09236_),
    .Y(_09237_));
 sky130_fd_sc_hd__a21o_1 _17773_ (.A1(_09235_),
    .A2(_09236_),
    .B1(_09221_),
    .X(_09238_));
 sky130_fd_sc_hd__o211ai_4 _17774_ (.A1(_09113_),
    .A2(_09115_),
    .B1(_09237_),
    .C1(_09238_),
    .Y(_09239_));
 sky130_fd_sc_hd__a211o_1 _17775_ (.A1(_09237_),
    .A2(_09238_),
    .B1(_09113_),
    .C1(_09115_),
    .X(_09240_));
 sky130_fd_sc_hd__nand2_1 _17776_ (.A(_09239_),
    .B(_09240_),
    .Y(_09241_));
 sky130_fd_sc_hd__nand2_1 _17777_ (.A(_09123_),
    .B(_09125_),
    .Y(_09242_));
 sky130_fd_sc_hd__nand4_2 _17778_ (.A(net247),
    .B(net629),
    .C(net169),
    .D(net162),
    .Y(_09243_));
 sky130_fd_sc_hd__a22o_1 _17779_ (.A1(net247),
    .A2(net169),
    .B1(net162),
    .B2(net630),
    .X(_09244_));
 sky130_fd_sc_hd__nand4_2 _17780_ (.A(net251),
    .B(net157),
    .C(_09243_),
    .D(_09244_),
    .Y(_09245_));
 sky130_fd_sc_hd__a22o_1 _17781_ (.A1(net251),
    .A2(net157),
    .B1(_09243_),
    .B2(_09244_),
    .X(_09246_));
 sky130_fd_sc_hd__o211a_1 _17782_ (.A1(_09132_),
    .A2(_09133_),
    .B1(_09245_),
    .C1(_09246_),
    .X(_09247_));
 sky130_fd_sc_hd__a211o_1 _17783_ (.A1(_09245_),
    .A2(_09246_),
    .B1(_09132_),
    .C1(_09133_),
    .X(_09248_));
 sky130_fd_sc_hd__nand2b_1 _17784_ (.A_N(_09247_),
    .B(_09248_),
    .Y(_09249_));
 sky130_fd_sc_hd__xnor2_2 _17785_ (.A(_09242_),
    .B(_09249_),
    .Y(_09250_));
 sky130_fd_sc_hd__nand2_1 _17786_ (.A(net173),
    .B(net240),
    .Y(_09251_));
 sky130_fd_sc_hd__a22o_1 _17787_ (.A1(net179),
    .A2(net235),
    .B1(net232),
    .B2(net184),
    .X(_09252_));
 sky130_fd_sc_hd__and3_1 _17788_ (.A(net184),
    .B(net179),
    .C(net235),
    .X(_09253_));
 sky130_fd_sc_hd__a21bo_1 _17789_ (.A1(net232),
    .A2(_09253_),
    .B1_N(_09252_),
    .X(_09254_));
 sky130_fd_sc_hd__xor2_2 _17790_ (.A(_09251_),
    .B(_09254_),
    .X(_09255_));
 sky130_fd_sc_hd__and2_1 _17791_ (.A(\mul1.b[2] ),
    .B(net227),
    .X(_09256_));
 sky130_fd_sc_hd__nand4_1 _17792_ (.A(net623),
    .B(net190),
    .C(net221),
    .D(net218),
    .Y(_09257_));
 sky130_fd_sc_hd__a22o_1 _17793_ (.A1(net190),
    .A2(net221),
    .B1(net215),
    .B2(net623),
    .X(_09258_));
 sky130_fd_sc_hd__nand3_1 _17794_ (.A(_09256_),
    .B(_09257_),
    .C(_09258_),
    .Y(_09259_));
 sky130_fd_sc_hd__a21o_1 _17795_ (.A1(_09257_),
    .A2(_09258_),
    .B1(_09256_),
    .X(_09260_));
 sky130_fd_sc_hd__a21bo_1 _17796_ (.A1(_09136_),
    .A2(_09138_),
    .B1_N(_09137_),
    .X(_09261_));
 sky130_fd_sc_hd__nand3_1 _17797_ (.A(_09259_),
    .B(_09260_),
    .C(_09261_),
    .Y(_09262_));
 sky130_fd_sc_hd__a21o_1 _17798_ (.A1(_09259_),
    .A2(_09260_),
    .B1(_09261_),
    .X(_09263_));
 sky130_fd_sc_hd__nand3_2 _17799_ (.A(_09255_),
    .B(_09262_),
    .C(_09263_),
    .Y(_09264_));
 sky130_fd_sc_hd__a21o_1 _17800_ (.A1(_09262_),
    .A2(_09263_),
    .B1(_09255_),
    .X(_09265_));
 sky130_fd_sc_hd__a21bo_1 _17801_ (.A1(_09135_),
    .A2(_09143_),
    .B1_N(_09142_),
    .X(_09266_));
 sky130_fd_sc_hd__nand3_4 _17802_ (.A(_09264_),
    .B(_09265_),
    .C(_09266_),
    .Y(_09267_));
 sky130_fd_sc_hd__a21o_1 _17803_ (.A1(_09264_),
    .A2(_09265_),
    .B1(_09266_),
    .X(_09268_));
 sky130_fd_sc_hd__and3_1 _17804_ (.A(_09250_),
    .B(_09267_),
    .C(_09268_),
    .X(_09269_));
 sky130_fd_sc_hd__nand3_2 _17805_ (.A(_09250_),
    .B(_09267_),
    .C(_09268_),
    .Y(_09270_));
 sky130_fd_sc_hd__a21oi_2 _17806_ (.A1(_09267_),
    .A2(_09268_),
    .B1(_09250_),
    .Y(_09271_));
 sky130_fd_sc_hd__a211oi_4 _17807_ (.A1(_09147_),
    .A2(_09150_),
    .B1(_09269_),
    .C1(_09271_),
    .Y(_09272_));
 sky130_fd_sc_hd__o211a_1 _17808_ (.A1(_09269_),
    .A2(_09271_),
    .B1(_09147_),
    .C1(_09150_),
    .X(_09273_));
 sky130_fd_sc_hd__nor3_1 _17809_ (.A(_09241_),
    .B(_09272_),
    .C(_09273_),
    .Y(_09274_));
 sky130_fd_sc_hd__or3_2 _17810_ (.A(_09241_),
    .B(_09272_),
    .C(_09273_),
    .X(_09275_));
 sky130_fd_sc_hd__o21ai_2 _17811_ (.A1(_09272_),
    .A2(_09273_),
    .B1(_09241_),
    .Y(_09276_));
 sky130_fd_sc_hd__o211a_1 _17812_ (.A1(_09152_),
    .A2(_09154_),
    .B1(_09275_),
    .C1(_09276_),
    .X(_09277_));
 sky130_fd_sc_hd__o211ai_2 _17813_ (.A1(_09152_),
    .A2(_09154_),
    .B1(_09275_),
    .C1(_09276_),
    .Y(_09278_));
 sky130_fd_sc_hd__a211o_1 _17814_ (.A1(_09275_),
    .A2(_09276_),
    .B1(_09152_),
    .C1(_09154_),
    .X(_09279_));
 sky130_fd_sc_hd__and4_2 _17815_ (.A(_09219_),
    .B(_09220_),
    .C(_09278_),
    .D(_09279_),
    .X(_09280_));
 sky130_fd_sc_hd__a22oi_2 _17816_ (.A1(_09219_),
    .A2(_09220_),
    .B1(_09278_),
    .B2(_09279_),
    .Y(_09281_));
 sky130_fd_sc_hd__a211o_2 _17817_ (.A1(_09157_),
    .A2(_09160_),
    .B1(_09280_),
    .C1(_09281_),
    .X(_09282_));
 sky130_fd_sc_hd__o211ai_2 _17818_ (.A1(_09280_),
    .A2(_09281_),
    .B1(_09157_),
    .C1(_09160_),
    .Y(_09283_));
 sky130_fd_sc_hd__nand3_2 _17819_ (.A(_09184_),
    .B(_09282_),
    .C(_09283_),
    .Y(_09284_));
 sky130_fd_sc_hd__a21o_1 _17820_ (.A1(_09282_),
    .A2(_09283_),
    .B1(_09184_),
    .X(_09285_));
 sky130_fd_sc_hd__nand2_1 _17821_ (.A(_09284_),
    .B(_09285_),
    .Y(_09286_));
 sky130_fd_sc_hd__o21ba_1 _17822_ (.A1(_09069_),
    .A2(_09163_),
    .B1_N(_09162_),
    .X(_09287_));
 sky130_fd_sc_hd__or2_1 _17823_ (.A(_09286_),
    .B(_09287_),
    .X(_09288_));
 sky130_fd_sc_hd__xor2_1 _17824_ (.A(_09286_),
    .B(_09287_),
    .X(_09289_));
 sky130_fd_sc_hd__xnor2_1 _17825_ (.A(_09067_),
    .B(_09289_),
    .Y(_09290_));
 sky130_fd_sc_hd__o21a_1 _17826_ (.A1(_08955_),
    .A2(_09169_),
    .B1(_09168_),
    .X(_09291_));
 sky130_fd_sc_hd__nor2_2 _17827_ (.A(_09290_),
    .B(_09291_),
    .Y(_09292_));
 sky130_fd_sc_hd__xnor2_1 _17828_ (.A(_09290_),
    .B(_09291_),
    .Y(_09293_));
 sky130_fd_sc_hd__o21ai_1 _17829_ (.A1(_09055_),
    .A2(_09170_),
    .B1(_09293_),
    .Y(_09294_));
 sky130_fd_sc_hd__or3_1 _17830_ (.A(_09055_),
    .B(_09170_),
    .C(_09293_),
    .X(_09295_));
 sky130_fd_sc_hd__nand2_2 _17831_ (.A(_09294_),
    .B(_09295_),
    .Y(_09296_));
 sky130_fd_sc_hd__xnor2_4 _17832_ (.A(_09178_),
    .B(_09296_),
    .Y(_09297_));
 sky130_fd_sc_hd__nor2_1 _17833_ (.A(_03049_),
    .B(_09297_),
    .Y(_09298_));
 sky130_fd_sc_hd__nor2_1 _17834_ (.A(net44),
    .B(_04449_),
    .Y(_09299_));
 sky130_fd_sc_hd__a21o_1 _17835_ (.A1(net742),
    .A2(net7),
    .B1(_03056_),
    .X(_09300_));
 sky130_fd_sc_hd__o32a_1 _17836_ (.A1(_09298_),
    .A2(_09299_),
    .A3(_09300_),
    .B1(net2),
    .B2(net726),
    .X(_00305_));
 sky130_fd_sc_hd__or2_2 _17837_ (.A(_09173_),
    .B(_09293_),
    .X(_09301_));
 sky130_fd_sc_hd__a211o_1 _17838_ (.A1(_09055_),
    .A2(_09293_),
    .B1(_09171_),
    .C1(_09170_),
    .X(_09302_));
 sky130_fd_sc_hd__o211a_1 _17839_ (.A1(_09174_),
    .A2(_09301_),
    .B1(_09302_),
    .C1(_09295_),
    .X(_09303_));
 sky130_fd_sc_hd__o31a_2 _17840_ (.A1(_08950_),
    .A2(_09059_),
    .A3(_09301_),
    .B1(_09303_),
    .X(_09304_));
 sky130_fd_sc_hd__o31ai_4 _17841_ (.A1(_08950_),
    .A2(_09059_),
    .A3(_09301_),
    .B1(_09303_),
    .Y(_09305_));
 sky130_fd_sc_hd__a21bo_2 _17842_ (.A1(_09067_),
    .A2(_09289_),
    .B1_N(_09288_),
    .X(_09306_));
 sky130_fd_sc_hd__o211a_1 _17843_ (.A1(_09185_),
    .A2(_09188_),
    .B1(net324),
    .C1(net82),
    .X(_09307_));
 sky130_fd_sc_hd__a211oi_1 _17844_ (.A1(net324),
    .A2(net82),
    .B1(_09185_),
    .C1(_09188_),
    .Y(_09308_));
 sky130_fd_sc_hd__or2_1 _17845_ (.A(_09307_),
    .B(_09308_),
    .X(_09309_));
 sky130_fd_sc_hd__a21oi_1 _17846_ (.A1(_09198_),
    .A2(_09200_),
    .B1(_09309_),
    .Y(_09310_));
 sky130_fd_sc_hd__and3_1 _17847_ (.A(_09198_),
    .B(_09200_),
    .C(_09309_),
    .X(_09311_));
 sky130_fd_sc_hd__nor2_1 _17848_ (.A(_09310_),
    .B(_09311_),
    .Y(_09312_));
 sky130_fd_sc_hd__nand2_1 _17849_ (.A(_09179_),
    .B(_09312_),
    .Y(_09313_));
 sky130_fd_sc_hd__xnor2_1 _17850_ (.A(_09179_),
    .B(_09312_),
    .Y(_09314_));
 sky130_fd_sc_hd__a21oi_2 _17851_ (.A1(_09217_),
    .A2(_09219_),
    .B1(_09314_),
    .Y(_09315_));
 sky130_fd_sc_hd__and3_1 _17852_ (.A(_09217_),
    .B(_09219_),
    .C(_09314_),
    .X(_09316_));
 sky130_fd_sc_hd__nor2_1 _17853_ (.A(_09315_),
    .B(_09316_),
    .Y(_09317_));
 sky130_fd_sc_hd__and4_1 _17854_ (.A(net312),
    .B(net317),
    .C(net94),
    .D(net89),
    .X(_09318_));
 sky130_fd_sc_hd__inv_2 _17855_ (.A(_09318_),
    .Y(_09319_));
 sky130_fd_sc_hd__a22o_1 _17856_ (.A1(net312),
    .A2(net94),
    .B1(net89),
    .B2(net317),
    .X(_09320_));
 sky130_fd_sc_hd__and4_1 _17857_ (.A(net321),
    .B(net85),
    .C(_09319_),
    .D(_09320_),
    .X(_09321_));
 sky130_fd_sc_hd__a22oi_1 _17858_ (.A1(net321),
    .A2(net85),
    .B1(_09319_),
    .B2(_09320_),
    .Y(_09322_));
 sky130_fd_sc_hd__or2_1 _17859_ (.A(_09321_),
    .B(_09322_),
    .X(_09323_));
 sky130_fd_sc_hd__nand2_1 _17860_ (.A(net307),
    .B(net100),
    .Y(_09324_));
 sky130_fd_sc_hd__and4_1 _17861_ (.A(net296),
    .B(net301),
    .C(net108),
    .D(net103),
    .X(_09325_));
 sky130_fd_sc_hd__a22o_1 _17862_ (.A1(net296),
    .A2(net108),
    .B1(net103),
    .B2(net301),
    .X(_09326_));
 sky130_fd_sc_hd__and2b_1 _17863_ (.A_N(_09325_),
    .B(_09326_),
    .X(_09327_));
 sky130_fd_sc_hd__xnor2_2 _17864_ (.A(_09324_),
    .B(_09327_),
    .Y(_09328_));
 sky130_fd_sc_hd__nor2_1 _17865_ (.A(_09191_),
    .B(_09194_),
    .Y(_09329_));
 sky130_fd_sc_hd__nand2b_1 _17866_ (.A_N(_09329_),
    .B(_09328_),
    .Y(_09330_));
 sky130_fd_sc_hd__xnor2_2 _17867_ (.A(_09328_),
    .B(_09329_),
    .Y(_09331_));
 sky130_fd_sc_hd__nand2b_1 _17868_ (.A_N(_09323_),
    .B(_09331_),
    .Y(_09332_));
 sky130_fd_sc_hd__xnor2_2 _17869_ (.A(_09323_),
    .B(_09331_),
    .Y(_09333_));
 sky130_fd_sc_hd__nand2_1 _17870_ (.A(_09204_),
    .B(_09206_),
    .Y(_09334_));
 sky130_fd_sc_hd__a32o_1 _17871_ (.A1(net282),
    .A2(net129),
    .A3(_09224_),
    .B1(_09223_),
    .B2(net138),
    .X(_09335_));
 sky130_fd_sc_hd__nand4_2 _17872_ (.A(net282),
    .B(net287),
    .C(net125),
    .D(net120),
    .Y(_09336_));
 sky130_fd_sc_hd__a22o_1 _17873_ (.A1(net282),
    .A2(net125),
    .B1(net120),
    .B2(net287),
    .X(_09337_));
 sky130_fd_sc_hd__nand4_2 _17874_ (.A(net292),
    .B(net116),
    .C(_09336_),
    .D(_09337_),
    .Y(_09338_));
 sky130_fd_sc_hd__a22o_1 _17875_ (.A1(net292),
    .A2(net114),
    .B1(_09336_),
    .B2(_09337_),
    .X(_09339_));
 sky130_fd_sc_hd__nand3_1 _17876_ (.A(_09335_),
    .B(_09338_),
    .C(_09339_),
    .Y(_09340_));
 sky130_fd_sc_hd__a21o_1 _17877_ (.A1(_09338_),
    .A2(_09339_),
    .B1(_09335_),
    .X(_09341_));
 sky130_fd_sc_hd__nand3_1 _17878_ (.A(_09334_),
    .B(_09340_),
    .C(_09341_),
    .Y(_09342_));
 sky130_fd_sc_hd__a21o_1 _17879_ (.A1(_09340_),
    .A2(_09341_),
    .B1(_09334_),
    .X(_09343_));
 sky130_fd_sc_hd__a21o_1 _17880_ (.A1(_09202_),
    .A2(_09209_),
    .B1(_09208_),
    .X(_09344_));
 sky130_fd_sc_hd__nand3_2 _17881_ (.A(_09342_),
    .B(_09343_),
    .C(_09344_),
    .Y(_09345_));
 sky130_fd_sc_hd__a21o_1 _17882_ (.A1(_09342_),
    .A2(_09343_),
    .B1(_09344_),
    .X(_09346_));
 sky130_fd_sc_hd__and3_1 _17883_ (.A(_09333_),
    .B(_09345_),
    .C(_09346_),
    .X(_09347_));
 sky130_fd_sc_hd__inv_2 _17884_ (.A(_09347_),
    .Y(_09348_));
 sky130_fd_sc_hd__a21oi_1 _17885_ (.A1(_09345_),
    .A2(_09346_),
    .B1(_09333_),
    .Y(_09349_));
 sky130_fd_sc_hd__a211o_1 _17886_ (.A1(_09237_),
    .A2(_09239_),
    .B1(_09347_),
    .C1(_09349_),
    .X(_09350_));
 sky130_fd_sc_hd__o211ai_2 _17887_ (.A1(_09347_),
    .A2(_09349_),
    .B1(_09237_),
    .C1(_09239_),
    .Y(_09351_));
 sky130_fd_sc_hd__o211ai_1 _17888_ (.A1(_09212_),
    .A2(_09215_),
    .B1(_09350_),
    .C1(_09351_),
    .Y(_09352_));
 sky130_fd_sc_hd__a211o_1 _17889_ (.A1(_09350_),
    .A2(_09351_),
    .B1(_09212_),
    .C1(_09215_),
    .X(_09353_));
 sky130_fd_sc_hd__nand2_1 _17890_ (.A(_09352_),
    .B(_09353_),
    .Y(_09354_));
 sky130_fd_sc_hd__nand2_1 _17891_ (.A(_09233_),
    .B(_09235_),
    .Y(_09355_));
 sky130_fd_sc_hd__a21o_1 _17892_ (.A1(_09242_),
    .A2(_09248_),
    .B1(_09247_),
    .X(_09356_));
 sky130_fd_sc_hd__nand2_1 _17893_ (.A(net277),
    .B(net129),
    .Y(_09357_));
 sky130_fd_sc_hd__and3_1 _17894_ (.A(net267),
    .B(net271),
    .C(net133),
    .X(_09358_));
 sky130_fd_sc_hd__a22o_1 _17895_ (.A1(net267),
    .A2(net138),
    .B1(net133),
    .B2(net271),
    .X(_09359_));
 sky130_fd_sc_hd__a21bo_1 _17896_ (.A1(net138),
    .A2(_09358_),
    .B1_N(_09359_),
    .X(_09360_));
 sky130_fd_sc_hd__xor2_1 _17897_ (.A(_09357_),
    .B(_09360_),
    .X(_09361_));
 sky130_fd_sc_hd__and2_1 _17898_ (.A(net262),
    .B(net144),
    .X(_09362_));
 sky130_fd_sc_hd__nand4_1 _17899_ (.A(net251),
    .B(net256),
    .C(net152),
    .D(net147),
    .Y(_09363_));
 sky130_fd_sc_hd__a22o_1 _17900_ (.A1(net251),
    .A2(net152),
    .B1(net147),
    .B2(net256),
    .X(_09364_));
 sky130_fd_sc_hd__nand3_1 _17901_ (.A(_09362_),
    .B(_09363_),
    .C(_09364_),
    .Y(_09365_));
 sky130_fd_sc_hd__a21o_1 _17902_ (.A1(_09363_),
    .A2(_09364_),
    .B1(_09362_),
    .X(_09366_));
 sky130_fd_sc_hd__a21bo_1 _17903_ (.A1(_09227_),
    .A2(_09229_),
    .B1_N(_09228_),
    .X(_09367_));
 sky130_fd_sc_hd__nand3_1 _17904_ (.A(_09365_),
    .B(_09366_),
    .C(_09367_),
    .Y(_09368_));
 sky130_fd_sc_hd__a21o_1 _17905_ (.A1(_09365_),
    .A2(_09366_),
    .B1(_09367_),
    .X(_09369_));
 sky130_fd_sc_hd__nand3_2 _17906_ (.A(_09361_),
    .B(_09368_),
    .C(_09369_),
    .Y(_09370_));
 sky130_fd_sc_hd__a21o_1 _17907_ (.A1(_09368_),
    .A2(_09369_),
    .B1(_09361_),
    .X(_09371_));
 sky130_fd_sc_hd__nand3_2 _17908_ (.A(_09356_),
    .B(_09370_),
    .C(_09371_),
    .Y(_09372_));
 sky130_fd_sc_hd__a21o_1 _17909_ (.A1(_09370_),
    .A2(_09371_),
    .B1(_09356_),
    .X(_09373_));
 sky130_fd_sc_hd__nand3_2 _17910_ (.A(_09355_),
    .B(_09372_),
    .C(_09373_),
    .Y(_09374_));
 sky130_fd_sc_hd__a21o_1 _17911_ (.A1(_09372_),
    .A2(_09373_),
    .B1(_09355_),
    .X(_09375_));
 sky130_fd_sc_hd__nand2_1 _17912_ (.A(_09374_),
    .B(_09375_),
    .Y(_09376_));
 sky130_fd_sc_hd__nand2_1 _17913_ (.A(_09243_),
    .B(_09245_),
    .Y(_09377_));
 sky130_fd_sc_hd__a32o_1 _17914_ (.A1(net173),
    .A2(net240),
    .A3(_09252_),
    .B1(_09253_),
    .B2(net232),
    .X(_09378_));
 sky130_fd_sc_hd__nand4_2 _17915_ (.A(net247),
    .B(net169),
    .C(net162),
    .D(net240),
    .Y(_09379_));
 sky130_fd_sc_hd__a22o_1 _17916_ (.A1(net247),
    .A2(net162),
    .B1(net240),
    .B2(net169),
    .X(_09380_));
 sky130_fd_sc_hd__nand4_2 _17917_ (.A(net629),
    .B(net157),
    .C(_09379_),
    .D(_09380_),
    .Y(_09381_));
 sky130_fd_sc_hd__a22o_1 _17918_ (.A1(net629),
    .A2(net157),
    .B1(_09379_),
    .B2(_09380_),
    .X(_09382_));
 sky130_fd_sc_hd__nand3_1 _17919_ (.A(_09378_),
    .B(_09381_),
    .C(_09382_),
    .Y(_09383_));
 sky130_fd_sc_hd__a21o_1 _17920_ (.A1(_09381_),
    .A2(_09382_),
    .B1(_09378_),
    .X(_09384_));
 sky130_fd_sc_hd__and3_1 _17921_ (.A(_09377_),
    .B(_09383_),
    .C(_09384_),
    .X(_09385_));
 sky130_fd_sc_hd__a21oi_1 _17922_ (.A1(_09383_),
    .A2(_09384_),
    .B1(_09377_),
    .Y(_09386_));
 sky130_fd_sc_hd__nor2_1 _17923_ (.A(_09385_),
    .B(_09386_),
    .Y(_09387_));
 sky130_fd_sc_hd__nand2_1 _17924_ (.A(net175),
    .B(net235),
    .Y(_09388_));
 sky130_fd_sc_hd__and4_1 _17925_ (.A(net184),
    .B(net179),
    .C(net229),
    .D(net225),
    .X(_09389_));
 sky130_fd_sc_hd__a22oi_2 _17926_ (.A1(net179),
    .A2(net229),
    .B1(net225),
    .B2(net184),
    .Y(_09390_));
 sky130_fd_sc_hd__nor2_1 _17927_ (.A(_09389_),
    .B(_09390_),
    .Y(_09391_));
 sky130_fd_sc_hd__xnor2_2 _17928_ (.A(_09388_),
    .B(_09391_),
    .Y(_09392_));
 sky130_fd_sc_hd__and2_1 _17929_ (.A(\mul1.b[2] ),
    .B(net219),
    .X(_09393_));
 sky130_fd_sc_hd__nand4_2 _17930_ (.A(net623),
    .B(net190),
    .C(net215),
    .D(net211),
    .Y(_09394_));
 sky130_fd_sc_hd__a22o_1 _17931_ (.A1(net190),
    .A2(net215),
    .B1(net211),
    .B2(net623),
    .X(_09395_));
 sky130_fd_sc_hd__nand3_1 _17932_ (.A(_09393_),
    .B(_09394_),
    .C(_09395_),
    .Y(_09396_));
 sky130_fd_sc_hd__a21o_1 _17933_ (.A1(_09394_),
    .A2(_09395_),
    .B1(_09393_),
    .X(_09397_));
 sky130_fd_sc_hd__a21bo_1 _17934_ (.A1(_09256_),
    .A2(_09258_),
    .B1_N(_09257_),
    .X(_09398_));
 sky130_fd_sc_hd__nand3_2 _17935_ (.A(_09396_),
    .B(_09397_),
    .C(_09398_),
    .Y(_09399_));
 sky130_fd_sc_hd__a21o_1 _17936_ (.A1(_09396_),
    .A2(_09397_),
    .B1(_09398_),
    .X(_09400_));
 sky130_fd_sc_hd__nand3_2 _17937_ (.A(_09392_),
    .B(_09399_),
    .C(_09400_),
    .Y(_09401_));
 sky130_fd_sc_hd__a21o_1 _17938_ (.A1(_09399_),
    .A2(_09400_),
    .B1(_09392_),
    .X(_09402_));
 sky130_fd_sc_hd__a21bo_1 _17939_ (.A1(_09255_),
    .A2(_09263_),
    .B1_N(_09262_),
    .X(_09403_));
 sky130_fd_sc_hd__nand3_4 _17940_ (.A(_09401_),
    .B(_09402_),
    .C(_09403_),
    .Y(_09404_));
 sky130_fd_sc_hd__a21o_1 _17941_ (.A1(_09401_),
    .A2(_09402_),
    .B1(_09403_),
    .X(_09405_));
 sky130_fd_sc_hd__and3_1 _17942_ (.A(_09387_),
    .B(_09404_),
    .C(_09405_),
    .X(_09406_));
 sky130_fd_sc_hd__nand3_2 _17943_ (.A(_09387_),
    .B(_09404_),
    .C(_09405_),
    .Y(_09407_));
 sky130_fd_sc_hd__a21oi_2 _17944_ (.A1(_09404_),
    .A2(_09405_),
    .B1(_09387_),
    .Y(_09408_));
 sky130_fd_sc_hd__a211oi_4 _17945_ (.A1(_09267_),
    .A2(_09270_),
    .B1(_09406_),
    .C1(_09408_),
    .Y(_09409_));
 sky130_fd_sc_hd__o211a_1 _17946_ (.A1(_09406_),
    .A2(_09408_),
    .B1(_09267_),
    .C1(_09270_),
    .X(_09410_));
 sky130_fd_sc_hd__nor3_2 _17947_ (.A(_09376_),
    .B(_09409_),
    .C(_09410_),
    .Y(_09411_));
 sky130_fd_sc_hd__or3_1 _17948_ (.A(_09376_),
    .B(_09409_),
    .C(_09410_),
    .X(_09412_));
 sky130_fd_sc_hd__o21ai_1 _17949_ (.A1(_09409_),
    .A2(_09410_),
    .B1(_09376_),
    .Y(_09413_));
 sky130_fd_sc_hd__o211a_2 _17950_ (.A1(_09272_),
    .A2(_09274_),
    .B1(_09412_),
    .C1(_09413_),
    .X(_09414_));
 sky130_fd_sc_hd__a211oi_2 _17951_ (.A1(_09412_),
    .A2(_09413_),
    .B1(_09272_),
    .C1(_09274_),
    .Y(_09415_));
 sky130_fd_sc_hd__nor3_2 _17952_ (.A(_09354_),
    .B(_09414_),
    .C(_09415_),
    .Y(_09416_));
 sky130_fd_sc_hd__or3_2 _17953_ (.A(_09354_),
    .B(_09414_),
    .C(_09415_),
    .X(_09417_));
 sky130_fd_sc_hd__o21ai_2 _17954_ (.A1(_09414_),
    .A2(_09415_),
    .B1(_09354_),
    .Y(_09418_));
 sky130_fd_sc_hd__o211ai_4 _17955_ (.A1(_09277_),
    .A2(_09280_),
    .B1(_09417_),
    .C1(_09418_),
    .Y(_09419_));
 sky130_fd_sc_hd__inv_2 _17956_ (.A(_09419_),
    .Y(_09420_));
 sky130_fd_sc_hd__a211o_1 _17957_ (.A1(_09417_),
    .A2(_09418_),
    .B1(_09277_),
    .C1(_09280_),
    .X(_09421_));
 sky130_fd_sc_hd__and3_2 _17958_ (.A(_09317_),
    .B(_09419_),
    .C(_09421_),
    .X(_09422_));
 sky130_fd_sc_hd__a21oi_2 _17959_ (.A1(_09419_),
    .A2(_09421_),
    .B1(_09317_),
    .Y(_09423_));
 sky130_fd_sc_hd__a211oi_4 _17960_ (.A1(_09282_),
    .A2(_09284_),
    .B1(_09422_),
    .C1(_09423_),
    .Y(_09424_));
 sky130_fd_sc_hd__o211a_1 _17961_ (.A1(_09422_),
    .A2(_09423_),
    .B1(_09282_),
    .C1(_09284_),
    .X(_09425_));
 sky130_fd_sc_hd__nor3_2 _17962_ (.A(_09182_),
    .B(_09424_),
    .C(_09425_),
    .Y(_09426_));
 sky130_fd_sc_hd__o21a_1 _17963_ (.A1(_09424_),
    .A2(_09425_),
    .B1(_09182_),
    .X(_09427_));
 sky130_fd_sc_hd__or2_1 _17964_ (.A(_09426_),
    .B(_09427_),
    .X(_09428_));
 sky130_fd_sc_hd__nand2b_1 _17965_ (.A_N(_09428_),
    .B(_09306_),
    .Y(_09429_));
 sky130_fd_sc_hd__xnor2_2 _17966_ (.A(_09306_),
    .B(_09428_),
    .Y(_09430_));
 sky130_fd_sc_hd__xnor2_1 _17967_ (.A(_09292_),
    .B(_09430_),
    .Y(_09431_));
 sky130_fd_sc_hd__nor2_1 _17968_ (.A(_09304_),
    .B(_09431_),
    .Y(_09432_));
 sky130_fd_sc_hd__nand2_1 _17969_ (.A(_09304_),
    .B(_09431_),
    .Y(_09433_));
 sky130_fd_sc_hd__and2b_2 _17970_ (.A_N(_09432_),
    .B(_09433_),
    .X(_09434_));
 sky130_fd_sc_hd__nor2_1 _17971_ (.A(net43),
    .B(_04588_),
    .Y(_09435_));
 sky130_fd_sc_hd__a221o_1 _17972_ (.A1(\temp[7] ),
    .A2(net8),
    .B1(_09434_),
    .B2(net10),
    .C1(_09435_),
    .X(_09436_));
 sky130_fd_sc_hd__mux2_1 _17973_ (.A0(net750),
    .A1(_09436_),
    .S(net2),
    .X(_00306_));
 sky130_fd_sc_hd__a21oi_2 _17974_ (.A1(_09292_),
    .A2(_09430_),
    .B1(_09432_),
    .Y(_09437_));
 sky130_fd_sc_hd__and2_1 _17975_ (.A(_09350_),
    .B(_09352_),
    .X(_09438_));
 sky130_fd_sc_hd__a22oi_1 _17976_ (.A1(net321),
    .A2(net82),
    .B1(\mul1.b[25] ),
    .B2(net324),
    .Y(_09439_));
 sky130_fd_sc_hd__and4_1 _17977_ (.A(\mul1.a[1] ),
    .B(net324),
    .C(net82),
    .D(net78),
    .X(_09440_));
 sky130_fd_sc_hd__nor2_1 _17978_ (.A(_09439_),
    .B(_09440_),
    .Y(_09441_));
 sky130_fd_sc_hd__o21ai_2 _17979_ (.A1(_09318_),
    .A2(_09321_),
    .B1(_09441_),
    .Y(_09442_));
 sky130_fd_sc_hd__or3_1 _17980_ (.A(_09318_),
    .B(_09321_),
    .C(_09441_),
    .X(_09443_));
 sky130_fd_sc_hd__nand2_1 _17981_ (.A(_09442_),
    .B(_09443_),
    .Y(_09444_));
 sky130_fd_sc_hd__nand3_2 _17982_ (.A(_09330_),
    .B(_09332_),
    .C(_09444_),
    .Y(_09445_));
 sky130_fd_sc_hd__inv_2 _17983_ (.A(_09445_),
    .Y(_09446_));
 sky130_fd_sc_hd__a21oi_1 _17984_ (.A1(_09330_),
    .A2(_09332_),
    .B1(_09444_),
    .Y(_09447_));
 sky130_fd_sc_hd__or2_1 _17985_ (.A(_09446_),
    .B(_09447_),
    .X(_09448_));
 sky130_fd_sc_hd__nor2_1 _17986_ (.A(_09307_),
    .B(_09310_),
    .Y(_09449_));
 sky130_fd_sc_hd__xnor2_2 _17987_ (.A(_09448_),
    .B(_09449_),
    .Y(_09450_));
 sky130_fd_sc_hd__nor2_1 _17988_ (.A(_09438_),
    .B(_09450_),
    .Y(_09451_));
 sky130_fd_sc_hd__xor2_2 _17989_ (.A(_09438_),
    .B(_09450_),
    .X(_09452_));
 sky130_fd_sc_hd__xnor2_2 _17990_ (.A(_09313_),
    .B(_09452_),
    .Y(_09453_));
 sky130_fd_sc_hd__and4_1 _17991_ (.A(net306),
    .B(net311),
    .C(net93),
    .D(net89),
    .X(_09454_));
 sky130_fd_sc_hd__a22o_1 _17992_ (.A1(net306),
    .A2(net93),
    .B1(net89),
    .B2(net311),
    .X(_09455_));
 sky130_fd_sc_hd__nand2b_1 _17993_ (.A_N(_09454_),
    .B(_09455_),
    .Y(_09456_));
 sky130_fd_sc_hd__nand2_1 _17994_ (.A(net316),
    .B(net85),
    .Y(_09457_));
 sky130_fd_sc_hd__xnor2_2 _17995_ (.A(_09456_),
    .B(_09457_),
    .Y(_09458_));
 sky130_fd_sc_hd__and2_1 _17996_ (.A(net301),
    .B(net99),
    .X(_09459_));
 sky130_fd_sc_hd__nand4_2 _17997_ (.A(net290),
    .B(net296),
    .C(net108),
    .D(net103),
    .Y(_09460_));
 sky130_fd_sc_hd__a22o_1 _17998_ (.A1(net290),
    .A2(net108),
    .B1(net103),
    .B2(net296),
    .X(_09461_));
 sky130_fd_sc_hd__nand3_1 _17999_ (.A(_09459_),
    .B(_09460_),
    .C(_09461_),
    .Y(_09462_));
 sky130_fd_sc_hd__a21o_1 _18000_ (.A1(_09460_),
    .A2(_09461_),
    .B1(_09459_),
    .X(_09463_));
 sky130_fd_sc_hd__a31o_1 _18001_ (.A1(net306),
    .A2(net100),
    .A3(_09326_),
    .B1(_09325_),
    .X(_09464_));
 sky130_fd_sc_hd__and3_1 _18002_ (.A(_09462_),
    .B(_09463_),
    .C(_09464_),
    .X(_09465_));
 sky130_fd_sc_hd__a21oi_1 _18003_ (.A1(_09462_),
    .A2(_09463_),
    .B1(_09464_),
    .Y(_09466_));
 sky130_fd_sc_hd__nor2_1 _18004_ (.A(_09465_),
    .B(_09466_),
    .Y(_09467_));
 sky130_fd_sc_hd__xnor2_2 _18005_ (.A(_09458_),
    .B(_09467_),
    .Y(_09468_));
 sky130_fd_sc_hd__nand2_1 _18006_ (.A(_09336_),
    .B(_09338_),
    .Y(_09469_));
 sky130_fd_sc_hd__a32o_1 _18007_ (.A1(net277),
    .A2(net129),
    .A3(_09359_),
    .B1(_09358_),
    .B2(net138),
    .X(_09470_));
 sky130_fd_sc_hd__nand4_2 _18008_ (.A(net277),
    .B(net282),
    .C(net125),
    .D(net120),
    .Y(_09471_));
 sky130_fd_sc_hd__a22o_1 _18009_ (.A1(net277),
    .A2(net125),
    .B1(net120),
    .B2(net282),
    .X(_09472_));
 sky130_fd_sc_hd__nand4_2 _18010_ (.A(net287),
    .B(net116),
    .C(_09471_),
    .D(_09472_),
    .Y(_09473_));
 sky130_fd_sc_hd__a22o_1 _18011_ (.A1(net287),
    .A2(net116),
    .B1(_09471_),
    .B2(_09472_),
    .X(_09474_));
 sky130_fd_sc_hd__nand3_1 _18012_ (.A(_09470_),
    .B(_09473_),
    .C(_09474_),
    .Y(_09475_));
 sky130_fd_sc_hd__a21o_1 _18013_ (.A1(_09473_),
    .A2(_09474_),
    .B1(_09470_),
    .X(_09476_));
 sky130_fd_sc_hd__nand3_1 _18014_ (.A(_09469_),
    .B(_09475_),
    .C(_09476_),
    .Y(_09477_));
 sky130_fd_sc_hd__a21o_1 _18015_ (.A1(_09475_),
    .A2(_09476_),
    .B1(_09469_),
    .X(_09478_));
 sky130_fd_sc_hd__a21bo_1 _18016_ (.A1(_09334_),
    .A2(_09341_),
    .B1_N(_09340_),
    .X(_09479_));
 sky130_fd_sc_hd__and3_1 _18017_ (.A(_09477_),
    .B(_09478_),
    .C(_09479_),
    .X(_09480_));
 sky130_fd_sc_hd__nand3_1 _18018_ (.A(_09477_),
    .B(_09478_),
    .C(_09479_),
    .Y(_09481_));
 sky130_fd_sc_hd__a21o_1 _18019_ (.A1(_09477_),
    .A2(_09478_),
    .B1(_09479_),
    .X(_09482_));
 sky130_fd_sc_hd__and3_1 _18020_ (.A(_09468_),
    .B(_09481_),
    .C(_09482_),
    .X(_09483_));
 sky130_fd_sc_hd__a21oi_1 _18021_ (.A1(_09481_),
    .A2(_09482_),
    .B1(_09468_),
    .Y(_09484_));
 sky130_fd_sc_hd__a211oi_2 _18022_ (.A1(_09372_),
    .A2(_09374_),
    .B1(_09483_),
    .C1(_09484_),
    .Y(_09485_));
 sky130_fd_sc_hd__o211a_1 _18023_ (.A1(_09483_),
    .A2(_09484_),
    .B1(_09372_),
    .C1(_09374_),
    .X(_09486_));
 sky130_fd_sc_hd__a211oi_4 _18024_ (.A1(_09345_),
    .A2(_09348_),
    .B1(_09485_),
    .C1(_09486_),
    .Y(_09487_));
 sky130_fd_sc_hd__o211a_1 _18025_ (.A1(_09485_),
    .A2(_09486_),
    .B1(_09345_),
    .C1(_09348_),
    .X(_09488_));
 sky130_fd_sc_hd__nand2_1 _18026_ (.A(_09368_),
    .B(_09370_),
    .Y(_09489_));
 sky130_fd_sc_hd__a21bo_1 _18027_ (.A1(_09377_),
    .A2(_09384_),
    .B1_N(_09383_),
    .X(_09490_));
 sky130_fd_sc_hd__and2_1 _18028_ (.A(net271),
    .B(net129),
    .X(_09491_));
 sky130_fd_sc_hd__a22o_1 _18029_ (.A1(net262),
    .A2(net138),
    .B1(net133),
    .B2(net267),
    .X(_09492_));
 sky130_fd_sc_hd__nand4_1 _18030_ (.A(net262),
    .B(net267),
    .C(net138),
    .D(net133),
    .Y(_09493_));
 sky130_fd_sc_hd__nand2_1 _18031_ (.A(_09492_),
    .B(_09493_),
    .Y(_09494_));
 sky130_fd_sc_hd__xnor2_1 _18032_ (.A(_09491_),
    .B(_09494_),
    .Y(_09495_));
 sky130_fd_sc_hd__nand4_1 _18033_ (.A(net629),
    .B(net249),
    .C(net152),
    .D(net147),
    .Y(_09496_));
 sky130_fd_sc_hd__a22o_1 _18034_ (.A1(net629),
    .A2(net152),
    .B1(net147),
    .B2(net251),
    .X(_09497_));
 sky130_fd_sc_hd__nand4_1 _18035_ (.A(net256),
    .B(net144),
    .C(_09496_),
    .D(_09497_),
    .Y(_09498_));
 sky130_fd_sc_hd__a22o_1 _18036_ (.A1(net256),
    .A2(net144),
    .B1(_09496_),
    .B2(_09497_),
    .X(_09499_));
 sky130_fd_sc_hd__a21bo_1 _18037_ (.A1(_09362_),
    .A2(_09364_),
    .B1_N(_09363_),
    .X(_09500_));
 sky130_fd_sc_hd__nand3_1 _18038_ (.A(_09498_),
    .B(_09499_),
    .C(_09500_),
    .Y(_09501_));
 sky130_fd_sc_hd__a21o_1 _18039_ (.A1(_09498_),
    .A2(_09499_),
    .B1(_09500_),
    .X(_09502_));
 sky130_fd_sc_hd__nand3_2 _18040_ (.A(_09495_),
    .B(_09501_),
    .C(_09502_),
    .Y(_09503_));
 sky130_fd_sc_hd__a21o_1 _18041_ (.A1(_09501_),
    .A2(_09502_),
    .B1(_09495_),
    .X(_09504_));
 sky130_fd_sc_hd__nand3_2 _18042_ (.A(_09490_),
    .B(_09503_),
    .C(_09504_),
    .Y(_09505_));
 sky130_fd_sc_hd__a21o_1 _18043_ (.A1(_09503_),
    .A2(_09504_),
    .B1(_09490_),
    .X(_09506_));
 sky130_fd_sc_hd__nand3_1 _18044_ (.A(_09489_),
    .B(_09505_),
    .C(_09506_),
    .Y(_09507_));
 sky130_fd_sc_hd__a21o_1 _18045_ (.A1(_09505_),
    .A2(_09506_),
    .B1(_09489_),
    .X(_09508_));
 sky130_fd_sc_hd__nand2_1 _18046_ (.A(_09507_),
    .B(_09508_),
    .Y(_09509_));
 sky130_fd_sc_hd__nand2_1 _18047_ (.A(_09379_),
    .B(_09381_),
    .Y(_09510_));
 sky130_fd_sc_hd__o21ba_1 _18048_ (.A1(_09388_),
    .A2(_09390_),
    .B1_N(_09389_),
    .X(_09511_));
 sky130_fd_sc_hd__a22oi_1 _18049_ (.A1(net162),
    .A2(net238),
    .B1(net233),
    .B2(net169),
    .Y(_09512_));
 sky130_fd_sc_hd__and4_1 _18050_ (.A(net169),
    .B(net162),
    .C(net238),
    .D(net233),
    .X(_09513_));
 sky130_fd_sc_hd__and4bb_1 _18051_ (.A_N(_09512_),
    .B_N(_09513_),
    .C(net244),
    .D(net157),
    .X(_09514_));
 sky130_fd_sc_hd__o2bb2a_1 _18052_ (.A1_N(net244),
    .A2_N(net157),
    .B1(_09512_),
    .B2(_09513_),
    .X(_09515_));
 sky130_fd_sc_hd__nor2_1 _18053_ (.A(_09514_),
    .B(_09515_),
    .Y(_09516_));
 sky130_fd_sc_hd__or3_1 _18054_ (.A(_09511_),
    .B(_09514_),
    .C(_09515_),
    .X(_09517_));
 sky130_fd_sc_hd__xnor2_2 _18055_ (.A(_09511_),
    .B(_09516_),
    .Y(_09518_));
 sky130_fd_sc_hd__nand2_1 _18056_ (.A(_09510_),
    .B(_09518_),
    .Y(_09519_));
 sky130_fd_sc_hd__xor2_2 _18057_ (.A(_09510_),
    .B(_09518_),
    .X(_09520_));
 sky130_fd_sc_hd__nand2_1 _18058_ (.A(net175),
    .B(net229),
    .Y(_09521_));
 sky130_fd_sc_hd__and4_1 _18059_ (.A(net184),
    .B(net179),
    .C(net225),
    .D(net219),
    .X(_09522_));
 sky130_fd_sc_hd__a22oi_2 _18060_ (.A1(net179),
    .A2(net225),
    .B1(net219),
    .B2(net184),
    .Y(_09523_));
 sky130_fd_sc_hd__nor2_1 _18061_ (.A(_09522_),
    .B(_09523_),
    .Y(_09524_));
 sky130_fd_sc_hd__xnor2_2 _18062_ (.A(_09521_),
    .B(_09524_),
    .Y(_09525_));
 sky130_fd_sc_hd__and2_1 _18063_ (.A(net187),
    .B(net215),
    .X(_09526_));
 sky130_fd_sc_hd__nand4_2 _18064_ (.A(net624),
    .B(net191),
    .C(net211),
    .D(net208),
    .Y(_09527_));
 sky130_fd_sc_hd__a22o_1 _18065_ (.A1(net191),
    .A2(net211),
    .B1(net208),
    .B2(net624),
    .X(_09528_));
 sky130_fd_sc_hd__nand3_1 _18066_ (.A(_09526_),
    .B(_09527_),
    .C(_09528_),
    .Y(_09529_));
 sky130_fd_sc_hd__a21o_1 _18067_ (.A1(_09527_),
    .A2(_09528_),
    .B1(_09526_),
    .X(_09530_));
 sky130_fd_sc_hd__a21bo_1 _18068_ (.A1(_09393_),
    .A2(_09395_),
    .B1_N(_09394_),
    .X(_09531_));
 sky130_fd_sc_hd__nand3_1 _18069_ (.A(_09529_),
    .B(_09530_),
    .C(_09531_),
    .Y(_09532_));
 sky130_fd_sc_hd__a21o_1 _18070_ (.A1(_09529_),
    .A2(_09530_),
    .B1(_09531_),
    .X(_09533_));
 sky130_fd_sc_hd__nand3_2 _18071_ (.A(_09525_),
    .B(_09532_),
    .C(_09533_),
    .Y(_09534_));
 sky130_fd_sc_hd__a21o_1 _18072_ (.A1(_09532_),
    .A2(_09533_),
    .B1(_09525_),
    .X(_09535_));
 sky130_fd_sc_hd__a21bo_1 _18073_ (.A1(_09392_),
    .A2(_09400_),
    .B1_N(_09399_),
    .X(_09536_));
 sky130_fd_sc_hd__nand3_4 _18074_ (.A(_09534_),
    .B(_09535_),
    .C(_09536_),
    .Y(_09537_));
 sky130_fd_sc_hd__a21o_1 _18075_ (.A1(_09534_),
    .A2(_09535_),
    .B1(_09536_),
    .X(_09538_));
 sky130_fd_sc_hd__and3_1 _18076_ (.A(_09520_),
    .B(_09537_),
    .C(_09538_),
    .X(_09539_));
 sky130_fd_sc_hd__nand3_2 _18077_ (.A(_09520_),
    .B(_09537_),
    .C(_09538_),
    .Y(_09540_));
 sky130_fd_sc_hd__a21oi_2 _18078_ (.A1(_09537_),
    .A2(_09538_),
    .B1(_09520_),
    .Y(_09541_));
 sky130_fd_sc_hd__a211oi_4 _18079_ (.A1(_09404_),
    .A2(_09407_),
    .B1(_09539_),
    .C1(_09541_),
    .Y(_09542_));
 sky130_fd_sc_hd__o211a_1 _18080_ (.A1(_09539_),
    .A2(_09541_),
    .B1(_09404_),
    .C1(_09407_),
    .X(_09543_));
 sky130_fd_sc_hd__nor3_1 _18081_ (.A(_09509_),
    .B(_09542_),
    .C(_09543_),
    .Y(_09544_));
 sky130_fd_sc_hd__or3_2 _18082_ (.A(_09509_),
    .B(_09542_),
    .C(_09543_),
    .X(_09545_));
 sky130_fd_sc_hd__o21ai_2 _18083_ (.A1(_09542_),
    .A2(_09543_),
    .B1(_09509_),
    .Y(_09546_));
 sky130_fd_sc_hd__o211a_2 _18084_ (.A1(_09409_),
    .A2(_09411_),
    .B1(_09545_),
    .C1(_09546_),
    .X(_09547_));
 sky130_fd_sc_hd__a211oi_4 _18085_ (.A1(_09545_),
    .A2(_09546_),
    .B1(_09409_),
    .C1(_09411_),
    .Y(_09548_));
 sky130_fd_sc_hd__nor4_2 _18086_ (.A(_09487_),
    .B(_09488_),
    .C(_09547_),
    .D(_09548_),
    .Y(_09549_));
 sky130_fd_sc_hd__or4_2 _18087_ (.A(_09487_),
    .B(_09488_),
    .C(_09547_),
    .D(_09548_),
    .X(_09550_));
 sky130_fd_sc_hd__o22ai_4 _18088_ (.A1(_09487_),
    .A2(_09488_),
    .B1(_09547_),
    .B2(_09548_),
    .Y(_09551_));
 sky130_fd_sc_hd__o211ai_4 _18089_ (.A1(_09414_),
    .A2(_09416_),
    .B1(_09550_),
    .C1(_09551_),
    .Y(_09552_));
 sky130_fd_sc_hd__a211o_1 _18090_ (.A1(_09550_),
    .A2(_09551_),
    .B1(_09414_),
    .C1(_09416_),
    .X(_09553_));
 sky130_fd_sc_hd__nand3_4 _18091_ (.A(_09453_),
    .B(_09552_),
    .C(_09553_),
    .Y(_09554_));
 sky130_fd_sc_hd__a21o_1 _18092_ (.A1(_09552_),
    .A2(_09553_),
    .B1(_09453_),
    .X(_09555_));
 sky130_fd_sc_hd__o211ai_4 _18093_ (.A1(_09420_),
    .A2(_09422_),
    .B1(_09554_),
    .C1(_09555_),
    .Y(_09556_));
 sky130_fd_sc_hd__a211o_1 _18094_ (.A1(_09554_),
    .A2(_09555_),
    .B1(_09420_),
    .C1(_09422_),
    .X(_09557_));
 sky130_fd_sc_hd__nand3_4 _18095_ (.A(_09315_),
    .B(_09556_),
    .C(_09557_),
    .Y(_09558_));
 sky130_fd_sc_hd__a21o_1 _18096_ (.A1(_09556_),
    .A2(_09557_),
    .B1(_09315_),
    .X(_09559_));
 sky130_fd_sc_hd__o211ai_4 _18097_ (.A1(_09424_),
    .A2(_09426_),
    .B1(_09558_),
    .C1(_09559_),
    .Y(_09560_));
 sky130_fd_sc_hd__a211o_1 _18098_ (.A1(_09558_),
    .A2(_09559_),
    .B1(_09424_),
    .C1(_09426_),
    .X(_09561_));
 sky130_fd_sc_hd__nand2_2 _18099_ (.A(_09560_),
    .B(_09561_),
    .Y(_09562_));
 sky130_fd_sc_hd__xnor2_2 _18100_ (.A(_09429_),
    .B(_09562_),
    .Y(_09563_));
 sky130_fd_sc_hd__xor2_4 _18101_ (.A(_09437_),
    .B(_09563_),
    .X(_09564_));
 sky130_fd_sc_hd__nor2_1 _18102_ (.A(net44),
    .B(_04719_),
    .Y(_09565_));
 sky130_fd_sc_hd__a221o_1 _18103_ (.A1(net709),
    .A2(net7),
    .B1(_09564_),
    .B2(_03050_),
    .C1(_09565_),
    .X(_09566_));
 sky130_fd_sc_hd__mux2_1 _18104_ (.A0(net704),
    .A1(_09566_),
    .S(net3),
    .X(_00307_));
 sky130_fd_sc_hd__a31o_1 _18105_ (.A1(_09179_),
    .A2(_09312_),
    .A3(_09452_),
    .B1(_09451_),
    .X(_09567_));
 sky130_fd_sc_hd__inv_2 _18106_ (.A(_09567_),
    .Y(_09568_));
 sky130_fd_sc_hd__or2_2 _18107_ (.A(_09485_),
    .B(_09487_),
    .X(_09569_));
 sky130_fd_sc_hd__o21ba_1 _18108_ (.A1(_09458_),
    .A2(_09466_),
    .B1_N(_09465_),
    .X(_09570_));
 sky130_fd_sc_hd__a31oi_1 _18109_ (.A1(net316),
    .A2(net85),
    .A3(_09455_),
    .B1(_09454_),
    .Y(_09571_));
 sky130_fd_sc_hd__and4_1 _18110_ (.A(net316),
    .B(\mul1.a[1] ),
    .C(net81),
    .D(net78),
    .X(_09572_));
 sky130_fd_sc_hd__a22oi_1 _18111_ (.A1(net316),
    .A2(net81),
    .B1(net78),
    .B2(\mul1.a[1] ),
    .Y(_09573_));
 sky130_fd_sc_hd__and4bb_1 _18112_ (.A_N(_09572_),
    .B_N(_09573_),
    .C(net324),
    .D(net75),
    .X(_09574_));
 sky130_fd_sc_hd__o2bb2a_1 _18113_ (.A1_N(net324),
    .A2_N(net75),
    .B1(_09572_),
    .B2(_09573_),
    .X(_09575_));
 sky130_fd_sc_hd__nor3_1 _18114_ (.A(_09571_),
    .B(_09574_),
    .C(_09575_),
    .Y(_09576_));
 sky130_fd_sc_hd__o21ai_1 _18115_ (.A1(_09574_),
    .A2(_09575_),
    .B1(_09571_),
    .Y(_09577_));
 sky130_fd_sc_hd__and2b_1 _18116_ (.A_N(_09576_),
    .B(_09577_),
    .X(_09578_));
 sky130_fd_sc_hd__xnor2_1 _18117_ (.A(_09440_),
    .B(_09578_),
    .Y(_09579_));
 sky130_fd_sc_hd__or2_1 _18118_ (.A(_09570_),
    .B(_09579_),
    .X(_09580_));
 sky130_fd_sc_hd__xnor2_1 _18119_ (.A(_09570_),
    .B(_09579_),
    .Y(_09581_));
 sky130_fd_sc_hd__xor2_1 _18120_ (.A(_09442_),
    .B(_09581_),
    .X(_09582_));
 sky130_fd_sc_hd__or2_1 _18121_ (.A(_09307_),
    .B(_09447_),
    .X(_09583_));
 sky130_fd_sc_hd__and3_1 _18122_ (.A(_09445_),
    .B(_09582_),
    .C(_09583_),
    .X(_09584_));
 sky130_fd_sc_hd__a21oi_1 _18123_ (.A1(_09445_),
    .A2(_09583_),
    .B1(_09582_),
    .Y(_09585_));
 sky130_fd_sc_hd__nor2_1 _18124_ (.A(_09584_),
    .B(_09585_),
    .Y(_09586_));
 sky130_fd_sc_hd__nand2_1 _18125_ (.A(_09569_),
    .B(_09586_),
    .Y(_09587_));
 sky130_fd_sc_hd__xor2_2 _18126_ (.A(_09569_),
    .B(_09586_),
    .X(_09588_));
 sky130_fd_sc_hd__and3b_1 _18127_ (.A_N(_09447_),
    .B(_09310_),
    .C(_09445_),
    .X(_09589_));
 sky130_fd_sc_hd__nand2_1 _18128_ (.A(_09588_),
    .B(_09589_),
    .Y(_09590_));
 sky130_fd_sc_hd__xor2_2 _18129_ (.A(_09588_),
    .B(_09589_),
    .X(_09591_));
 sky130_fd_sc_hd__a22o_1 _18130_ (.A1(net301),
    .A2(net93),
    .B1(net89),
    .B2(net306),
    .X(_09592_));
 sky130_fd_sc_hd__and3_1 _18131_ (.A(net301),
    .B(net306),
    .C(net89),
    .X(_09593_));
 sky130_fd_sc_hd__a21bo_1 _18132_ (.A1(net93),
    .A2(_09593_),
    .B1_N(_09592_),
    .X(_09594_));
 sky130_fd_sc_hd__nand2_1 _18133_ (.A(net311),
    .B(net85),
    .Y(_09595_));
 sky130_fd_sc_hd__xnor2_2 _18134_ (.A(_09594_),
    .B(_09595_),
    .Y(_09596_));
 sky130_fd_sc_hd__nand4_1 _18135_ (.A(net286),
    .B(net290),
    .C(net108),
    .D(net103),
    .Y(_09597_));
 sky130_fd_sc_hd__a22o_1 _18136_ (.A1(net286),
    .A2(net108),
    .B1(net103),
    .B2(net290),
    .X(_09598_));
 sky130_fd_sc_hd__nand4_1 _18137_ (.A(net296),
    .B(net99),
    .C(_09597_),
    .D(_09598_),
    .Y(_09599_));
 sky130_fd_sc_hd__a22o_1 _18138_ (.A1(net296),
    .A2(net99),
    .B1(_09597_),
    .B2(_09598_),
    .X(_09600_));
 sky130_fd_sc_hd__a21bo_1 _18139_ (.A1(_09459_),
    .A2(_09461_),
    .B1_N(_09460_),
    .X(_09601_));
 sky130_fd_sc_hd__and3_1 _18140_ (.A(_09599_),
    .B(_09600_),
    .C(_09601_),
    .X(_09602_));
 sky130_fd_sc_hd__a21oi_1 _18141_ (.A1(_09599_),
    .A2(_09600_),
    .B1(_09601_),
    .Y(_09603_));
 sky130_fd_sc_hd__nor2_1 _18142_ (.A(_09602_),
    .B(_09603_),
    .Y(_09604_));
 sky130_fd_sc_hd__xnor2_2 _18143_ (.A(_09596_),
    .B(_09604_),
    .Y(_09605_));
 sky130_fd_sc_hd__nand2_2 _18144_ (.A(_09471_),
    .B(_09473_),
    .Y(_09606_));
 sky130_fd_sc_hd__a21boi_2 _18145_ (.A1(_09491_),
    .A2(_09492_),
    .B1_N(_09493_),
    .Y(_09607_));
 sky130_fd_sc_hd__and4_1 _18146_ (.A(net270),
    .B(net276),
    .C(net124),
    .D(net119),
    .X(_09608_));
 sky130_fd_sc_hd__a22oi_1 _18147_ (.A1(net270),
    .A2(net124),
    .B1(net119),
    .B2(net276),
    .Y(_09609_));
 sky130_fd_sc_hd__and4bb_1 _18148_ (.A_N(_09608_),
    .B_N(_09609_),
    .C(net281),
    .D(net115),
    .X(_09610_));
 sky130_fd_sc_hd__o2bb2a_1 _18149_ (.A1_N(net281),
    .A2_N(net115),
    .B1(_09608_),
    .B2(_09609_),
    .X(_09611_));
 sky130_fd_sc_hd__or3_4 _18150_ (.A(_09607_),
    .B(_09610_),
    .C(_09611_),
    .X(_09612_));
 sky130_fd_sc_hd__o21ai_2 _18151_ (.A1(_09610_),
    .A2(_09611_),
    .B1(_09607_),
    .Y(_09613_));
 sky130_fd_sc_hd__nand3_4 _18152_ (.A(_09606_),
    .B(_09612_),
    .C(_09613_),
    .Y(_09614_));
 sky130_fd_sc_hd__a21o_1 _18153_ (.A1(_09612_),
    .A2(_09613_),
    .B1(_09606_),
    .X(_09615_));
 sky130_fd_sc_hd__a21bo_1 _18154_ (.A1(_09469_),
    .A2(_09476_),
    .B1_N(_09475_),
    .X(_09616_));
 sky130_fd_sc_hd__and3_2 _18155_ (.A(_09614_),
    .B(_09615_),
    .C(_09616_),
    .X(_09617_));
 sky130_fd_sc_hd__a21oi_2 _18156_ (.A1(_09614_),
    .A2(_09615_),
    .B1(_09616_),
    .Y(_09618_));
 sky130_fd_sc_hd__nor3b_4 _18157_ (.A(_09617_),
    .B(_09618_),
    .C_N(_09605_),
    .Y(_09619_));
 sky130_fd_sc_hd__o21ba_1 _18158_ (.A1(_09617_),
    .A2(_09618_),
    .B1_N(_09605_),
    .X(_09620_));
 sky130_fd_sc_hd__a211o_1 _18159_ (.A1(_09505_),
    .A2(_09507_),
    .B1(_09619_),
    .C1(_09620_),
    .X(_09621_));
 sky130_fd_sc_hd__o211ai_1 _18160_ (.A1(_09619_),
    .A2(_09620_),
    .B1(_09505_),
    .C1(_09507_),
    .Y(_09622_));
 sky130_fd_sc_hd__o211ai_1 _18161_ (.A1(_09480_),
    .A2(_09483_),
    .B1(_09621_),
    .C1(_09622_),
    .Y(_09623_));
 sky130_fd_sc_hd__a211o_1 _18162_ (.A1(_09621_),
    .A2(_09622_),
    .B1(_09480_),
    .C1(_09483_),
    .X(_09624_));
 sky130_fd_sc_hd__nand2_1 _18163_ (.A(_09623_),
    .B(_09624_),
    .Y(_09625_));
 sky130_fd_sc_hd__nand2_1 _18164_ (.A(_09501_),
    .B(_09503_),
    .Y(_09626_));
 sky130_fd_sc_hd__a22o_1 _18165_ (.A1(net256),
    .A2(net140),
    .B1(net133),
    .B2(net260),
    .X(_09627_));
 sky130_fd_sc_hd__nand4_2 _18166_ (.A(net257),
    .B(net260),
    .C(net140),
    .D(net133),
    .Y(_09628_));
 sky130_fd_sc_hd__nand4_1 _18167_ (.A(net264),
    .B(net129),
    .C(_09627_),
    .D(_09628_),
    .Y(_09629_));
 sky130_fd_sc_hd__a22o_1 _18168_ (.A1(net264),
    .A2(net129),
    .B1(_09627_),
    .B2(_09628_),
    .X(_09630_));
 sky130_fd_sc_hd__and2_1 _18169_ (.A(_09629_),
    .B(_09630_),
    .X(_09631_));
 sky130_fd_sc_hd__a22oi_1 _18170_ (.A1(net243),
    .A2(net152),
    .B1(net147),
    .B2(net626),
    .Y(_09632_));
 sky130_fd_sc_hd__and4_1 _18171_ (.A(net243),
    .B(net626),
    .C(net152),
    .D(net147),
    .X(_09633_));
 sky130_fd_sc_hd__and4bb_1 _18172_ (.A_N(_09632_),
    .B_N(_09633_),
    .C(net249),
    .D(net144),
    .X(_09634_));
 sky130_fd_sc_hd__o2bb2a_1 _18173_ (.A1_N(net249),
    .A2_N(net144),
    .B1(_09632_),
    .B2(_09633_),
    .X(_09635_));
 sky130_fd_sc_hd__nor2_1 _18174_ (.A(_09634_),
    .B(_09635_),
    .Y(_09636_));
 sky130_fd_sc_hd__and2_1 _18175_ (.A(_09496_),
    .B(_09498_),
    .X(_09637_));
 sky130_fd_sc_hd__and2b_2 _18176_ (.A_N(_09637_),
    .B(_09636_),
    .X(_09638_));
 sky130_fd_sc_hd__xnor2_1 _18177_ (.A(_09636_),
    .B(_09637_),
    .Y(_09639_));
 sky130_fd_sc_hd__and2_2 _18178_ (.A(_09631_),
    .B(_09639_),
    .X(_09640_));
 sky130_fd_sc_hd__xnor2_1 _18179_ (.A(_09631_),
    .B(_09639_),
    .Y(_09641_));
 sky130_fd_sc_hd__a21o_2 _18180_ (.A1(_09517_),
    .A2(_09519_),
    .B1(_09641_),
    .X(_09642_));
 sky130_fd_sc_hd__nand3_2 _18181_ (.A(_09517_),
    .B(_09519_),
    .C(_09641_),
    .Y(_09643_));
 sky130_fd_sc_hd__and3_1 _18182_ (.A(_09626_),
    .B(_09642_),
    .C(_09643_),
    .X(_09644_));
 sky130_fd_sc_hd__nand3_2 _18183_ (.A(_09626_),
    .B(_09642_),
    .C(_09643_),
    .Y(_09645_));
 sky130_fd_sc_hd__a21oi_2 _18184_ (.A1(_09642_),
    .A2(_09643_),
    .B1(_09626_),
    .Y(_09646_));
 sky130_fd_sc_hd__or2_1 _18185_ (.A(_09513_),
    .B(_09514_),
    .X(_09647_));
 sky130_fd_sc_hd__o21ba_1 _18186_ (.A1(_09521_),
    .A2(_09523_),
    .B1_N(_09522_),
    .X(_09648_));
 sky130_fd_sc_hd__a22oi_1 _18187_ (.A1(net162),
    .A2(net233),
    .B1(net228),
    .B2(net169),
    .Y(_09649_));
 sky130_fd_sc_hd__and4_1 _18188_ (.A(net169),
    .B(net162),
    .C(net233),
    .D(net228),
    .X(_09650_));
 sky130_fd_sc_hd__and4bb_1 _18189_ (.A_N(_09649_),
    .B_N(_09650_),
    .C(net157),
    .D(net238),
    .X(_09651_));
 sky130_fd_sc_hd__o2bb2a_1 _18190_ (.A1_N(net157),
    .A2_N(net238),
    .B1(_09649_),
    .B2(_09650_),
    .X(_09652_));
 sky130_fd_sc_hd__nor2_1 _18191_ (.A(_09651_),
    .B(_09652_),
    .Y(_09653_));
 sky130_fd_sc_hd__or3_1 _18192_ (.A(_09648_),
    .B(_09651_),
    .C(_09652_),
    .X(_09654_));
 sky130_fd_sc_hd__xnor2_2 _18193_ (.A(_09648_),
    .B(_09653_),
    .Y(_09655_));
 sky130_fd_sc_hd__nand2_1 _18194_ (.A(_09647_),
    .B(_09655_),
    .Y(_09656_));
 sky130_fd_sc_hd__xor2_2 _18195_ (.A(_09647_),
    .B(_09655_),
    .X(_09657_));
 sky130_fd_sc_hd__nand2_1 _18196_ (.A(net174),
    .B(net225),
    .Y(_09658_));
 sky130_fd_sc_hd__and4_1 _18197_ (.A(net184),
    .B(net179),
    .C(net219),
    .D(net215),
    .X(_09659_));
 sky130_fd_sc_hd__a22o_1 _18198_ (.A1(net179),
    .A2(net219),
    .B1(net216),
    .B2(net184),
    .X(_09660_));
 sky130_fd_sc_hd__and2b_1 _18199_ (.A_N(_09659_),
    .B(_09660_),
    .X(_09661_));
 sky130_fd_sc_hd__xnor2_2 _18200_ (.A(_09658_),
    .B(_09661_),
    .Y(_09662_));
 sky130_fd_sc_hd__and2_1 _18201_ (.A(net187),
    .B(net211),
    .X(_09663_));
 sky130_fd_sc_hd__nand4_2 _18202_ (.A(net624),
    .B(net191),
    .C(net208),
    .D(net205),
    .Y(_09664_));
 sky130_fd_sc_hd__a22o_1 _18203_ (.A1(net191),
    .A2(net208),
    .B1(net205),
    .B2(net624),
    .X(_09665_));
 sky130_fd_sc_hd__nand3_1 _18204_ (.A(_09663_),
    .B(_09664_),
    .C(_09665_),
    .Y(_09666_));
 sky130_fd_sc_hd__a21o_1 _18205_ (.A1(_09664_),
    .A2(_09665_),
    .B1(_09663_),
    .X(_09667_));
 sky130_fd_sc_hd__a21bo_1 _18206_ (.A1(_09526_),
    .A2(_09528_),
    .B1_N(_09527_),
    .X(_09668_));
 sky130_fd_sc_hd__nand3_1 _18207_ (.A(_09666_),
    .B(_09667_),
    .C(_09668_),
    .Y(_09669_));
 sky130_fd_sc_hd__a21o_1 _18208_ (.A1(_09666_),
    .A2(_09667_),
    .B1(_09668_),
    .X(_09670_));
 sky130_fd_sc_hd__nand3_2 _18209_ (.A(_09662_),
    .B(_09669_),
    .C(_09670_),
    .Y(_09671_));
 sky130_fd_sc_hd__a21o_1 _18210_ (.A1(_09669_),
    .A2(_09670_),
    .B1(_09662_),
    .X(_09672_));
 sky130_fd_sc_hd__a21bo_1 _18211_ (.A1(_09525_),
    .A2(_09533_),
    .B1_N(_09532_),
    .X(_09673_));
 sky130_fd_sc_hd__nand3_4 _18212_ (.A(_09671_),
    .B(_09672_),
    .C(_09673_),
    .Y(_09674_));
 sky130_fd_sc_hd__a21o_1 _18213_ (.A1(_09671_),
    .A2(_09672_),
    .B1(_09673_),
    .X(_09675_));
 sky130_fd_sc_hd__and3_1 _18214_ (.A(_09657_),
    .B(_09674_),
    .C(_09675_),
    .X(_09676_));
 sky130_fd_sc_hd__nand3_2 _18215_ (.A(_09657_),
    .B(_09674_),
    .C(_09675_),
    .Y(_09677_));
 sky130_fd_sc_hd__a21oi_2 _18216_ (.A1(_09674_),
    .A2(_09675_),
    .B1(_09657_),
    .Y(_09678_));
 sky130_fd_sc_hd__a211oi_4 _18217_ (.A1(_09537_),
    .A2(_09540_),
    .B1(_09676_),
    .C1(_09678_),
    .Y(_09679_));
 sky130_fd_sc_hd__o211a_1 _18218_ (.A1(_09676_),
    .A2(_09678_),
    .B1(_09537_),
    .C1(_09540_),
    .X(_09680_));
 sky130_fd_sc_hd__nor4_2 _18219_ (.A(_09644_),
    .B(_09646_),
    .C(_09679_),
    .D(_09680_),
    .Y(_09681_));
 sky130_fd_sc_hd__or4_1 _18220_ (.A(_09644_),
    .B(_09646_),
    .C(_09679_),
    .D(_09680_),
    .X(_09682_));
 sky130_fd_sc_hd__o22ai_2 _18221_ (.A1(_09644_),
    .A2(_09646_),
    .B1(_09679_),
    .B2(_09680_),
    .Y(_09683_));
 sky130_fd_sc_hd__o211a_2 _18222_ (.A1(_09542_),
    .A2(_09544_),
    .B1(_09682_),
    .C1(_09683_),
    .X(_09684_));
 sky130_fd_sc_hd__a211oi_2 _18223_ (.A1(_09682_),
    .A2(_09683_),
    .B1(_09542_),
    .C1(_09544_),
    .Y(_09685_));
 sky130_fd_sc_hd__nor3_2 _18224_ (.A(_09625_),
    .B(_09684_),
    .C(_09685_),
    .Y(_09686_));
 sky130_fd_sc_hd__or3_2 _18225_ (.A(_09625_),
    .B(_09684_),
    .C(_09685_),
    .X(_09687_));
 sky130_fd_sc_hd__o21ai_2 _18226_ (.A1(_09684_),
    .A2(_09685_),
    .B1(_09625_),
    .Y(_09688_));
 sky130_fd_sc_hd__o211ai_4 _18227_ (.A1(_09547_),
    .A2(_09549_),
    .B1(_09687_),
    .C1(_09688_),
    .Y(_09689_));
 sky130_fd_sc_hd__a211o_1 _18228_ (.A1(_09687_),
    .A2(_09688_),
    .B1(_09547_),
    .C1(_09549_),
    .X(_09690_));
 sky130_fd_sc_hd__and3_1 _18229_ (.A(_09591_),
    .B(_09689_),
    .C(_09690_),
    .X(_09691_));
 sky130_fd_sc_hd__nand3_2 _18230_ (.A(_09591_),
    .B(_09689_),
    .C(_09690_),
    .Y(_09692_));
 sky130_fd_sc_hd__a21oi_2 _18231_ (.A1(_09689_),
    .A2(_09690_),
    .B1(_09591_),
    .Y(_09693_));
 sky130_fd_sc_hd__a211oi_4 _18232_ (.A1(_09552_),
    .A2(_09554_),
    .B1(_09691_),
    .C1(_09693_),
    .Y(_09694_));
 sky130_fd_sc_hd__o211a_1 _18233_ (.A1(_09691_),
    .A2(_09693_),
    .B1(_09552_),
    .C1(_09554_),
    .X(_09695_));
 sky130_fd_sc_hd__nor3_2 _18234_ (.A(_09568_),
    .B(_09694_),
    .C(_09695_),
    .Y(_09696_));
 sky130_fd_sc_hd__o21a_1 _18235_ (.A1(_09694_),
    .A2(_09695_),
    .B1(_09568_),
    .X(_09697_));
 sky130_fd_sc_hd__a211o_2 _18236_ (.A1(_09556_),
    .A2(_09558_),
    .B1(_09696_),
    .C1(_09697_),
    .X(_09698_));
 sky130_fd_sc_hd__o211a_1 _18237_ (.A1(_09696_),
    .A2(_09697_),
    .B1(_09556_),
    .C1(_09558_),
    .X(_09699_));
 sky130_fd_sc_hd__o211ai_1 _18238_ (.A1(_09696_),
    .A2(_09697_),
    .B1(_09556_),
    .C1(_09558_),
    .Y(_09700_));
 sky130_fd_sc_hd__nand2_2 _18239_ (.A(_09698_),
    .B(_09700_),
    .Y(_09701_));
 sky130_fd_sc_hd__or3b_2 _18240_ (.A(_09699_),
    .B(_09560_),
    .C_N(_09698_),
    .X(_09702_));
 sky130_fd_sc_hd__xnor2_4 _18241_ (.A(_09560_),
    .B(_09701_),
    .Y(_09703_));
 sky130_fd_sc_hd__a21boi_2 _18242_ (.A1(_09292_),
    .A2(_09430_),
    .B1_N(_09429_),
    .Y(_09704_));
 sky130_fd_sc_hd__or2_1 _18243_ (.A(_09431_),
    .B(_09563_),
    .X(_09705_));
 sky130_fd_sc_hd__o22a_2 _18244_ (.A1(_09562_),
    .A2(_09704_),
    .B1(_09705_),
    .B2(_09304_),
    .X(_09706_));
 sky130_fd_sc_hd__xnor2_4 _18245_ (.A(_09703_),
    .B(_09706_),
    .Y(_09707_));
 sky130_fd_sc_hd__o2bb2a_1 _18246_ (.A1_N(\temp[9] ),
    .A2_N(net8),
    .B1(_04862_),
    .B2(net43),
    .X(_09708_));
 sky130_fd_sc_hd__o21ai_1 _18247_ (.A1(_03049_),
    .A2(_09707_),
    .B1(_09708_),
    .Y(_09709_));
 sky130_fd_sc_hd__mux2_1 _18248_ (.A0(net768),
    .A1(_09709_),
    .S(net2),
    .X(_00308_));
 sky130_fd_sc_hd__o21ai_4 _18249_ (.A1(_09703_),
    .A2(_09706_),
    .B1(_09702_),
    .Y(_09710_));
 sky130_fd_sc_hd__nand2_1 _18250_ (.A(_09621_),
    .B(_09623_),
    .Y(_09711_));
 sky130_fd_sc_hd__a21o_1 _18251_ (.A1(_09440_),
    .A2(_09577_),
    .B1(_09576_),
    .X(_09712_));
 sky130_fd_sc_hd__o21ba_1 _18252_ (.A1(_09596_),
    .A2(_09603_),
    .B1_N(_09602_),
    .X(_09713_));
 sky130_fd_sc_hd__or2_1 _18253_ (.A(_09572_),
    .B(_09574_),
    .X(_09714_));
 sky130_fd_sc_hd__a32oi_2 _18254_ (.A1(net311),
    .A2(net85),
    .A3(_09592_),
    .B1(_09593_),
    .B2(net93),
    .Y(_09715_));
 sky130_fd_sc_hd__a22oi_1 _18255_ (.A1(net311),
    .A2(net81),
    .B1(net78),
    .B2(net316),
    .Y(_09716_));
 sky130_fd_sc_hd__and4_1 _18256_ (.A(net311),
    .B(net316),
    .C(net81),
    .D(net78),
    .X(_09717_));
 sky130_fd_sc_hd__o2bb2a_1 _18257_ (.A1_N(net321),
    .A2_N(net75),
    .B1(_09716_),
    .B2(_09717_),
    .X(_09718_));
 sky130_fd_sc_hd__and4bb_1 _18258_ (.A_N(_09716_),
    .B_N(_09717_),
    .C(net321),
    .D(net75),
    .X(_09719_));
 sky130_fd_sc_hd__or2_1 _18259_ (.A(_09718_),
    .B(_09719_),
    .X(_09720_));
 sky130_fd_sc_hd__or2_1 _18260_ (.A(_09715_),
    .B(_09720_),
    .X(_09721_));
 sky130_fd_sc_hd__xor2_1 _18261_ (.A(_09715_),
    .B(_09720_),
    .X(_09722_));
 sky130_fd_sc_hd__nand2_1 _18262_ (.A(_09714_),
    .B(_09722_),
    .Y(_09723_));
 sky130_fd_sc_hd__xnor2_1 _18263_ (.A(_09714_),
    .B(_09722_),
    .Y(_09724_));
 sky130_fd_sc_hd__or2_1 _18264_ (.A(_09713_),
    .B(_09724_),
    .X(_09725_));
 sky130_fd_sc_hd__xor2_1 _18265_ (.A(_09713_),
    .B(_09724_),
    .X(_09726_));
 sky130_fd_sc_hd__nand2_1 _18266_ (.A(_09712_),
    .B(_09726_),
    .Y(_09727_));
 sky130_fd_sc_hd__xor2_1 _18267_ (.A(_09712_),
    .B(_09726_),
    .X(_09728_));
 sky130_fd_sc_hd__o21ai_1 _18268_ (.A1(_09442_),
    .A2(_09581_),
    .B1(_09580_),
    .Y(_09729_));
 sky130_fd_sc_hd__nand2_1 _18269_ (.A(_09728_),
    .B(_09729_),
    .Y(_09730_));
 sky130_fd_sc_hd__xnor2_1 _18270_ (.A(_09728_),
    .B(_09729_),
    .Y(_09731_));
 sky130_fd_sc_hd__nand2_1 _18271_ (.A(net324),
    .B(net74),
    .Y(_09732_));
 sky130_fd_sc_hd__or2_1 _18272_ (.A(_09731_),
    .B(_09732_),
    .X(_09733_));
 sky130_fd_sc_hd__xnor2_1 _18273_ (.A(_09731_),
    .B(_09732_),
    .Y(_09734_));
 sky130_fd_sc_hd__and2b_1 _18274_ (.A_N(_09734_),
    .B(_09711_),
    .X(_09735_));
 sky130_fd_sc_hd__xnor2_1 _18275_ (.A(_09711_),
    .B(_09734_),
    .Y(_09736_));
 sky130_fd_sc_hd__and2_1 _18276_ (.A(_09584_),
    .B(_09736_),
    .X(_09737_));
 sky130_fd_sc_hd__nor2_1 _18277_ (.A(_09584_),
    .B(_09736_),
    .Y(_09738_));
 sky130_fd_sc_hd__a22o_1 _18278_ (.A1(net296),
    .A2(net93),
    .B1(net89),
    .B2(net301),
    .X(_09739_));
 sky130_fd_sc_hd__nand4_2 _18279_ (.A(net296),
    .B(net301),
    .C(net93),
    .D(net89),
    .Y(_09740_));
 sky130_fd_sc_hd__a22o_1 _18280_ (.A1(net306),
    .A2(net85),
    .B1(_09739_),
    .B2(_09740_),
    .X(_09741_));
 sky130_fd_sc_hd__nand4_2 _18281_ (.A(net306),
    .B(net85),
    .C(_09739_),
    .D(_09740_),
    .Y(_09742_));
 sky130_fd_sc_hd__nand2_1 _18282_ (.A(_09741_),
    .B(_09742_),
    .Y(_09743_));
 sky130_fd_sc_hd__nand2_1 _18283_ (.A(net290),
    .B(net99),
    .Y(_09744_));
 sky130_fd_sc_hd__a22o_1 _18284_ (.A1(net281),
    .A2(net108),
    .B1(net103),
    .B2(net286),
    .X(_09745_));
 sky130_fd_sc_hd__nand4_1 _18285_ (.A(net281),
    .B(net286),
    .C(net108),
    .D(net103),
    .Y(_09746_));
 sky130_fd_sc_hd__nand2_1 _18286_ (.A(_09745_),
    .B(_09746_),
    .Y(_09747_));
 sky130_fd_sc_hd__xor2_2 _18287_ (.A(_09744_),
    .B(_09747_),
    .X(_09748_));
 sky130_fd_sc_hd__and2_1 _18288_ (.A(_09597_),
    .B(_09599_),
    .X(_09749_));
 sky130_fd_sc_hd__nand2b_1 _18289_ (.A_N(_09749_),
    .B(_09748_),
    .Y(_09750_));
 sky130_fd_sc_hd__xnor2_2 _18290_ (.A(_09748_),
    .B(_09749_),
    .Y(_09751_));
 sky130_fd_sc_hd__nand2b_1 _18291_ (.A_N(_09743_),
    .B(_09751_),
    .Y(_09752_));
 sky130_fd_sc_hd__xnor2_2 _18292_ (.A(_09743_),
    .B(_09751_),
    .Y(_09753_));
 sky130_fd_sc_hd__or2_1 _18293_ (.A(_09608_),
    .B(_09610_),
    .X(_09754_));
 sky130_fd_sc_hd__a22oi_1 _18294_ (.A1(net264),
    .A2(net124),
    .B1(net119),
    .B2(net270),
    .Y(_09755_));
 sky130_fd_sc_hd__and4_1 _18295_ (.A(net264),
    .B(net270),
    .C(net124),
    .D(net119),
    .X(_09756_));
 sky130_fd_sc_hd__o2bb2a_1 _18296_ (.A1_N(net276),
    .A2_N(net115),
    .B1(_09755_),
    .B2(_09756_),
    .X(_09757_));
 sky130_fd_sc_hd__and4bb_1 _18297_ (.A_N(_09755_),
    .B_N(_09756_),
    .C(net276),
    .D(net115),
    .X(_09758_));
 sky130_fd_sc_hd__a211o_1 _18298_ (.A1(_09628_),
    .A2(_09629_),
    .B1(_09757_),
    .C1(_09758_),
    .X(_09759_));
 sky130_fd_sc_hd__o211ai_1 _18299_ (.A1(_09757_),
    .A2(_09758_),
    .B1(_09628_),
    .C1(_09629_),
    .Y(_09760_));
 sky130_fd_sc_hd__and2_1 _18300_ (.A(_09759_),
    .B(_09760_),
    .X(_09761_));
 sky130_fd_sc_hd__nand2_1 _18301_ (.A(_09754_),
    .B(_09761_),
    .Y(_09762_));
 sky130_fd_sc_hd__xnor2_2 _18302_ (.A(_09754_),
    .B(_09761_),
    .Y(_09763_));
 sky130_fd_sc_hd__a21oi_4 _18303_ (.A1(_09612_),
    .A2(_09614_),
    .B1(_09763_),
    .Y(_09764_));
 sky130_fd_sc_hd__and3_1 _18304_ (.A(_09612_),
    .B(_09614_),
    .C(_09763_),
    .X(_09765_));
 sky130_fd_sc_hd__nor3b_4 _18305_ (.A(_09764_),
    .B(_09765_),
    .C_N(_09753_),
    .Y(_09766_));
 sky130_fd_sc_hd__o21ba_1 _18306_ (.A1(_09764_),
    .A2(_09765_),
    .B1_N(_09753_),
    .X(_09767_));
 sky130_fd_sc_hd__a211o_2 _18307_ (.A1(_09642_),
    .A2(_09645_),
    .B1(_09766_),
    .C1(_09767_),
    .X(_09768_));
 sky130_fd_sc_hd__o211ai_4 _18308_ (.A1(_09766_),
    .A2(_09767_),
    .B1(_09642_),
    .C1(_09645_),
    .Y(_09769_));
 sky130_fd_sc_hd__o211a_1 _18309_ (.A1(_09617_),
    .A2(_09619_),
    .B1(_09768_),
    .C1(_09769_),
    .X(_09770_));
 sky130_fd_sc_hd__o211ai_2 _18310_ (.A1(_09617_),
    .A2(_09619_),
    .B1(_09768_),
    .C1(_09769_),
    .Y(_09771_));
 sky130_fd_sc_hd__a211oi_2 _18311_ (.A1(_09768_),
    .A2(_09769_),
    .B1(_09617_),
    .C1(_09619_),
    .Y(_09772_));
 sky130_fd_sc_hd__a22o_1 _18312_ (.A1(net248),
    .A2(net140),
    .B1(net133),
    .B2(net253),
    .X(_09773_));
 sky130_fd_sc_hd__nand4_2 _18313_ (.A(net248),
    .B(net253),
    .C(net140),
    .D(net133),
    .Y(_09774_));
 sky130_fd_sc_hd__nand4_2 _18314_ (.A(net259),
    .B(net129),
    .C(_09773_),
    .D(_09774_),
    .Y(_09775_));
 sky130_fd_sc_hd__a22o_1 _18315_ (.A1(net259),
    .A2(net129),
    .B1(_09773_),
    .B2(_09774_),
    .X(_09776_));
 sky130_fd_sc_hd__and2_1 _18316_ (.A(_09775_),
    .B(_09776_),
    .X(_09777_));
 sky130_fd_sc_hd__nand2_1 _18317_ (.A(net626),
    .B(net144),
    .Y(_09778_));
 sky130_fd_sc_hd__a22o_1 _18318_ (.A1(net243),
    .A2(net147),
    .B1(net238),
    .B2(net152),
    .X(_09779_));
 sky130_fd_sc_hd__nand4_1 _18319_ (.A(net243),
    .B(net152),
    .C(net147),
    .D(net238),
    .Y(_09780_));
 sky130_fd_sc_hd__nand2_1 _18320_ (.A(_09779_),
    .B(_09780_),
    .Y(_09781_));
 sky130_fd_sc_hd__xor2_1 _18321_ (.A(_09778_),
    .B(_09781_),
    .X(_09782_));
 sky130_fd_sc_hd__or2_1 _18322_ (.A(_09633_),
    .B(_09634_),
    .X(_09783_));
 sky130_fd_sc_hd__and2_1 _18323_ (.A(_09782_),
    .B(_09783_),
    .X(_09784_));
 sky130_fd_sc_hd__xor2_1 _18324_ (.A(_09782_),
    .B(_09783_),
    .X(_09785_));
 sky130_fd_sc_hd__and2_1 _18325_ (.A(_09777_),
    .B(_09785_),
    .X(_09786_));
 sky130_fd_sc_hd__xnor2_1 _18326_ (.A(_09777_),
    .B(_09785_),
    .Y(_09787_));
 sky130_fd_sc_hd__a21o_2 _18327_ (.A1(_09654_),
    .A2(_09656_),
    .B1(_09787_),
    .X(_09788_));
 sky130_fd_sc_hd__nand3_2 _18328_ (.A(_09654_),
    .B(_09656_),
    .C(_09787_),
    .Y(_09789_));
 sky130_fd_sc_hd__o211a_1 _18329_ (.A1(_09638_),
    .A2(_09640_),
    .B1(_09788_),
    .C1(_09789_),
    .X(_09790_));
 sky130_fd_sc_hd__o211ai_4 _18330_ (.A1(_09638_),
    .A2(_09640_),
    .B1(_09788_),
    .C1(_09789_),
    .Y(_09791_));
 sky130_fd_sc_hd__a211oi_2 _18331_ (.A1(_09788_),
    .A2(_09789_),
    .B1(_09638_),
    .C1(_09640_),
    .Y(_09792_));
 sky130_fd_sc_hd__or2_1 _18332_ (.A(_09650_),
    .B(_09651_),
    .X(_09793_));
 sky130_fd_sc_hd__a31o_1 _18333_ (.A1(net174),
    .A2(net225),
    .A3(_09660_),
    .B1(_09659_),
    .X(_09794_));
 sky130_fd_sc_hd__a22o_1 _18334_ (.A1(net162),
    .A2(net228),
    .B1(net224),
    .B2(net169),
    .X(_09795_));
 sky130_fd_sc_hd__and4_1 _18335_ (.A(net169),
    .B(net162),
    .C(net228),
    .D(net224),
    .X(_09796_));
 sky130_fd_sc_hd__nand4_1 _18336_ (.A(net170),
    .B(net163),
    .C(net228),
    .D(net224),
    .Y(_09797_));
 sky130_fd_sc_hd__a22oi_1 _18337_ (.A1(net157),
    .A2(net233),
    .B1(_09795_),
    .B2(_09797_),
    .Y(_09798_));
 sky130_fd_sc_hd__and4_1 _18338_ (.A(net157),
    .B(net233),
    .C(_09795_),
    .D(_09797_),
    .X(_09799_));
 sky130_fd_sc_hd__or2_1 _18339_ (.A(_09798_),
    .B(_09799_),
    .X(_09800_));
 sky130_fd_sc_hd__and2b_1 _18340_ (.A_N(_09800_),
    .B(_09794_),
    .X(_09801_));
 sky130_fd_sc_hd__xnor2_2 _18341_ (.A(_09794_),
    .B(_09800_),
    .Y(_09802_));
 sky130_fd_sc_hd__and2_1 _18342_ (.A(_09793_),
    .B(_09802_),
    .X(_09803_));
 sky130_fd_sc_hd__xor2_2 _18343_ (.A(_09793_),
    .B(_09802_),
    .X(_09804_));
 sky130_fd_sc_hd__nand2_1 _18344_ (.A(net174),
    .B(net219),
    .Y(_09805_));
 sky130_fd_sc_hd__and4_1 _18345_ (.A(net184),
    .B(net179),
    .C(net215),
    .D(net211),
    .X(_09806_));
 sky130_fd_sc_hd__a22o_1 _18346_ (.A1(net179),
    .A2(net216),
    .B1(net211),
    .B2(net184),
    .X(_09807_));
 sky130_fd_sc_hd__and2b_1 _18347_ (.A_N(_09806_),
    .B(_09807_),
    .X(_09808_));
 sky130_fd_sc_hd__xnor2_2 _18348_ (.A(_09805_),
    .B(_09808_),
    .Y(_09809_));
 sky130_fd_sc_hd__and2_1 _18349_ (.A(net187),
    .B(net208),
    .X(_09810_));
 sky130_fd_sc_hd__nand4_2 _18350_ (.A(net624),
    .B(net191),
    .C(net205),
    .D(net203),
    .Y(_09811_));
 sky130_fd_sc_hd__a22o_1 _18351_ (.A1(net191),
    .A2(net205),
    .B1(net203),
    .B2(net624),
    .X(_09812_));
 sky130_fd_sc_hd__nand3_1 _18352_ (.A(_09810_),
    .B(_09811_),
    .C(_09812_),
    .Y(_09813_));
 sky130_fd_sc_hd__a21o_1 _18353_ (.A1(_09811_),
    .A2(_09812_),
    .B1(_09810_),
    .X(_09814_));
 sky130_fd_sc_hd__a21bo_1 _18354_ (.A1(_09663_),
    .A2(_09665_),
    .B1_N(_09664_),
    .X(_09815_));
 sky130_fd_sc_hd__nand3_2 _18355_ (.A(_09813_),
    .B(_09814_),
    .C(_09815_),
    .Y(_09816_));
 sky130_fd_sc_hd__a21o_1 _18356_ (.A1(_09813_),
    .A2(_09814_),
    .B1(_09815_),
    .X(_09817_));
 sky130_fd_sc_hd__nand3_2 _18357_ (.A(_09809_),
    .B(_09816_),
    .C(_09817_),
    .Y(_09818_));
 sky130_fd_sc_hd__a21o_1 _18358_ (.A1(_09816_),
    .A2(_09817_),
    .B1(_09809_),
    .X(_09819_));
 sky130_fd_sc_hd__a21bo_1 _18359_ (.A1(_09662_),
    .A2(_09670_),
    .B1_N(_09669_),
    .X(_09820_));
 sky130_fd_sc_hd__nand3_4 _18360_ (.A(_09818_),
    .B(_09819_),
    .C(_09820_),
    .Y(_09821_));
 sky130_fd_sc_hd__a21o_1 _18361_ (.A1(_09818_),
    .A2(_09819_),
    .B1(_09820_),
    .X(_09822_));
 sky130_fd_sc_hd__and3_1 _18362_ (.A(_09804_),
    .B(_09821_),
    .C(_09822_),
    .X(_09823_));
 sky130_fd_sc_hd__nand3_2 _18363_ (.A(_09804_),
    .B(_09821_),
    .C(_09822_),
    .Y(_09824_));
 sky130_fd_sc_hd__a21oi_2 _18364_ (.A1(_09821_),
    .A2(_09822_),
    .B1(_09804_),
    .Y(_09825_));
 sky130_fd_sc_hd__a211oi_4 _18365_ (.A1(_09674_),
    .A2(_09677_),
    .B1(_09823_),
    .C1(_09825_),
    .Y(_09826_));
 sky130_fd_sc_hd__o211a_1 _18366_ (.A1(_09823_),
    .A2(_09825_),
    .B1(_09674_),
    .C1(_09677_),
    .X(_09827_));
 sky130_fd_sc_hd__nor4_1 _18367_ (.A(_09790_),
    .B(_09792_),
    .C(_09826_),
    .D(_09827_),
    .Y(_09828_));
 sky130_fd_sc_hd__or4_1 _18368_ (.A(_09790_),
    .B(_09792_),
    .C(_09826_),
    .D(_09827_),
    .X(_09829_));
 sky130_fd_sc_hd__o22ai_2 _18369_ (.A1(_09790_),
    .A2(_09792_),
    .B1(_09826_),
    .B2(_09827_),
    .Y(_09830_));
 sky130_fd_sc_hd__o211a_2 _18370_ (.A1(_09679_),
    .A2(_09681_),
    .B1(_09829_),
    .C1(_09830_),
    .X(_09831_));
 sky130_fd_sc_hd__a211oi_2 _18371_ (.A1(_09829_),
    .A2(_09830_),
    .B1(_09679_),
    .C1(_09681_),
    .Y(_09832_));
 sky130_fd_sc_hd__nor4_1 _18372_ (.A(_09770_),
    .B(_09772_),
    .C(_09831_),
    .D(_09832_),
    .Y(_09833_));
 sky130_fd_sc_hd__or4_2 _18373_ (.A(_09770_),
    .B(_09772_),
    .C(_09831_),
    .D(_09832_),
    .X(_09834_));
 sky130_fd_sc_hd__o22ai_4 _18374_ (.A1(_09770_),
    .A2(_09772_),
    .B1(_09831_),
    .B2(_09832_),
    .Y(_09835_));
 sky130_fd_sc_hd__o211ai_4 _18375_ (.A1(_09684_),
    .A2(_09686_),
    .B1(_09834_),
    .C1(_09835_),
    .Y(_09836_));
 sky130_fd_sc_hd__a211o_1 _18376_ (.A1(_09834_),
    .A2(_09835_),
    .B1(_09684_),
    .C1(_09686_),
    .X(_09837_));
 sky130_fd_sc_hd__and4bb_1 _18377_ (.A_N(_09737_),
    .B_N(_09738_),
    .C(_09836_),
    .D(_09837_),
    .X(_09838_));
 sky130_fd_sc_hd__or4bb_1 _18378_ (.A(_09737_),
    .B(_09738_),
    .C_N(_09836_),
    .D_N(_09837_),
    .X(_09839_));
 sky130_fd_sc_hd__a2bb2oi_2 _18379_ (.A1_N(_09737_),
    .A2_N(_09738_),
    .B1(_09836_),
    .B2(_09837_),
    .Y(_09840_));
 sky130_fd_sc_hd__a211oi_4 _18380_ (.A1(_09689_),
    .A2(_09692_),
    .B1(_09838_),
    .C1(_09840_),
    .Y(_09841_));
 sky130_fd_sc_hd__o211a_1 _18381_ (.A1(_09838_),
    .A2(_09840_),
    .B1(_09689_),
    .C1(_09692_),
    .X(_09842_));
 sky130_fd_sc_hd__a211oi_2 _18382_ (.A1(_09587_),
    .A2(_09590_),
    .B1(_09841_),
    .C1(_09842_),
    .Y(_09843_));
 sky130_fd_sc_hd__a211o_1 _18383_ (.A1(_09587_),
    .A2(_09590_),
    .B1(_09841_),
    .C1(_09842_),
    .X(_09844_));
 sky130_fd_sc_hd__o211ai_2 _18384_ (.A1(_09841_),
    .A2(_09842_),
    .B1(_09587_),
    .C1(_09590_),
    .Y(_09845_));
 sky130_fd_sc_hd__nand2_2 _18385_ (.A(_09844_),
    .B(_09845_),
    .Y(_09846_));
 sky130_fd_sc_hd__nor2_2 _18386_ (.A(_09694_),
    .B(_09696_),
    .Y(_09847_));
 sky130_fd_sc_hd__o211a_1 _18387_ (.A1(_09694_),
    .A2(_09696_),
    .B1(_09844_),
    .C1(_09845_),
    .X(_09848_));
 sky130_fd_sc_hd__xor2_4 _18388_ (.A(_09846_),
    .B(_09847_),
    .X(_09849_));
 sky130_fd_sc_hd__xor2_4 _18389_ (.A(_09698_),
    .B(_09849_),
    .X(_09850_));
 sky130_fd_sc_hd__xnor2_4 _18390_ (.A(_09710_),
    .B(_09850_),
    .Y(_09851_));
 sky130_fd_sc_hd__nor2_1 _18391_ (.A(net43),
    .B(_05006_),
    .Y(_09852_));
 sky130_fd_sc_hd__a221o_1 _18392_ (.A1(\temp[10] ),
    .A2(net8),
    .B1(_09851_),
    .B2(net10),
    .C1(_09852_),
    .X(_09853_));
 sky130_fd_sc_hd__mux2_1 _18393_ (.A0(net680),
    .A1(_09853_),
    .S(net2),
    .X(_00309_));
 sky130_fd_sc_hd__nor3_2 _18394_ (.A(_09703_),
    .B(_09705_),
    .C(_09850_),
    .Y(_09854_));
 sky130_fd_sc_hd__a21bo_1 _18395_ (.A1(_09698_),
    .A2(_09702_),
    .B1_N(_09849_),
    .X(_09855_));
 sky130_fd_sc_hd__o41ai_4 _18396_ (.A1(_09562_),
    .A2(_09703_),
    .A3(_09704_),
    .A4(_09850_),
    .B1(_09855_),
    .Y(_09856_));
 sky130_fd_sc_hd__a21oi_4 _18397_ (.A1(_09305_),
    .A2(_09854_),
    .B1(_09856_),
    .Y(_09857_));
 sky130_fd_sc_hd__nor2_1 _18398_ (.A(_09735_),
    .B(_09737_),
    .Y(_09858_));
 sky130_fd_sc_hd__a22oi_2 _18399_ (.A1(\mul1.a[1] ),
    .A2(net74),
    .B1(net71),
    .B2(net324),
    .Y(_09859_));
 sky130_fd_sc_hd__and4_1 _18400_ (.A(\mul1.a[1] ),
    .B(net324),
    .C(net74),
    .D(net71),
    .X(_09860_));
 sky130_fd_sc_hd__inv_2 _18401_ (.A(_09860_),
    .Y(_09861_));
 sky130_fd_sc_hd__or2_1 _18402_ (.A(_09717_),
    .B(_09719_),
    .X(_09862_));
 sky130_fd_sc_hd__a22oi_1 _18403_ (.A1(net306),
    .A2(net81),
    .B1(net78),
    .B2(net311),
    .Y(_09863_));
 sky130_fd_sc_hd__and4_1 _18404_ (.A(net306),
    .B(net311),
    .C(net81),
    .D(net78),
    .X(_09864_));
 sky130_fd_sc_hd__o2bb2a_1 _18405_ (.A1_N(net316),
    .A2_N(net75),
    .B1(_09863_),
    .B2(_09864_),
    .X(_09865_));
 sky130_fd_sc_hd__and4bb_1 _18406_ (.A_N(_09863_),
    .B_N(_09864_),
    .C(net316),
    .D(net75),
    .X(_09866_));
 sky130_fd_sc_hd__a211o_1 _18407_ (.A1(_09740_),
    .A2(_09742_),
    .B1(_09865_),
    .C1(_09866_),
    .X(_09867_));
 sky130_fd_sc_hd__o211ai_1 _18408_ (.A1(_09865_),
    .A2(_09866_),
    .B1(_09740_),
    .C1(_09742_),
    .Y(_09868_));
 sky130_fd_sc_hd__and2_1 _18409_ (.A(_09867_),
    .B(_09868_),
    .X(_09869_));
 sky130_fd_sc_hd__nand2_1 _18410_ (.A(_09862_),
    .B(_09869_),
    .Y(_09870_));
 sky130_fd_sc_hd__xnor2_1 _18411_ (.A(_09862_),
    .B(_09869_),
    .Y(_09871_));
 sky130_fd_sc_hd__a21oi_2 _18412_ (.A1(_09750_),
    .A2(_09752_),
    .B1(_09871_),
    .Y(_09872_));
 sky130_fd_sc_hd__inv_2 _18413_ (.A(_09872_),
    .Y(_09873_));
 sky130_fd_sc_hd__and3_1 _18414_ (.A(_09750_),
    .B(_09752_),
    .C(_09871_),
    .X(_09874_));
 sky130_fd_sc_hd__a211oi_2 _18415_ (.A1(_09721_),
    .A2(_09723_),
    .B1(_09872_),
    .C1(_09874_),
    .Y(_09875_));
 sky130_fd_sc_hd__a211o_1 _18416_ (.A1(_09721_),
    .A2(_09723_),
    .B1(_09872_),
    .C1(_09874_),
    .X(_09876_));
 sky130_fd_sc_hd__o211a_1 _18417_ (.A1(_09872_),
    .A2(_09874_),
    .B1(_09721_),
    .C1(_09723_),
    .X(_09877_));
 sky130_fd_sc_hd__a211oi_2 _18418_ (.A1(_09725_),
    .A2(_09727_),
    .B1(_09875_),
    .C1(_09877_),
    .Y(_09878_));
 sky130_fd_sc_hd__o211a_1 _18419_ (.A1(_09875_),
    .A2(_09877_),
    .B1(_09725_),
    .C1(_09727_),
    .X(_09879_));
 sky130_fd_sc_hd__nor4_2 _18420_ (.A(_09859_),
    .B(_09860_),
    .C(_09878_),
    .D(_09879_),
    .Y(_09880_));
 sky130_fd_sc_hd__o22a_1 _18421_ (.A1(_09859_),
    .A2(_09860_),
    .B1(_09878_),
    .B2(_09879_),
    .X(_09881_));
 sky130_fd_sc_hd__a211oi_2 _18422_ (.A1(_09768_),
    .A2(_09771_),
    .B1(_09880_),
    .C1(_09881_),
    .Y(_09882_));
 sky130_fd_sc_hd__o211a_1 _18423_ (.A1(_09880_),
    .A2(_09881_),
    .B1(_09768_),
    .C1(_09771_),
    .X(_09883_));
 sky130_fd_sc_hd__a211oi_2 _18424_ (.A1(_09730_),
    .A2(_09733_),
    .B1(_09882_),
    .C1(_09883_),
    .Y(_09884_));
 sky130_fd_sc_hd__o211a_1 _18425_ (.A1(_09882_),
    .A2(_09883_),
    .B1(_09730_),
    .C1(_09733_),
    .X(_09885_));
 sky130_fd_sc_hd__a22o_1 _18426_ (.A1(net290),
    .A2(net93),
    .B1(net89),
    .B2(net296),
    .X(_09886_));
 sky130_fd_sc_hd__nand4_2 _18427_ (.A(net290),
    .B(net296),
    .C(net93),
    .D(net89),
    .Y(_09887_));
 sky130_fd_sc_hd__a22o_1 _18428_ (.A1(net301),
    .A2(net85),
    .B1(_09886_),
    .B2(_09887_),
    .X(_09888_));
 sky130_fd_sc_hd__nand4_2 _18429_ (.A(net301),
    .B(net85),
    .C(_09886_),
    .D(_09887_),
    .Y(_09889_));
 sky130_fd_sc_hd__nand2_1 _18430_ (.A(_09888_),
    .B(_09889_),
    .Y(_09890_));
 sky130_fd_sc_hd__a22oi_1 _18431_ (.A1(net276),
    .A2(net108),
    .B1(net103),
    .B2(net281),
    .Y(_09891_));
 sky130_fd_sc_hd__and4_1 _18432_ (.A(net276),
    .B(net281),
    .C(net108),
    .D(net103),
    .X(_09892_));
 sky130_fd_sc_hd__o2bb2a_1 _18433_ (.A1_N(net286),
    .A2_N(net99),
    .B1(_09891_),
    .B2(_09892_),
    .X(_09893_));
 sky130_fd_sc_hd__and4bb_1 _18434_ (.A_N(_09891_),
    .B_N(_09892_),
    .C(net286),
    .D(net99),
    .X(_09894_));
 sky130_fd_sc_hd__or2_1 _18435_ (.A(_09893_),
    .B(_09894_),
    .X(_09895_));
 sky130_fd_sc_hd__o21ai_1 _18436_ (.A1(_09744_),
    .A2(_09747_),
    .B1(_09746_),
    .Y(_09896_));
 sky130_fd_sc_hd__nand2b_1 _18437_ (.A_N(_09895_),
    .B(_09896_),
    .Y(_09897_));
 sky130_fd_sc_hd__xor2_1 _18438_ (.A(_09895_),
    .B(_09896_),
    .X(_09898_));
 sky130_fd_sc_hd__or2_1 _18439_ (.A(_09890_),
    .B(_09898_),
    .X(_09899_));
 sky130_fd_sc_hd__nand2_1 _18440_ (.A(_09890_),
    .B(_09898_),
    .Y(_09900_));
 sky130_fd_sc_hd__and2_1 _18441_ (.A(_09899_),
    .B(_09900_),
    .X(_09901_));
 sky130_fd_sc_hd__or2_1 _18442_ (.A(_09756_),
    .B(_09758_),
    .X(_09902_));
 sky130_fd_sc_hd__a22oi_1 _18443_ (.A1(net259),
    .A2(net124),
    .B1(net119),
    .B2(net264),
    .Y(_09903_));
 sky130_fd_sc_hd__and4_1 _18444_ (.A(net259),
    .B(net266),
    .C(net124),
    .D(net119),
    .X(_09904_));
 sky130_fd_sc_hd__o2bb2a_1 _18445_ (.A1_N(net270),
    .A2_N(net115),
    .B1(_09903_),
    .B2(_09904_),
    .X(_09905_));
 sky130_fd_sc_hd__and4bb_1 _18446_ (.A_N(_09903_),
    .B_N(_09904_),
    .C(net270),
    .D(net115),
    .X(_09906_));
 sky130_fd_sc_hd__a211o_1 _18447_ (.A1(_09774_),
    .A2(_09775_),
    .B1(_09905_),
    .C1(_09906_),
    .X(_09907_));
 sky130_fd_sc_hd__o211ai_1 _18448_ (.A1(_09905_),
    .A2(_09906_),
    .B1(_09774_),
    .C1(_09775_),
    .Y(_09908_));
 sky130_fd_sc_hd__and2_1 _18449_ (.A(_09907_),
    .B(_09908_),
    .X(_09909_));
 sky130_fd_sc_hd__nand2_1 _18450_ (.A(_09902_),
    .B(_09909_),
    .Y(_09910_));
 sky130_fd_sc_hd__xnor2_2 _18451_ (.A(_09902_),
    .B(_09909_),
    .Y(_09911_));
 sky130_fd_sc_hd__a21oi_4 _18452_ (.A1(_09759_),
    .A2(_09762_),
    .B1(_09911_),
    .Y(_09912_));
 sky130_fd_sc_hd__and3_1 _18453_ (.A(_09759_),
    .B(_09762_),
    .C(_09911_),
    .X(_09913_));
 sky130_fd_sc_hd__nor3b_4 _18454_ (.A(_09912_),
    .B(_09913_),
    .C_N(_09901_),
    .Y(_09914_));
 sky130_fd_sc_hd__o21ba_1 _18455_ (.A1(_09912_),
    .A2(_09913_),
    .B1_N(_09901_),
    .X(_09915_));
 sky130_fd_sc_hd__a211o_2 _18456_ (.A1(_09788_),
    .A2(_09791_),
    .B1(_09914_),
    .C1(_09915_),
    .X(_09916_));
 sky130_fd_sc_hd__o211ai_4 _18457_ (.A1(_09914_),
    .A2(_09915_),
    .B1(_09788_),
    .C1(_09791_),
    .Y(_09917_));
 sky130_fd_sc_hd__o211a_1 _18458_ (.A1(_09764_),
    .A2(_09766_),
    .B1(_09916_),
    .C1(_09917_),
    .X(_09918_));
 sky130_fd_sc_hd__o211ai_2 _18459_ (.A1(_09764_),
    .A2(_09766_),
    .B1(_09916_),
    .C1(_09917_),
    .Y(_09919_));
 sky130_fd_sc_hd__a211oi_2 _18460_ (.A1(_09916_),
    .A2(_09917_),
    .B1(_09764_),
    .C1(_09766_),
    .Y(_09920_));
 sky130_fd_sc_hd__a22o_1 _18461_ (.A1(net626),
    .A2(net140),
    .B1(net133),
    .B2(net248),
    .X(_09921_));
 sky130_fd_sc_hd__nand4_4 _18462_ (.A(net626),
    .B(net248),
    .C(net138),
    .D(net133),
    .Y(_09922_));
 sky130_fd_sc_hd__a22o_1 _18463_ (.A1(net253),
    .A2(net129),
    .B1(_09921_),
    .B2(_09922_),
    .X(_09923_));
 sky130_fd_sc_hd__nand4_2 _18464_ (.A(net253),
    .B(net129),
    .C(_09921_),
    .D(_09922_),
    .Y(_09924_));
 sky130_fd_sc_hd__nand2_1 _18465_ (.A(_09923_),
    .B(_09924_),
    .Y(_09925_));
 sky130_fd_sc_hd__a22oi_1 _18466_ (.A1(net149),
    .A2(net238),
    .B1(net233),
    .B2(net152),
    .Y(_09926_));
 sky130_fd_sc_hd__and4_1 _18467_ (.A(net154),
    .B(net149),
    .C(net238),
    .D(net233),
    .X(_09927_));
 sky130_fd_sc_hd__o2bb2a_1 _18468_ (.A1_N(net243),
    .A2_N(net144),
    .B1(_09926_),
    .B2(_09927_),
    .X(_09928_));
 sky130_fd_sc_hd__and4bb_1 _18469_ (.A_N(_09926_),
    .B_N(_09927_),
    .C(net243),
    .D(net144),
    .X(_09929_));
 sky130_fd_sc_hd__or2_1 _18470_ (.A(_09928_),
    .B(_09929_),
    .X(_09930_));
 sky130_fd_sc_hd__o21ai_1 _18471_ (.A1(_09778_),
    .A2(_09781_),
    .B1(_09780_),
    .Y(_09931_));
 sky130_fd_sc_hd__nand2b_1 _18472_ (.A_N(_09930_),
    .B(_09931_),
    .Y(_09932_));
 sky130_fd_sc_hd__xor2_1 _18473_ (.A(_09930_),
    .B(_09931_),
    .X(_09933_));
 sky130_fd_sc_hd__or2_1 _18474_ (.A(_09925_),
    .B(_09933_),
    .X(_09934_));
 sky130_fd_sc_hd__xor2_1 _18475_ (.A(_09925_),
    .B(_09933_),
    .X(_09935_));
 sky130_fd_sc_hd__o21a_1 _18476_ (.A1(_09801_),
    .A2(_09803_),
    .B1(_09935_),
    .X(_09936_));
 sky130_fd_sc_hd__o21ai_1 _18477_ (.A1(_09801_),
    .A2(_09803_),
    .B1(_09935_),
    .Y(_09937_));
 sky130_fd_sc_hd__or3_1 _18478_ (.A(_09801_),
    .B(_09803_),
    .C(_09935_),
    .X(_09938_));
 sky130_fd_sc_hd__o211a_2 _18479_ (.A1(_09784_),
    .A2(_09786_),
    .B1(_09937_),
    .C1(_09938_),
    .X(_09939_));
 sky130_fd_sc_hd__a211oi_2 _18480_ (.A1(_09937_),
    .A2(_09938_),
    .B1(_09784_),
    .C1(_09786_),
    .Y(_09940_));
 sky130_fd_sc_hd__nor2_1 _18481_ (.A(_09796_),
    .B(_09799_),
    .Y(_09941_));
 sky130_fd_sc_hd__a31o_1 _18482_ (.A1(net174),
    .A2(net219),
    .A3(_09807_),
    .B1(_09806_),
    .X(_09942_));
 sky130_fd_sc_hd__a22o_1 _18483_ (.A1(net162),
    .A2(net225),
    .B1(net219),
    .B2(net169),
    .X(_09943_));
 sky130_fd_sc_hd__nand4_1 _18484_ (.A(net169),
    .B(net163),
    .C(net225),
    .D(net219),
    .Y(_09944_));
 sky130_fd_sc_hd__a22oi_1 _18485_ (.A1(net158),
    .A2(net229),
    .B1(_09943_),
    .B2(_09944_),
    .Y(_09945_));
 sky130_fd_sc_hd__and4_1 _18486_ (.A(net158),
    .B(net229),
    .C(_09943_),
    .D(_09944_),
    .X(_09946_));
 sky130_fd_sc_hd__or2_1 _18487_ (.A(_09945_),
    .B(_09946_),
    .X(_09947_));
 sky130_fd_sc_hd__and2b_1 _18488_ (.A_N(_09947_),
    .B(_09942_),
    .X(_09948_));
 sky130_fd_sc_hd__xnor2_2 _18489_ (.A(_09942_),
    .B(_09947_),
    .Y(_09949_));
 sky130_fd_sc_hd__and2b_1 _18490_ (.A_N(_09941_),
    .B(_09949_),
    .X(_09950_));
 sky130_fd_sc_hd__xnor2_2 _18491_ (.A(_09941_),
    .B(_09949_),
    .Y(_09951_));
 sky130_fd_sc_hd__nand2_1 _18492_ (.A(net174),
    .B(net215),
    .Y(_09952_));
 sky130_fd_sc_hd__and4_1 _18493_ (.A(net184),
    .B(net179),
    .C(net211),
    .D(net208),
    .X(_09953_));
 sky130_fd_sc_hd__a22o_1 _18494_ (.A1(net179),
    .A2(net211),
    .B1(net208),
    .B2(net184),
    .X(_09954_));
 sky130_fd_sc_hd__and2b_1 _18495_ (.A_N(_09953_),
    .B(_09954_),
    .X(_09955_));
 sky130_fd_sc_hd__xnor2_2 _18496_ (.A(_09952_),
    .B(_09955_),
    .Y(_09956_));
 sky130_fd_sc_hd__and2_1 _18497_ (.A(net187),
    .B(net205),
    .X(_09957_));
 sky130_fd_sc_hd__nand4_1 _18498_ (.A(net623),
    .B(net191),
    .C(net203),
    .D(net200),
    .Y(_09958_));
 sky130_fd_sc_hd__a22o_1 _18499_ (.A1(net190),
    .A2(net203),
    .B1(net200),
    .B2(net623),
    .X(_09959_));
 sky130_fd_sc_hd__nand3_1 _18500_ (.A(_09957_),
    .B(_09958_),
    .C(_09959_),
    .Y(_09960_));
 sky130_fd_sc_hd__a21o_1 _18501_ (.A1(_09958_),
    .A2(_09959_),
    .B1(_09957_),
    .X(_09961_));
 sky130_fd_sc_hd__a21bo_1 _18502_ (.A1(_09810_),
    .A2(_09812_),
    .B1_N(_09811_),
    .X(_09962_));
 sky130_fd_sc_hd__nand3_1 _18503_ (.A(_09960_),
    .B(_09961_),
    .C(_09962_),
    .Y(_09963_));
 sky130_fd_sc_hd__a21o_1 _18504_ (.A1(_09960_),
    .A2(_09961_),
    .B1(_09962_),
    .X(_09964_));
 sky130_fd_sc_hd__nand3_2 _18505_ (.A(_09956_),
    .B(_09963_),
    .C(_09964_),
    .Y(_09965_));
 sky130_fd_sc_hd__a21o_1 _18506_ (.A1(_09963_),
    .A2(_09964_),
    .B1(_09956_),
    .X(_09966_));
 sky130_fd_sc_hd__a21bo_1 _18507_ (.A1(_09809_),
    .A2(_09817_),
    .B1_N(_09816_),
    .X(_09967_));
 sky130_fd_sc_hd__nand3_4 _18508_ (.A(_09965_),
    .B(_09966_),
    .C(_09967_),
    .Y(_09968_));
 sky130_fd_sc_hd__a21o_1 _18509_ (.A1(_09965_),
    .A2(_09966_),
    .B1(_09967_),
    .X(_09969_));
 sky130_fd_sc_hd__and3_1 _18510_ (.A(_09951_),
    .B(_09968_),
    .C(_09969_),
    .X(_09970_));
 sky130_fd_sc_hd__nand3_2 _18511_ (.A(_09951_),
    .B(_09968_),
    .C(_09969_),
    .Y(_09971_));
 sky130_fd_sc_hd__a21oi_2 _18512_ (.A1(_09968_),
    .A2(_09969_),
    .B1(_09951_),
    .Y(_09972_));
 sky130_fd_sc_hd__a211oi_4 _18513_ (.A1(_09821_),
    .A2(_09824_),
    .B1(_09970_),
    .C1(_09972_),
    .Y(_09973_));
 sky130_fd_sc_hd__o211a_1 _18514_ (.A1(_09970_),
    .A2(_09972_),
    .B1(_09821_),
    .C1(_09824_),
    .X(_09974_));
 sky130_fd_sc_hd__nor4_1 _18515_ (.A(_09939_),
    .B(_09940_),
    .C(_09973_),
    .D(_09974_),
    .Y(_09975_));
 sky130_fd_sc_hd__or4_1 _18516_ (.A(_09939_),
    .B(_09940_),
    .C(_09973_),
    .D(_09974_),
    .X(_09976_));
 sky130_fd_sc_hd__o22ai_2 _18517_ (.A1(_09939_),
    .A2(_09940_),
    .B1(_09973_),
    .B2(_09974_),
    .Y(_09977_));
 sky130_fd_sc_hd__o211a_2 _18518_ (.A1(_09826_),
    .A2(_09828_),
    .B1(_09976_),
    .C1(_09977_),
    .X(_09978_));
 sky130_fd_sc_hd__a211oi_2 _18519_ (.A1(_09976_),
    .A2(_09977_),
    .B1(_09826_),
    .C1(_09828_),
    .Y(_09979_));
 sky130_fd_sc_hd__nor4_1 _18520_ (.A(_09918_),
    .B(_09920_),
    .C(_09978_),
    .D(_09979_),
    .Y(_09980_));
 sky130_fd_sc_hd__or4_1 _18521_ (.A(_09918_),
    .B(_09920_),
    .C(_09978_),
    .D(_09979_),
    .X(_09981_));
 sky130_fd_sc_hd__o22ai_1 _18522_ (.A1(_09918_),
    .A2(_09920_),
    .B1(_09978_),
    .B2(_09979_),
    .Y(_09982_));
 sky130_fd_sc_hd__o211a_1 _18523_ (.A1(_09831_),
    .A2(_09833_),
    .B1(_09981_),
    .C1(_09982_),
    .X(_09983_));
 sky130_fd_sc_hd__a211oi_1 _18524_ (.A1(_09981_),
    .A2(_09982_),
    .B1(_09831_),
    .C1(_09833_),
    .Y(_09984_));
 sky130_fd_sc_hd__nor4_2 _18525_ (.A(_09884_),
    .B(_09885_),
    .C(_09983_),
    .D(_09984_),
    .Y(_09985_));
 sky130_fd_sc_hd__o22a_1 _18526_ (.A1(_09884_),
    .A2(_09885_),
    .B1(_09983_),
    .B2(_09984_),
    .X(_09986_));
 sky130_fd_sc_hd__a211oi_2 _18527_ (.A1(_09836_),
    .A2(_09839_),
    .B1(_09985_),
    .C1(_09986_),
    .Y(_09987_));
 sky130_fd_sc_hd__o211a_1 _18528_ (.A1(_09985_),
    .A2(_09986_),
    .B1(_09836_),
    .C1(_09839_),
    .X(_09988_));
 sky130_fd_sc_hd__or3_2 _18529_ (.A(_09858_),
    .B(_09987_),
    .C(_09988_),
    .X(_09989_));
 sky130_fd_sc_hd__o21ai_2 _18530_ (.A1(_09987_),
    .A2(_09988_),
    .B1(_09858_),
    .Y(_09990_));
 sky130_fd_sc_hd__o211ai_4 _18531_ (.A1(_09841_),
    .A2(_09843_),
    .B1(_09989_),
    .C1(_09990_),
    .Y(_09991_));
 sky130_fd_sc_hd__a211o_1 _18532_ (.A1(_09989_),
    .A2(_09990_),
    .B1(_09841_),
    .C1(_09843_),
    .X(_09992_));
 sky130_fd_sc_hd__and3_1 _18533_ (.A(_09848_),
    .B(_09991_),
    .C(_09992_),
    .X(_09993_));
 sky130_fd_sc_hd__nand3_1 _18534_ (.A(_09848_),
    .B(_09991_),
    .C(_09992_),
    .Y(_09994_));
 sky130_fd_sc_hd__a21oi_1 _18535_ (.A1(_09991_),
    .A2(_09992_),
    .B1(_09848_),
    .Y(_09995_));
 sky130_fd_sc_hd__nor2_2 _18536_ (.A(_09993_),
    .B(_09995_),
    .Y(_09996_));
 sky130_fd_sc_hd__xnor2_4 _18537_ (.A(_09857_),
    .B(_09996_),
    .Y(_09997_));
 sky130_fd_sc_hd__nor2_1 _18538_ (.A(net43),
    .B(_05156_),
    .Y(_09998_));
 sky130_fd_sc_hd__a221o_1 _18539_ (.A1(net740),
    .A2(net8),
    .B1(_09997_),
    .B2(net10),
    .C1(_09998_),
    .X(_09999_));
 sky130_fd_sc_hd__mux2_1 _18540_ (.A0(net797),
    .A1(_09999_),
    .S(net1),
    .X(_00310_));
 sky130_fd_sc_hd__o21a_1 _18541_ (.A1(_09857_),
    .A2(_09995_),
    .B1(_09994_),
    .X(_10000_));
 sky130_fd_sc_hd__or2_4 _18542_ (.A(_09882_),
    .B(_09884_),
    .X(_10001_));
 sky130_fd_sc_hd__nor2_1 _18543_ (.A(_09878_),
    .B(_09880_),
    .Y(_10002_));
 sky130_fd_sc_hd__a22o_1 _18544_ (.A1(net316),
    .A2(net74),
    .B1(net71),
    .B2(net321),
    .X(_10003_));
 sky130_fd_sc_hd__and3_1 _18545_ (.A(net316),
    .B(net321),
    .C(net71),
    .X(_10004_));
 sky130_fd_sc_hd__a21bo_1 _18546_ (.A1(net74),
    .A2(_10004_),
    .B1_N(_10003_),
    .X(_10005_));
 sky130_fd_sc_hd__nand2_1 _18547_ (.A(net324),
    .B(net68),
    .Y(_10006_));
 sky130_fd_sc_hd__xnor2_1 _18548_ (.A(_10005_),
    .B(_10006_),
    .Y(_10007_));
 sky130_fd_sc_hd__nor2_1 _18549_ (.A(_09861_),
    .B(_10007_),
    .Y(_10008_));
 sky130_fd_sc_hd__and2_1 _18550_ (.A(_09861_),
    .B(_10007_),
    .X(_10009_));
 sky130_fd_sc_hd__or2_1 _18551_ (.A(_10008_),
    .B(_10009_),
    .X(_10010_));
 sky130_fd_sc_hd__or2_1 _18552_ (.A(_09864_),
    .B(_09866_),
    .X(_10011_));
 sky130_fd_sc_hd__a22oi_1 _18553_ (.A1(net301),
    .A2(net81),
    .B1(net78),
    .B2(net306),
    .Y(_10012_));
 sky130_fd_sc_hd__and4_1 _18554_ (.A(net301),
    .B(net306),
    .C(net81),
    .D(net78),
    .X(_10013_));
 sky130_fd_sc_hd__o2bb2a_1 _18555_ (.A1_N(net311),
    .A2_N(net75),
    .B1(_10012_),
    .B2(_10013_),
    .X(_10014_));
 sky130_fd_sc_hd__and4bb_1 _18556_ (.A_N(_10012_),
    .B_N(_10013_),
    .C(net311),
    .D(net75),
    .X(_10015_));
 sky130_fd_sc_hd__a211o_1 _18557_ (.A1(_09887_),
    .A2(_09889_),
    .B1(_10014_),
    .C1(_10015_),
    .X(_10016_));
 sky130_fd_sc_hd__o211ai_1 _18558_ (.A1(_10014_),
    .A2(_10015_),
    .B1(_09887_),
    .C1(_09889_),
    .Y(_10017_));
 sky130_fd_sc_hd__and2_1 _18559_ (.A(_10016_),
    .B(_10017_),
    .X(_10018_));
 sky130_fd_sc_hd__nand2_1 _18560_ (.A(_10011_),
    .B(_10018_),
    .Y(_10019_));
 sky130_fd_sc_hd__xnor2_1 _18561_ (.A(_10011_),
    .B(_10018_),
    .Y(_10020_));
 sky130_fd_sc_hd__a21oi_2 _18562_ (.A1(_09897_),
    .A2(_09899_),
    .B1(_10020_),
    .Y(_10021_));
 sky130_fd_sc_hd__inv_2 _18563_ (.A(_10021_),
    .Y(_10022_));
 sky130_fd_sc_hd__and3_1 _18564_ (.A(_09897_),
    .B(_09899_),
    .C(_10020_),
    .X(_10023_));
 sky130_fd_sc_hd__a211oi_1 _18565_ (.A1(_09867_),
    .A2(_09870_),
    .B1(_10021_),
    .C1(_10023_),
    .Y(_10024_));
 sky130_fd_sc_hd__a211o_1 _18566_ (.A1(_09867_),
    .A2(_09870_),
    .B1(_10021_),
    .C1(_10023_),
    .X(_10025_));
 sky130_fd_sc_hd__o211a_1 _18567_ (.A1(_10021_),
    .A2(_10023_),
    .B1(_09867_),
    .C1(_09870_),
    .X(_10026_));
 sky130_fd_sc_hd__a211oi_2 _18568_ (.A1(_09873_),
    .A2(_09876_),
    .B1(_10024_),
    .C1(_10026_),
    .Y(_10027_));
 sky130_fd_sc_hd__inv_2 _18569_ (.A(_10027_),
    .Y(_10028_));
 sky130_fd_sc_hd__o211a_1 _18570_ (.A1(_10024_),
    .A2(_10026_),
    .B1(_09873_),
    .C1(_09876_),
    .X(_10029_));
 sky130_fd_sc_hd__nor3_1 _18571_ (.A(_10010_),
    .B(_10027_),
    .C(_10029_),
    .Y(_10030_));
 sky130_fd_sc_hd__or3_1 _18572_ (.A(_10010_),
    .B(_10027_),
    .C(_10029_),
    .X(_10031_));
 sky130_fd_sc_hd__o21a_1 _18573_ (.A1(_10027_),
    .A2(_10029_),
    .B1(_10010_),
    .X(_10032_));
 sky130_fd_sc_hd__a211oi_2 _18574_ (.A1(_09916_),
    .A2(_09919_),
    .B1(_10030_),
    .C1(_10032_),
    .Y(_10033_));
 sky130_fd_sc_hd__o211a_1 _18575_ (.A1(_10030_),
    .A2(_10032_),
    .B1(_09916_),
    .C1(_09919_),
    .X(_10034_));
 sky130_fd_sc_hd__nor3_1 _18576_ (.A(_10002_),
    .B(_10033_),
    .C(_10034_),
    .Y(_10035_));
 sky130_fd_sc_hd__o21a_1 _18577_ (.A1(_10033_),
    .A2(_10034_),
    .B1(_10002_),
    .X(_10036_));
 sky130_fd_sc_hd__a22o_1 _18578_ (.A1(net286),
    .A2(net93),
    .B1(net89),
    .B2(net290),
    .X(_10037_));
 sky130_fd_sc_hd__nand4_2 _18579_ (.A(net286),
    .B(net290),
    .C(net93),
    .D(net90),
    .Y(_10038_));
 sky130_fd_sc_hd__a22o_1 _18580_ (.A1(net296),
    .A2(net85),
    .B1(_10037_),
    .B2(_10038_),
    .X(_10039_));
 sky130_fd_sc_hd__nand4_2 _18581_ (.A(net296),
    .B(net85),
    .C(_10037_),
    .D(_10038_),
    .Y(_10040_));
 sky130_fd_sc_hd__nand2_1 _18582_ (.A(_10039_),
    .B(_10040_),
    .Y(_10041_));
 sky130_fd_sc_hd__a22oi_1 _18583_ (.A1(net270),
    .A2(net109),
    .B1(net104),
    .B2(net276),
    .Y(_10042_));
 sky130_fd_sc_hd__and4_1 _18584_ (.A(net270),
    .B(net276),
    .C(net109),
    .D(net104),
    .X(_10043_));
 sky130_fd_sc_hd__o2bb2a_1 _18585_ (.A1_N(net281),
    .A2_N(net99),
    .B1(_10042_),
    .B2(_10043_),
    .X(_10044_));
 sky130_fd_sc_hd__and4bb_1 _18586_ (.A_N(_10042_),
    .B_N(_10043_),
    .C(net281),
    .D(net100),
    .X(_10045_));
 sky130_fd_sc_hd__nor2_1 _18587_ (.A(_10044_),
    .B(_10045_),
    .Y(_10046_));
 sky130_fd_sc_hd__or2_1 _18588_ (.A(_09892_),
    .B(_09894_),
    .X(_10047_));
 sky130_fd_sc_hd__nand2_1 _18589_ (.A(_10046_),
    .B(_10047_),
    .Y(_10048_));
 sky130_fd_sc_hd__xnor2_1 _18590_ (.A(_10046_),
    .B(_10047_),
    .Y(_10049_));
 sky130_fd_sc_hd__or2_2 _18591_ (.A(_10041_),
    .B(_10049_),
    .X(_10050_));
 sky130_fd_sc_hd__nand2_1 _18592_ (.A(_10041_),
    .B(_10049_),
    .Y(_10051_));
 sky130_fd_sc_hd__and2_1 _18593_ (.A(_10050_),
    .B(_10051_),
    .X(_10052_));
 sky130_fd_sc_hd__or2_1 _18594_ (.A(_09904_),
    .B(_09906_),
    .X(_10053_));
 sky130_fd_sc_hd__a22o_1 _18595_ (.A1(net253),
    .A2(net124),
    .B1(net119),
    .B2(net259),
    .X(_10054_));
 sky130_fd_sc_hd__nand4_1 _18596_ (.A(net253),
    .B(net259),
    .C(net124),
    .D(net119),
    .Y(_10055_));
 sky130_fd_sc_hd__a22oi_2 _18597_ (.A1(net266),
    .A2(net115),
    .B1(_10054_),
    .B2(_10055_),
    .Y(_10056_));
 sky130_fd_sc_hd__and4_1 _18598_ (.A(net266),
    .B(net115),
    .C(_10054_),
    .D(_10055_),
    .X(_10057_));
 sky130_fd_sc_hd__a211o_1 _18599_ (.A1(_09922_),
    .A2(_09924_),
    .B1(_10056_),
    .C1(_10057_),
    .X(_10058_));
 sky130_fd_sc_hd__o211ai_1 _18600_ (.A1(_10056_),
    .A2(_10057_),
    .B1(_09922_),
    .C1(_09924_),
    .Y(_10059_));
 sky130_fd_sc_hd__and2_1 _18601_ (.A(_10058_),
    .B(_10059_),
    .X(_10060_));
 sky130_fd_sc_hd__nand2_1 _18602_ (.A(_10053_),
    .B(_10060_),
    .Y(_10061_));
 sky130_fd_sc_hd__xnor2_2 _18603_ (.A(_10053_),
    .B(_10060_),
    .Y(_10062_));
 sky130_fd_sc_hd__a21oi_2 _18604_ (.A1(_09907_),
    .A2(_09910_),
    .B1(_10062_),
    .Y(_10063_));
 sky130_fd_sc_hd__a21o_1 _18605_ (.A1(_09907_),
    .A2(_09910_),
    .B1(_10062_),
    .X(_10064_));
 sky130_fd_sc_hd__nand3_1 _18606_ (.A(_09907_),
    .B(_09910_),
    .C(_10062_),
    .Y(_10065_));
 sky130_fd_sc_hd__and3_1 _18607_ (.A(_10052_),
    .B(_10064_),
    .C(_10065_),
    .X(_10066_));
 sky130_fd_sc_hd__nand3_2 _18608_ (.A(_10052_),
    .B(_10064_),
    .C(_10065_),
    .Y(_10067_));
 sky130_fd_sc_hd__a21o_1 _18609_ (.A1(_10064_),
    .A2(_10065_),
    .B1(_10052_),
    .X(_10068_));
 sky130_fd_sc_hd__o211ai_4 _18610_ (.A1(_09936_),
    .A2(_09939_),
    .B1(_10067_),
    .C1(_10068_),
    .Y(_10069_));
 sky130_fd_sc_hd__a211o_1 _18611_ (.A1(_10067_),
    .A2(_10068_),
    .B1(_09936_),
    .C1(_09939_),
    .X(_10070_));
 sky130_fd_sc_hd__o211a_1 _18612_ (.A1(_09912_),
    .A2(_09914_),
    .B1(_10069_),
    .C1(_10070_),
    .X(_10071_));
 sky130_fd_sc_hd__o211ai_2 _18613_ (.A1(_09912_),
    .A2(_09914_),
    .B1(_10069_),
    .C1(_10070_),
    .Y(_10072_));
 sky130_fd_sc_hd__a211oi_2 _18614_ (.A1(_10069_),
    .A2(_10070_),
    .B1(_09912_),
    .C1(_09914_),
    .Y(_10073_));
 sky130_fd_sc_hd__a22o_1 _18615_ (.A1(net243),
    .A2(net140),
    .B1(net135),
    .B2(net626),
    .X(_10074_));
 sky130_fd_sc_hd__and4_1 _18616_ (.A(net243),
    .B(net626),
    .C(net140),
    .D(net133),
    .X(_10075_));
 sky130_fd_sc_hd__inv_2 _18617_ (.A(_10075_),
    .Y(_10076_));
 sky130_fd_sc_hd__nand2_1 _18618_ (.A(_10074_),
    .B(_10076_),
    .Y(_10077_));
 sky130_fd_sc_hd__nand2_1 _18619_ (.A(net248),
    .B(net129),
    .Y(_10078_));
 sky130_fd_sc_hd__xnor2_1 _18620_ (.A(_10077_),
    .B(_10078_),
    .Y(_10079_));
 sky130_fd_sc_hd__a22o_1 _18621_ (.A1(net147),
    .A2(net233),
    .B1(net228),
    .B2(net154),
    .X(_10080_));
 sky130_fd_sc_hd__nand4_4 _18622_ (.A(net154),
    .B(net147),
    .C(net233),
    .D(net228),
    .Y(_10081_));
 sky130_fd_sc_hd__a22o_1 _18623_ (.A1(net144),
    .A2(net238),
    .B1(_10080_),
    .B2(_10081_),
    .X(_10082_));
 sky130_fd_sc_hd__nand4_2 _18624_ (.A(net144),
    .B(net238),
    .C(_10080_),
    .D(_10081_),
    .Y(_10083_));
 sky130_fd_sc_hd__nand2_1 _18625_ (.A(_10082_),
    .B(_10083_),
    .Y(_10084_));
 sky130_fd_sc_hd__or2_1 _18626_ (.A(_09927_),
    .B(_09929_),
    .X(_10085_));
 sky130_fd_sc_hd__nand2b_1 _18627_ (.A_N(_10084_),
    .B(_10085_),
    .Y(_10086_));
 sky130_fd_sc_hd__xor2_1 _18628_ (.A(_10084_),
    .B(_10085_),
    .X(_10087_));
 sky130_fd_sc_hd__or2_1 _18629_ (.A(_10079_),
    .B(_10087_),
    .X(_10088_));
 sky130_fd_sc_hd__xor2_1 _18630_ (.A(_10079_),
    .B(_10087_),
    .X(_10089_));
 sky130_fd_sc_hd__o21a_2 _18631_ (.A1(_09948_),
    .A2(_09950_),
    .B1(_10089_),
    .X(_10090_));
 sky130_fd_sc_hd__nor3_2 _18632_ (.A(_09948_),
    .B(_09950_),
    .C(_10089_),
    .Y(_10091_));
 sky130_fd_sc_hd__a211oi_4 _18633_ (.A1(_09932_),
    .A2(_09934_),
    .B1(_10090_),
    .C1(_10091_),
    .Y(_10092_));
 sky130_fd_sc_hd__o211a_1 _18634_ (.A1(_10090_),
    .A2(_10091_),
    .B1(_09932_),
    .C1(_09934_),
    .X(_10093_));
 sky130_fd_sc_hd__a41o_1 _18635_ (.A1(net169),
    .A2(net163),
    .A3(net225),
    .A4(net219),
    .B1(_09946_),
    .X(_10094_));
 sky130_fd_sc_hd__a31o_1 _18636_ (.A1(net174),
    .A2(net215),
    .A3(_09954_),
    .B1(_09953_),
    .X(_10095_));
 sky130_fd_sc_hd__a22o_1 _18637_ (.A1(net162),
    .A2(net219),
    .B1(net215),
    .B2(net169),
    .X(_10096_));
 sky130_fd_sc_hd__nand4_1 _18638_ (.A(net170),
    .B(net162),
    .C(net219),
    .D(net215),
    .Y(_10097_));
 sky130_fd_sc_hd__a22o_1 _18639_ (.A1(net157),
    .A2(net225),
    .B1(_10096_),
    .B2(_10097_),
    .X(_10098_));
 sky130_fd_sc_hd__nand4_1 _18640_ (.A(net157),
    .B(net225),
    .C(_10096_),
    .D(_10097_),
    .Y(_10099_));
 sky130_fd_sc_hd__and3_1 _18641_ (.A(_10095_),
    .B(_10098_),
    .C(_10099_),
    .X(_10100_));
 sky130_fd_sc_hd__a21o_1 _18642_ (.A1(_10098_),
    .A2(_10099_),
    .B1(_10095_),
    .X(_10101_));
 sky130_fd_sc_hd__and2b_1 _18643_ (.A_N(_10100_),
    .B(_10101_),
    .X(_10102_));
 sky130_fd_sc_hd__xor2_1 _18644_ (.A(_10094_),
    .B(_10102_),
    .X(_10103_));
 sky130_fd_sc_hd__nand2_1 _18645_ (.A(net173),
    .B(net211),
    .Y(_10104_));
 sky130_fd_sc_hd__a22o_1 _18646_ (.A1(net178),
    .A2(net208),
    .B1(net205),
    .B2(net183),
    .X(_10105_));
 sky130_fd_sc_hd__and3_1 _18647_ (.A(net183),
    .B(net178),
    .C(net208),
    .X(_10106_));
 sky130_fd_sc_hd__a21bo_1 _18648_ (.A1(net205),
    .A2(_10106_),
    .B1_N(_10105_),
    .X(_10107_));
 sky130_fd_sc_hd__xor2_1 _18649_ (.A(_10104_),
    .B(_10107_),
    .X(_10108_));
 sky130_fd_sc_hd__and2_1 _18650_ (.A(net187),
    .B(net203),
    .X(_10109_));
 sky130_fd_sc_hd__a22o_1 _18651_ (.A1(net190),
    .A2(net200),
    .B1(net198),
    .B2(net624),
    .X(_10110_));
 sky130_fd_sc_hd__nand4_1 _18652_ (.A(net624),
    .B(net190),
    .C(net200),
    .D(net198),
    .Y(_10111_));
 sky130_fd_sc_hd__nand3_1 _18653_ (.A(_10109_),
    .B(_10110_),
    .C(_10111_),
    .Y(_10112_));
 sky130_fd_sc_hd__a21o_1 _18654_ (.A1(_10110_),
    .A2(_10111_),
    .B1(_10109_),
    .X(_10113_));
 sky130_fd_sc_hd__a21bo_1 _18655_ (.A1(_09957_),
    .A2(_09959_),
    .B1_N(_09958_),
    .X(_10114_));
 sky130_fd_sc_hd__nand3_1 _18656_ (.A(_10112_),
    .B(_10113_),
    .C(_10114_),
    .Y(_10115_));
 sky130_fd_sc_hd__a21o_1 _18657_ (.A1(_10112_),
    .A2(_10113_),
    .B1(_10114_),
    .X(_10116_));
 sky130_fd_sc_hd__nand3_1 _18658_ (.A(_10108_),
    .B(_10115_),
    .C(_10116_),
    .Y(_10117_));
 sky130_fd_sc_hd__a21o_1 _18659_ (.A1(_10115_),
    .A2(_10116_),
    .B1(_10108_),
    .X(_10118_));
 sky130_fd_sc_hd__a21bo_1 _18660_ (.A1(_09956_),
    .A2(_09964_),
    .B1_N(_09963_),
    .X(_10119_));
 sky130_fd_sc_hd__nand3_2 _18661_ (.A(_10117_),
    .B(_10118_),
    .C(_10119_),
    .Y(_10120_));
 sky130_fd_sc_hd__a21o_1 _18662_ (.A1(_10117_),
    .A2(_10118_),
    .B1(_10119_),
    .X(_10121_));
 sky130_fd_sc_hd__and3_1 _18663_ (.A(_10103_),
    .B(_10120_),
    .C(_10121_),
    .X(_10122_));
 sky130_fd_sc_hd__nand3_1 _18664_ (.A(_10103_),
    .B(_10120_),
    .C(_10121_),
    .Y(_10123_));
 sky130_fd_sc_hd__a21oi_2 _18665_ (.A1(_10120_),
    .A2(_10121_),
    .B1(_10103_),
    .Y(_10124_));
 sky130_fd_sc_hd__a211oi_4 _18666_ (.A1(_09968_),
    .A2(_09971_),
    .B1(_10122_),
    .C1(_10124_),
    .Y(_10125_));
 sky130_fd_sc_hd__o211a_1 _18667_ (.A1(_10122_),
    .A2(_10124_),
    .B1(_09968_),
    .C1(_09971_),
    .X(_10126_));
 sky130_fd_sc_hd__nor4_2 _18668_ (.A(_10092_),
    .B(_10093_),
    .C(_10125_),
    .D(_10126_),
    .Y(_10127_));
 sky130_fd_sc_hd__or4_1 _18669_ (.A(_10092_),
    .B(_10093_),
    .C(_10125_),
    .D(_10126_),
    .X(_10128_));
 sky130_fd_sc_hd__o22ai_2 _18670_ (.A1(_10092_),
    .A2(_10093_),
    .B1(_10125_),
    .B2(_10126_),
    .Y(_10129_));
 sky130_fd_sc_hd__o211a_2 _18671_ (.A1(_09973_),
    .A2(_09975_),
    .B1(_10128_),
    .C1(_10129_),
    .X(_10130_));
 sky130_fd_sc_hd__a211oi_2 _18672_ (.A1(_10128_),
    .A2(_10129_),
    .B1(_09973_),
    .C1(_09975_),
    .Y(_10131_));
 sky130_fd_sc_hd__nor4_1 _18673_ (.A(_10071_),
    .B(_10073_),
    .C(_10130_),
    .D(_10131_),
    .Y(_10132_));
 sky130_fd_sc_hd__or4_1 _18674_ (.A(_10071_),
    .B(_10073_),
    .C(_10130_),
    .D(_10131_),
    .X(_10133_));
 sky130_fd_sc_hd__o22ai_2 _18675_ (.A1(_10071_),
    .A2(_10073_),
    .B1(_10130_),
    .B2(_10131_),
    .Y(_10134_));
 sky130_fd_sc_hd__o211ai_2 _18676_ (.A1(_09978_),
    .A2(_09980_),
    .B1(_10133_),
    .C1(_10134_),
    .Y(_10135_));
 sky130_fd_sc_hd__a211o_1 _18677_ (.A1(_10133_),
    .A2(_10134_),
    .B1(_09978_),
    .C1(_09980_),
    .X(_10136_));
 sky130_fd_sc_hd__or4bb_2 _18678_ (.A(_10035_),
    .B(_10036_),
    .C_N(_10135_),
    .D_N(_10136_),
    .X(_10137_));
 sky130_fd_sc_hd__a2bb2o_1 _18679_ (.A1_N(_10035_),
    .A2_N(_10036_),
    .B1(_10135_),
    .B2(_10136_),
    .X(_10138_));
 sky130_fd_sc_hd__o211a_1 _18680_ (.A1(_09983_),
    .A2(_09985_),
    .B1(_10137_),
    .C1(_10138_),
    .X(_10139_));
 sky130_fd_sc_hd__a211oi_1 _18681_ (.A1(_10137_),
    .A2(_10138_),
    .B1(_09983_),
    .C1(_09985_),
    .Y(_10140_));
 sky130_fd_sc_hd__nor2_2 _18682_ (.A(_10139_),
    .B(_10140_),
    .Y(_10141_));
 sky130_fd_sc_hd__xnor2_4 _18683_ (.A(_10001_),
    .B(_10141_),
    .Y(_10142_));
 sky130_fd_sc_hd__and2b_2 _18684_ (.A_N(_09987_),
    .B(_09989_),
    .X(_10143_));
 sky130_fd_sc_hd__or2_2 _18685_ (.A(_10142_),
    .B(_10143_),
    .X(_10144_));
 sky130_fd_sc_hd__xnor2_4 _18686_ (.A(_10142_),
    .B(_10143_),
    .Y(_10145_));
 sky130_fd_sc_hd__xor2_4 _18687_ (.A(_09991_),
    .B(_10145_),
    .X(_10146_));
 sky130_fd_sc_hd__xnor2_4 _18688_ (.A(_10000_),
    .B(_10146_),
    .Y(_10147_));
 sky130_fd_sc_hd__nor2_1 _18689_ (.A(net43),
    .B(_05305_),
    .Y(_10148_));
 sky130_fd_sc_hd__a221o_1 _18690_ (.A1(\temp[12] ),
    .A2(net8),
    .B1(_10147_),
    .B2(net10),
    .C1(_10148_),
    .X(_10149_));
 sky130_fd_sc_hd__mux2_1 _18691_ (.A0(net668),
    .A1(_10149_),
    .S(net1),
    .X(_00311_));
 sky130_fd_sc_hd__a21oi_4 _18692_ (.A1(_10001_),
    .A2(_10141_),
    .B1(_10139_),
    .Y(_10150_));
 sky130_fd_sc_hd__nor2_1 _18693_ (.A(_10033_),
    .B(_10035_),
    .Y(_10151_));
 sky130_fd_sc_hd__a22o_1 _18694_ (.A1(net311),
    .A2(net74),
    .B1(net71),
    .B2(net316),
    .X(_10152_));
 sky130_fd_sc_hd__inv_2 _18695_ (.A(_10152_),
    .Y(_10153_));
 sky130_fd_sc_hd__and4_1 _18696_ (.A(net311),
    .B(net316),
    .C(net74),
    .D(net71),
    .X(_10154_));
 sky130_fd_sc_hd__o2bb2a_1 _18697_ (.A1_N(net321),
    .A2_N(net68),
    .B1(_10153_),
    .B2(_10154_),
    .X(_10155_));
 sky130_fd_sc_hd__and4b_1 _18698_ (.A_N(_10154_),
    .B(net68),
    .C(net321),
    .D(_10152_),
    .X(_10156_));
 sky130_fd_sc_hd__or2_1 _18699_ (.A(_10155_),
    .B(_10156_),
    .X(_10157_));
 sky130_fd_sc_hd__a32o_1 _18700_ (.A1(net324),
    .A2(net68),
    .A3(_10003_),
    .B1(_10004_),
    .B2(net74),
    .X(_10158_));
 sky130_fd_sc_hd__or3b_1 _18701_ (.A(_10155_),
    .B(_10156_),
    .C_N(_10158_),
    .X(_10159_));
 sky130_fd_sc_hd__xor2_1 _18702_ (.A(_10157_),
    .B(_10158_),
    .X(_10160_));
 sky130_fd_sc_hd__nand2_1 _18703_ (.A(net324),
    .B(net65),
    .Y(_10161_));
 sky130_fd_sc_hd__or2_1 _18704_ (.A(_10160_),
    .B(_10161_),
    .X(_10162_));
 sky130_fd_sc_hd__xor2_1 _18705_ (.A(_10160_),
    .B(_10161_),
    .X(_10163_));
 sky130_fd_sc_hd__and2_1 _18706_ (.A(_10008_),
    .B(_10163_),
    .X(_10164_));
 sky130_fd_sc_hd__nor2_1 _18707_ (.A(_10008_),
    .B(_10163_),
    .Y(_10165_));
 sky130_fd_sc_hd__or2_1 _18708_ (.A(_10164_),
    .B(_10165_),
    .X(_10166_));
 sky130_fd_sc_hd__or2_1 _18709_ (.A(_10013_),
    .B(_10015_),
    .X(_10167_));
 sky130_fd_sc_hd__a22o_1 _18710_ (.A1(net296),
    .A2(net81),
    .B1(net78),
    .B2(net302),
    .X(_10168_));
 sky130_fd_sc_hd__nand4_1 _18711_ (.A(net296),
    .B(net302),
    .C(net81),
    .D(net78),
    .Y(_10169_));
 sky130_fd_sc_hd__a22oi_2 _18712_ (.A1(net307),
    .A2(net75),
    .B1(_10168_),
    .B2(_10169_),
    .Y(_10170_));
 sky130_fd_sc_hd__and4_1 _18713_ (.A(net307),
    .B(net75),
    .C(_10168_),
    .D(_10169_),
    .X(_10171_));
 sky130_fd_sc_hd__a211o_1 _18714_ (.A1(_10038_),
    .A2(_10040_),
    .B1(_10170_),
    .C1(_10171_),
    .X(_10172_));
 sky130_fd_sc_hd__o211ai_1 _18715_ (.A1(_10170_),
    .A2(_10171_),
    .B1(_10038_),
    .C1(_10040_),
    .Y(_10173_));
 sky130_fd_sc_hd__and2_1 _18716_ (.A(_10172_),
    .B(_10173_),
    .X(_10174_));
 sky130_fd_sc_hd__nand2_1 _18717_ (.A(_10167_),
    .B(_10174_),
    .Y(_10175_));
 sky130_fd_sc_hd__xnor2_2 _18718_ (.A(_10167_),
    .B(_10174_),
    .Y(_10176_));
 sky130_fd_sc_hd__a21oi_4 _18719_ (.A1(_10048_),
    .A2(_10050_),
    .B1(_10176_),
    .Y(_10177_));
 sky130_fd_sc_hd__and3_1 _18720_ (.A(_10048_),
    .B(_10050_),
    .C(_10176_),
    .X(_10178_));
 sky130_fd_sc_hd__a211oi_4 _18721_ (.A1(_10016_),
    .A2(_10019_),
    .B1(_10177_),
    .C1(_10178_),
    .Y(_10179_));
 sky130_fd_sc_hd__o211a_1 _18722_ (.A1(_10177_),
    .A2(_10178_),
    .B1(_10016_),
    .C1(_10019_),
    .X(_10180_));
 sky130_fd_sc_hd__a211oi_2 _18723_ (.A1(_10022_),
    .A2(_10025_),
    .B1(_10179_),
    .C1(_10180_),
    .Y(_10181_));
 sky130_fd_sc_hd__o211a_1 _18724_ (.A1(_10179_),
    .A2(_10180_),
    .B1(_10022_),
    .C1(_10025_),
    .X(_10182_));
 sky130_fd_sc_hd__nor3_1 _18725_ (.A(_10166_),
    .B(_10181_),
    .C(_10182_),
    .Y(_10183_));
 sky130_fd_sc_hd__o21a_1 _18726_ (.A1(_10181_),
    .A2(_10182_),
    .B1(_10166_),
    .X(_10184_));
 sky130_fd_sc_hd__a211oi_2 _18727_ (.A1(_10069_),
    .A2(_10072_),
    .B1(_10183_),
    .C1(_10184_),
    .Y(_10185_));
 sky130_fd_sc_hd__o211a_1 _18728_ (.A1(_10183_),
    .A2(_10184_),
    .B1(_10069_),
    .C1(_10072_),
    .X(_10186_));
 sky130_fd_sc_hd__a211oi_2 _18729_ (.A1(_10028_),
    .A2(_10031_),
    .B1(_10185_),
    .C1(_10186_),
    .Y(_10187_));
 sky130_fd_sc_hd__o211a_1 _18730_ (.A1(_10185_),
    .A2(_10186_),
    .B1(_10028_),
    .C1(_10031_),
    .X(_10188_));
 sky130_fd_sc_hd__a22oi_1 _18731_ (.A1(net281),
    .A2(net93),
    .B1(net90),
    .B2(net286),
    .Y(_10189_));
 sky130_fd_sc_hd__and4_1 _18732_ (.A(net281),
    .B(net286),
    .C(net93),
    .D(net90),
    .X(_10190_));
 sky130_fd_sc_hd__nor2_1 _18733_ (.A(_10189_),
    .B(_10190_),
    .Y(_10191_));
 sky130_fd_sc_hd__nand2_1 _18734_ (.A(net290),
    .B(net88),
    .Y(_10192_));
 sky130_fd_sc_hd__xnor2_1 _18735_ (.A(_10191_),
    .B(_10192_),
    .Y(_10193_));
 sky130_fd_sc_hd__a22o_1 _18736_ (.A1(net264),
    .A2(net109),
    .B1(net104),
    .B2(net270),
    .X(_10194_));
 sky130_fd_sc_hd__and4_1 _18737_ (.A(net264),
    .B(net270),
    .C(net109),
    .D(net104),
    .X(_10195_));
 sky130_fd_sc_hd__nand4_1 _18738_ (.A(net266),
    .B(net270),
    .C(net108),
    .D(net104),
    .Y(_10196_));
 sky130_fd_sc_hd__a22o_1 _18739_ (.A1(net276),
    .A2(net100),
    .B1(_10194_),
    .B2(_10196_),
    .X(_10197_));
 sky130_fd_sc_hd__and4_1 _18740_ (.A(net276),
    .B(net99),
    .C(_10194_),
    .D(_10196_),
    .X(_10198_));
 sky130_fd_sc_hd__nand4_1 _18741_ (.A(net276),
    .B(net99),
    .C(_10194_),
    .D(_10196_),
    .Y(_10199_));
 sky130_fd_sc_hd__o211a_1 _18742_ (.A1(_10043_),
    .A2(_10045_),
    .B1(_10197_),
    .C1(_10199_),
    .X(_10200_));
 sky130_fd_sc_hd__a211o_1 _18743_ (.A1(_10197_),
    .A2(_10199_),
    .B1(_10043_),
    .C1(_10045_),
    .X(_10201_));
 sky130_fd_sc_hd__nand2b_1 _18744_ (.A_N(_10200_),
    .B(_10201_),
    .Y(_10202_));
 sky130_fd_sc_hd__xnor2_1 _18745_ (.A(_10193_),
    .B(_10202_),
    .Y(_10203_));
 sky130_fd_sc_hd__a41o_1 _18746_ (.A1(net253),
    .A2(net259),
    .A3(net124),
    .A4(net119),
    .B1(_10057_),
    .X(_10204_));
 sky130_fd_sc_hd__a31o_1 _18747_ (.A1(net248),
    .A2(net129),
    .A3(_10074_),
    .B1(_10075_),
    .X(_10205_));
 sky130_fd_sc_hd__a22o_1 _18748_ (.A1(net248),
    .A2(net124),
    .B1(net119),
    .B2(net253),
    .X(_10206_));
 sky130_fd_sc_hd__nand4_2 _18749_ (.A(net248),
    .B(net253),
    .C(net124),
    .D(net120),
    .Y(_10207_));
 sky130_fd_sc_hd__a22o_1 _18750_ (.A1(net259),
    .A2(net116),
    .B1(_10206_),
    .B2(_10207_),
    .X(_10208_));
 sky130_fd_sc_hd__nand4_2 _18751_ (.A(net259),
    .B(net115),
    .C(_10206_),
    .D(_10207_),
    .Y(_10209_));
 sky130_fd_sc_hd__and3_1 _18752_ (.A(_10205_),
    .B(_10208_),
    .C(_10209_),
    .X(_10210_));
 sky130_fd_sc_hd__a21o_1 _18753_ (.A1(_10208_),
    .A2(_10209_),
    .B1(_10205_),
    .X(_10211_));
 sky130_fd_sc_hd__and2b_1 _18754_ (.A_N(_10210_),
    .B(_10211_),
    .X(_10212_));
 sky130_fd_sc_hd__xnor2_1 _18755_ (.A(_10204_),
    .B(_10212_),
    .Y(_10213_));
 sky130_fd_sc_hd__a21o_1 _18756_ (.A1(_10058_),
    .A2(_10061_),
    .B1(_10213_),
    .X(_10214_));
 sky130_fd_sc_hd__nand3_1 _18757_ (.A(_10058_),
    .B(_10061_),
    .C(_10213_),
    .Y(_10215_));
 sky130_fd_sc_hd__nand3_2 _18758_ (.A(_10203_),
    .B(_10214_),
    .C(_10215_),
    .Y(_10216_));
 sky130_fd_sc_hd__a21o_1 _18759_ (.A1(_10214_),
    .A2(_10215_),
    .B1(_10203_),
    .X(_10217_));
 sky130_fd_sc_hd__o211ai_4 _18760_ (.A1(_10090_),
    .A2(_10092_),
    .B1(_10216_),
    .C1(_10217_),
    .Y(_10218_));
 sky130_fd_sc_hd__a211o_1 _18761_ (.A1(_10216_),
    .A2(_10217_),
    .B1(_10090_),
    .C1(_10092_),
    .X(_10219_));
 sky130_fd_sc_hd__o211a_1 _18762_ (.A1(_10063_),
    .A2(_10066_),
    .B1(_10218_),
    .C1(_10219_),
    .X(_10220_));
 sky130_fd_sc_hd__o211ai_2 _18763_ (.A1(_10063_),
    .A2(_10066_),
    .B1(_10218_),
    .C1(_10219_),
    .Y(_10221_));
 sky130_fd_sc_hd__a211oi_2 _18764_ (.A1(_10218_),
    .A2(_10219_),
    .B1(_10063_),
    .C1(_10066_),
    .Y(_10222_));
 sky130_fd_sc_hd__a21o_1 _18765_ (.A1(_10094_),
    .A2(_10101_),
    .B1(_10100_),
    .X(_10223_));
 sky130_fd_sc_hd__a22o_1 _18766_ (.A1(net243),
    .A2(net135),
    .B1(net238),
    .B2(net138),
    .X(_10224_));
 sky130_fd_sc_hd__and3_1 _18767_ (.A(net243),
    .B(net138),
    .C(net135),
    .X(_10225_));
 sky130_fd_sc_hd__a21bo_1 _18768_ (.A1(net238),
    .A2(_10225_),
    .B1_N(_10224_),
    .X(_10226_));
 sky130_fd_sc_hd__nand2_1 _18769_ (.A(net626),
    .B(net129),
    .Y(_10227_));
 sky130_fd_sc_hd__xor2_1 _18770_ (.A(_10226_),
    .B(_10227_),
    .X(_10228_));
 sky130_fd_sc_hd__a22o_1 _18771_ (.A1(net149),
    .A2(net228),
    .B1(net224),
    .B2(net153),
    .X(_10229_));
 sky130_fd_sc_hd__nand4_1 _18772_ (.A(net153),
    .B(net148),
    .C(net228),
    .D(net224),
    .Y(_10230_));
 sky130_fd_sc_hd__and2_1 _18773_ (.A(net143),
    .B(net233),
    .X(_10231_));
 sky130_fd_sc_hd__a21oi_1 _18774_ (.A1(_10229_),
    .A2(_10230_),
    .B1(_10231_),
    .Y(_10232_));
 sky130_fd_sc_hd__and3_1 _18775_ (.A(_10229_),
    .B(_10230_),
    .C(_10231_),
    .X(_10233_));
 sky130_fd_sc_hd__a211o_1 _18776_ (.A1(_10081_),
    .A2(_10083_),
    .B1(_10232_),
    .C1(_10233_),
    .X(_10234_));
 sky130_fd_sc_hd__o211ai_1 _18777_ (.A1(_10232_),
    .A2(_10233_),
    .B1(_10081_),
    .C1(_10083_),
    .Y(_10235_));
 sky130_fd_sc_hd__nand3_1 _18778_ (.A(_10228_),
    .B(_10234_),
    .C(_10235_),
    .Y(_10236_));
 sky130_fd_sc_hd__a21o_1 _18779_ (.A1(_10234_),
    .A2(_10235_),
    .B1(_10228_),
    .X(_10237_));
 sky130_fd_sc_hd__and3_1 _18780_ (.A(_10223_),
    .B(_10236_),
    .C(_10237_),
    .X(_10238_));
 sky130_fd_sc_hd__a21oi_1 _18781_ (.A1(_10236_),
    .A2(_10237_),
    .B1(_10223_),
    .Y(_10239_));
 sky130_fd_sc_hd__a211oi_2 _18782_ (.A1(_10086_),
    .A2(_10088_),
    .B1(_10238_),
    .C1(_10239_),
    .Y(_10240_));
 sky130_fd_sc_hd__o211a_1 _18783_ (.A1(_10238_),
    .A2(_10239_),
    .B1(_10086_),
    .C1(_10088_),
    .X(_10241_));
 sky130_fd_sc_hd__nand2_1 _18784_ (.A(_10097_),
    .B(_10099_),
    .Y(_10242_));
 sky130_fd_sc_hd__a32o_1 _18785_ (.A1(net173),
    .A2(net211),
    .A3(_10105_),
    .B1(_10106_),
    .B2(net205),
    .X(_10243_));
 sky130_fd_sc_hd__a22o_1 _18786_ (.A1(net162),
    .A2(net218),
    .B1(net212),
    .B2(net169),
    .X(_10244_));
 sky130_fd_sc_hd__nand4_2 _18787_ (.A(net169),
    .B(net162),
    .C(net218),
    .D(net212),
    .Y(_10245_));
 sky130_fd_sc_hd__a22o_1 _18788_ (.A1(net157),
    .A2(net221),
    .B1(_10244_),
    .B2(_10245_),
    .X(_10246_));
 sky130_fd_sc_hd__nand4_1 _18789_ (.A(net157),
    .B(net221),
    .C(_10244_),
    .D(_10245_),
    .Y(_10247_));
 sky130_fd_sc_hd__and3_1 _18790_ (.A(_10243_),
    .B(_10246_),
    .C(_10247_),
    .X(_10248_));
 sky130_fd_sc_hd__a21o_1 _18791_ (.A1(_10246_),
    .A2(_10247_),
    .B1(_10243_),
    .X(_10249_));
 sky130_fd_sc_hd__and2b_1 _18792_ (.A_N(_10248_),
    .B(_10249_),
    .X(_10250_));
 sky130_fd_sc_hd__xor2_2 _18793_ (.A(_10242_),
    .B(_10250_),
    .X(_10251_));
 sky130_fd_sc_hd__a22oi_1 _18794_ (.A1(net178),
    .A2(net206),
    .B1(net202),
    .B2(net183),
    .Y(_10252_));
 sky130_fd_sc_hd__and4_1 _18795_ (.A(net183),
    .B(net178),
    .C(net206),
    .D(net202),
    .X(_10253_));
 sky130_fd_sc_hd__and4bb_1 _18796_ (.A_N(_10252_),
    .B_N(_10253_),
    .C(net174),
    .D(net209),
    .X(_10254_));
 sky130_fd_sc_hd__o2bb2a_1 _18797_ (.A1_N(net174),
    .A2_N(net209),
    .B1(_10252_),
    .B2(_10253_),
    .X(_10255_));
 sky130_fd_sc_hd__nor2_1 _18798_ (.A(_10254_),
    .B(_10255_),
    .Y(_10256_));
 sky130_fd_sc_hd__and2_1 _18799_ (.A(net187),
    .B(net200),
    .X(_10257_));
 sky130_fd_sc_hd__a22o_1 _18800_ (.A1(net190),
    .A2(net197),
    .B1(net195),
    .B2(net623),
    .X(_10258_));
 sky130_fd_sc_hd__nand4_2 _18801_ (.A(net623),
    .B(net190),
    .C(net198),
    .D(net195),
    .Y(_10259_));
 sky130_fd_sc_hd__nand3_1 _18802_ (.A(_10257_),
    .B(_10258_),
    .C(_10259_),
    .Y(_10260_));
 sky130_fd_sc_hd__a21o_1 _18803_ (.A1(_10258_),
    .A2(_10259_),
    .B1(_10257_),
    .X(_10261_));
 sky130_fd_sc_hd__a21bo_1 _18804_ (.A1(_10109_),
    .A2(_10110_),
    .B1_N(_10111_),
    .X(_10262_));
 sky130_fd_sc_hd__nand3_1 _18805_ (.A(_10260_),
    .B(_10261_),
    .C(_10262_),
    .Y(_10263_));
 sky130_fd_sc_hd__a21o_1 _18806_ (.A1(_10260_),
    .A2(_10261_),
    .B1(_10262_),
    .X(_10264_));
 sky130_fd_sc_hd__nand3_2 _18807_ (.A(_10256_),
    .B(_10263_),
    .C(_10264_),
    .Y(_10265_));
 sky130_fd_sc_hd__a21o_1 _18808_ (.A1(_10263_),
    .A2(_10264_),
    .B1(_10256_),
    .X(_10266_));
 sky130_fd_sc_hd__a21bo_1 _18809_ (.A1(_10108_),
    .A2(_10116_),
    .B1_N(_10115_),
    .X(_10267_));
 sky130_fd_sc_hd__nand3_4 _18810_ (.A(_10265_),
    .B(_10266_),
    .C(_10267_),
    .Y(_10268_));
 sky130_fd_sc_hd__a21o_1 _18811_ (.A1(_10265_),
    .A2(_10266_),
    .B1(_10267_),
    .X(_10269_));
 sky130_fd_sc_hd__and3_1 _18812_ (.A(_10251_),
    .B(_10268_),
    .C(_10269_),
    .X(_10270_));
 sky130_fd_sc_hd__nand3_2 _18813_ (.A(_10251_),
    .B(_10268_),
    .C(_10269_),
    .Y(_10271_));
 sky130_fd_sc_hd__a21oi_1 _18814_ (.A1(_10268_),
    .A2(_10269_),
    .B1(_10251_),
    .Y(_10272_));
 sky130_fd_sc_hd__a211o_2 _18815_ (.A1(_10120_),
    .A2(_10123_),
    .B1(_10270_),
    .C1(_10272_),
    .X(_10273_));
 sky130_fd_sc_hd__o211ai_2 _18816_ (.A1(_10270_),
    .A2(_10272_),
    .B1(_10120_),
    .C1(_10123_),
    .Y(_10274_));
 sky130_fd_sc_hd__or4bb_4 _18817_ (.A(_10240_),
    .B(_10241_),
    .C_N(_10273_),
    .D_N(_10274_),
    .X(_10275_));
 sky130_fd_sc_hd__a2bb2o_1 _18818_ (.A1_N(_10240_),
    .A2_N(_10241_),
    .B1(_10273_),
    .B2(_10274_),
    .X(_10276_));
 sky130_fd_sc_hd__o211a_2 _18819_ (.A1(_10125_),
    .A2(_10127_),
    .B1(_10275_),
    .C1(_10276_),
    .X(_10277_));
 sky130_fd_sc_hd__a211oi_4 _18820_ (.A1(_10275_),
    .A2(_10276_),
    .B1(_10125_),
    .C1(_10127_),
    .Y(_10278_));
 sky130_fd_sc_hd__nor4_2 _18821_ (.A(_10220_),
    .B(_10222_),
    .C(_10277_),
    .D(_10278_),
    .Y(_10279_));
 sky130_fd_sc_hd__or4_1 _18822_ (.A(_10220_),
    .B(_10222_),
    .C(_10277_),
    .D(_10278_),
    .X(_10280_));
 sky130_fd_sc_hd__o22ai_2 _18823_ (.A1(_10220_),
    .A2(_10222_),
    .B1(_10277_),
    .B2(_10278_),
    .Y(_10281_));
 sky130_fd_sc_hd__o211a_1 _18824_ (.A1(_10130_),
    .A2(_10132_),
    .B1(_10280_),
    .C1(_10281_),
    .X(_10282_));
 sky130_fd_sc_hd__a211oi_2 _18825_ (.A1(_10280_),
    .A2(_10281_),
    .B1(_10130_),
    .C1(_10132_),
    .Y(_10283_));
 sky130_fd_sc_hd__nor4_2 _18826_ (.A(_10187_),
    .B(_10188_),
    .C(_10282_),
    .D(_10283_),
    .Y(_10284_));
 sky130_fd_sc_hd__o22a_1 _18827_ (.A1(_10187_),
    .A2(_10188_),
    .B1(_10282_),
    .B2(_10283_),
    .X(_10285_));
 sky130_fd_sc_hd__a211oi_2 _18828_ (.A1(_10135_),
    .A2(_10137_),
    .B1(_10284_),
    .C1(_10285_),
    .Y(_10286_));
 sky130_fd_sc_hd__o211a_1 _18829_ (.A1(_10284_),
    .A2(_10285_),
    .B1(_10135_),
    .C1(_10137_),
    .X(_10287_));
 sky130_fd_sc_hd__nor3_2 _18830_ (.A(_10151_),
    .B(_10286_),
    .C(_10287_),
    .Y(_10288_));
 sky130_fd_sc_hd__o21a_1 _18831_ (.A1(_10286_),
    .A2(_10287_),
    .B1(_10151_),
    .X(_10289_));
 sky130_fd_sc_hd__nor2_2 _18832_ (.A(_10288_),
    .B(_10289_),
    .Y(_10290_));
 sky130_fd_sc_hd__or3_1 _18833_ (.A(_10150_),
    .B(_10288_),
    .C(_10289_),
    .X(_10291_));
 sky130_fd_sc_hd__xnor2_4 _18834_ (.A(_10150_),
    .B(_10290_),
    .Y(_10292_));
 sky130_fd_sc_hd__nand2b_1 _18835_ (.A_N(_10144_),
    .B(_10292_),
    .Y(_10293_));
 sky130_fd_sc_hd__xnor2_1 _18836_ (.A(_10144_),
    .B(_10292_),
    .Y(_10294_));
 sky130_fd_sc_hd__xor2_4 _18837_ (.A(_10144_),
    .B(_10292_),
    .X(_10295_));
 sky130_fd_sc_hd__a21oi_1 _18838_ (.A1(_09991_),
    .A2(_09994_),
    .B1(_10145_),
    .Y(_10296_));
 sky130_fd_sc_hd__nand2_1 _18839_ (.A(_09996_),
    .B(_10146_),
    .Y(_10297_));
 sky130_fd_sc_hd__o21ba_2 _18840_ (.A1(_09857_),
    .A2(_10297_),
    .B1_N(_10296_),
    .X(_10298_));
 sky130_fd_sc_hd__xnor2_4 _18841_ (.A(_10295_),
    .B(_10298_),
    .Y(_10299_));
 sky130_fd_sc_hd__nor2_1 _18842_ (.A(_03049_),
    .B(_10299_),
    .Y(_10300_));
 sky130_fd_sc_hd__a221o_1 _18843_ (.A1(net693),
    .A2(net8),
    .B1(_05457_),
    .B2(_03052_),
    .C1(_10300_),
    .X(_10301_));
 sky130_fd_sc_hd__mux2_1 _18844_ (.A0(net761),
    .A1(_10301_),
    .S(net1),
    .X(_00312_));
 sky130_fd_sc_hd__o21a_1 _18845_ (.A1(_10295_),
    .A2(_10298_),
    .B1(_10293_),
    .X(_10302_));
 sky130_fd_sc_hd__nor2_1 _18846_ (.A(_10185_),
    .B(_10187_),
    .Y(_10303_));
 sky130_fd_sc_hd__or2_1 _18847_ (.A(_10181_),
    .B(_10183_),
    .X(_10304_));
 sky130_fd_sc_hd__a22oi_1 _18848_ (.A1(net301),
    .A2(net75),
    .B1(net74),
    .B2(net306),
    .Y(_10305_));
 sky130_fd_sc_hd__and4_1 _18849_ (.A(net301),
    .B(net306),
    .C(\mul1.b[26] ),
    .D(net74),
    .X(_10306_));
 sky130_fd_sc_hd__o2bb2a_1 _18850_ (.A1_N(net312),
    .A2_N(net71),
    .B1(_10305_),
    .B2(_10306_),
    .X(_10307_));
 sky130_fd_sc_hd__and4bb_1 _18851_ (.A_N(_10305_),
    .B_N(_10306_),
    .C(net312),
    .D(net71),
    .X(_10308_));
 sky130_fd_sc_hd__nor2_1 _18852_ (.A(_10307_),
    .B(_10308_),
    .Y(_10309_));
 sky130_fd_sc_hd__nor2_1 _18853_ (.A(_10154_),
    .B(_10156_),
    .Y(_10310_));
 sky130_fd_sc_hd__or3_1 _18854_ (.A(_10307_),
    .B(_10308_),
    .C(_10310_),
    .X(_10311_));
 sky130_fd_sc_hd__xnor2_1 _18855_ (.A(_10309_),
    .B(_10310_),
    .Y(_10312_));
 sky130_fd_sc_hd__a22oi_2 _18856_ (.A1(net316),
    .A2(net68),
    .B1(net65),
    .B2(net321),
    .Y(_10313_));
 sky130_fd_sc_hd__and4_1 _18857_ (.A(net316),
    .B(net321),
    .C(net68),
    .D(net65),
    .X(_10314_));
 sky130_fd_sc_hd__o22a_1 _18858_ (.A1(net325),
    .A2(net56),
    .B1(_10313_),
    .B2(_10314_),
    .X(_10315_));
 sky130_fd_sc_hd__nor4_1 _18859_ (.A(net325),
    .B(net56),
    .C(_10313_),
    .D(_10314_),
    .Y(_10316_));
 sky130_fd_sc_hd__or2_1 _18860_ (.A(_10315_),
    .B(_10316_),
    .X(_10317_));
 sky130_fd_sc_hd__inv_2 _18861_ (.A(_10317_),
    .Y(_10318_));
 sky130_fd_sc_hd__nand2_1 _18862_ (.A(_10312_),
    .B(_10318_),
    .Y(_10319_));
 sky130_fd_sc_hd__or2_1 _18863_ (.A(_10312_),
    .B(_10318_),
    .X(_10320_));
 sky130_fd_sc_hd__nand2_1 _18864_ (.A(_10319_),
    .B(_10320_),
    .Y(_10321_));
 sky130_fd_sc_hd__a21oi_2 _18865_ (.A1(_10159_),
    .A2(_10162_),
    .B1(_10321_),
    .Y(_10322_));
 sky130_fd_sc_hd__and3_1 _18866_ (.A(_10159_),
    .B(_10162_),
    .C(_10321_),
    .X(_10323_));
 sky130_fd_sc_hd__a21oi_1 _18867_ (.A1(_10193_),
    .A2(_10201_),
    .B1(_10200_),
    .Y(_10324_));
 sky130_fd_sc_hd__a41o_1 _18868_ (.A1(net297),
    .A2(net301),
    .A3(net82),
    .A4(\mul1.b[25] ),
    .B1(_10171_),
    .X(_10325_));
 sky130_fd_sc_hd__o21bai_1 _18869_ (.A1(_10189_),
    .A2(_10192_),
    .B1_N(_10190_),
    .Y(_10326_));
 sky130_fd_sc_hd__a22o_1 _18870_ (.A1(net285),
    .A2(net85),
    .B1(net81),
    .B2(net290),
    .X(_10327_));
 sky130_fd_sc_hd__nand4_2 _18871_ (.A(net285),
    .B(net290),
    .C(net88),
    .D(net81),
    .Y(_10328_));
 sky130_fd_sc_hd__a22o_1 _18872_ (.A1(net296),
    .A2(net78),
    .B1(_10327_),
    .B2(_10328_),
    .X(_10329_));
 sky130_fd_sc_hd__nand4_2 _18873_ (.A(net296),
    .B(\mul1.b[25] ),
    .C(_10327_),
    .D(_10328_),
    .Y(_10330_));
 sky130_fd_sc_hd__nand3_2 _18874_ (.A(_10326_),
    .B(_10329_),
    .C(_10330_),
    .Y(_10331_));
 sky130_fd_sc_hd__a21o_1 _18875_ (.A1(_10329_),
    .A2(_10330_),
    .B1(_10326_),
    .X(_10332_));
 sky130_fd_sc_hd__nand3_2 _18876_ (.A(_10325_),
    .B(_10331_),
    .C(_10332_),
    .Y(_10333_));
 sky130_fd_sc_hd__a21o_1 _18877_ (.A1(_10331_),
    .A2(_10332_),
    .B1(_10325_),
    .X(_10334_));
 sky130_fd_sc_hd__and3b_2 _18878_ (.A_N(_10324_),
    .B(_10333_),
    .C(_10334_),
    .X(_10335_));
 sky130_fd_sc_hd__a21boi_2 _18879_ (.A1(_10333_),
    .A2(_10334_),
    .B1_N(_10324_),
    .Y(_10336_));
 sky130_fd_sc_hd__a211oi_2 _18880_ (.A1(_10172_),
    .A2(_10175_),
    .B1(_10335_),
    .C1(_10336_),
    .Y(_10337_));
 sky130_fd_sc_hd__inv_2 _18881_ (.A(_10337_),
    .Y(_10338_));
 sky130_fd_sc_hd__o211ai_2 _18882_ (.A1(_10335_),
    .A2(_10336_),
    .B1(_10172_),
    .C1(_10175_),
    .Y(_10339_));
 sky130_fd_sc_hd__o211a_1 _18883_ (.A1(_10177_),
    .A2(_10179_),
    .B1(_10338_),
    .C1(_10339_),
    .X(_10340_));
 sky130_fd_sc_hd__a211oi_2 _18884_ (.A1(_10338_),
    .A2(_10339_),
    .B1(_10177_),
    .C1(_10179_),
    .Y(_10341_));
 sky130_fd_sc_hd__nor4_2 _18885_ (.A(_10322_),
    .B(_10323_),
    .C(_10340_),
    .D(_10341_),
    .Y(_10342_));
 sky130_fd_sc_hd__o22a_1 _18886_ (.A1(_10322_),
    .A2(_10323_),
    .B1(_10340_),
    .B2(_10341_),
    .X(_10343_));
 sky130_fd_sc_hd__a211o_1 _18887_ (.A1(_10218_),
    .A2(_10221_),
    .B1(_10342_),
    .C1(_10343_),
    .X(_10344_));
 sky130_fd_sc_hd__o211ai_2 _18888_ (.A1(_10342_),
    .A2(_10343_),
    .B1(_10218_),
    .C1(_10221_),
    .Y(_10345_));
 sky130_fd_sc_hd__and3_1 _18889_ (.A(_10304_),
    .B(_10344_),
    .C(_10345_),
    .X(_10346_));
 sky130_fd_sc_hd__a21oi_1 _18890_ (.A1(_10344_),
    .A2(_10345_),
    .B1(_10304_),
    .Y(_10347_));
 sky130_fd_sc_hd__a22o_1 _18891_ (.A1(net270),
    .A2(net99),
    .B1(net94),
    .B2(net276),
    .X(_10348_));
 sky130_fd_sc_hd__nand4_4 _18892_ (.A(net270),
    .B(net275),
    .C(net100),
    .D(net94),
    .Y(_10349_));
 sky130_fd_sc_hd__a22o_1 _18893_ (.A1(net280),
    .A2(net90),
    .B1(_10348_),
    .B2(_10349_),
    .X(_10350_));
 sky130_fd_sc_hd__nand4_2 _18894_ (.A(net280),
    .B(net90),
    .C(_10348_),
    .D(_10349_),
    .Y(_10351_));
 sky130_fd_sc_hd__and2_1 _18895_ (.A(_10350_),
    .B(_10351_),
    .X(_10352_));
 sky130_fd_sc_hd__a22o_1 _18896_ (.A1(net253),
    .A2(net115),
    .B1(net109),
    .B2(net260),
    .X(_10353_));
 sky130_fd_sc_hd__and4_1 _18897_ (.A(net253),
    .B(net259),
    .C(net115),
    .D(net109),
    .X(_10354_));
 sky130_fd_sc_hd__nand4_1 _18898_ (.A(net254),
    .B(net260),
    .C(net115),
    .D(net109),
    .Y(_10355_));
 sky130_fd_sc_hd__a22o_1 _18899_ (.A1(net264),
    .A2(net104),
    .B1(_10353_),
    .B2(_10355_),
    .X(_10356_));
 sky130_fd_sc_hd__and4_1 _18900_ (.A(net264),
    .B(net104),
    .C(_10353_),
    .D(_10355_),
    .X(_10357_));
 sky130_fd_sc_hd__nand4_1 _18901_ (.A(net264),
    .B(net103),
    .C(_10353_),
    .D(_10355_),
    .Y(_10358_));
 sky130_fd_sc_hd__o211a_1 _18902_ (.A1(_10195_),
    .A2(_10198_),
    .B1(_10356_),
    .C1(_10358_),
    .X(_10359_));
 sky130_fd_sc_hd__a211o_1 _18903_ (.A1(_10356_),
    .A2(_10358_),
    .B1(_10195_),
    .C1(_10198_),
    .X(_10360_));
 sky130_fd_sc_hd__and2b_1 _18904_ (.A_N(_10359_),
    .B(_10360_),
    .X(_10361_));
 sky130_fd_sc_hd__xnor2_1 _18905_ (.A(_10352_),
    .B(_10361_),
    .Y(_10362_));
 sky130_fd_sc_hd__nand2_1 _18906_ (.A(_10207_),
    .B(_10209_),
    .Y(_10363_));
 sky130_fd_sc_hd__a32o_1 _18907_ (.A1(net626),
    .A2(net130),
    .A3(_10224_),
    .B1(_10225_),
    .B2(net238),
    .X(_10364_));
 sky130_fd_sc_hd__a22o_1 _18908_ (.A1(net243),
    .A2(net130),
    .B1(net124),
    .B2(net626),
    .X(_10365_));
 sky130_fd_sc_hd__nand4_2 _18909_ (.A(net243),
    .B(net626),
    .C(net130),
    .D(net125),
    .Y(_10366_));
 sky130_fd_sc_hd__a22o_1 _18910_ (.A1(net249),
    .A2(net119),
    .B1(_10365_),
    .B2(_10366_),
    .X(_10367_));
 sky130_fd_sc_hd__nand4_1 _18911_ (.A(net248),
    .B(net119),
    .C(_10365_),
    .D(_10366_),
    .Y(_10368_));
 sky130_fd_sc_hd__nand3_1 _18912_ (.A(_10364_),
    .B(_10367_),
    .C(_10368_),
    .Y(_10369_));
 sky130_fd_sc_hd__a21o_1 _18913_ (.A1(_10367_),
    .A2(_10368_),
    .B1(_10364_),
    .X(_10370_));
 sky130_fd_sc_hd__nand3_1 _18914_ (.A(_10363_),
    .B(_10369_),
    .C(_10370_),
    .Y(_10371_));
 sky130_fd_sc_hd__a21o_1 _18915_ (.A1(_10369_),
    .A2(_10370_),
    .B1(_10363_),
    .X(_10372_));
 sky130_fd_sc_hd__a21o_1 _18916_ (.A1(_10204_),
    .A2(_10211_),
    .B1(_10210_),
    .X(_10373_));
 sky130_fd_sc_hd__and3_1 _18917_ (.A(_10371_),
    .B(_10372_),
    .C(_10373_),
    .X(_10374_));
 sky130_fd_sc_hd__a21oi_1 _18918_ (.A1(_10371_),
    .A2(_10372_),
    .B1(_10373_),
    .Y(_10375_));
 sky130_fd_sc_hd__or3_1 _18919_ (.A(_10362_),
    .B(_10374_),
    .C(_10375_),
    .X(_10376_));
 sky130_fd_sc_hd__o21ai_1 _18920_ (.A1(_10374_),
    .A2(_10375_),
    .B1(_10362_),
    .Y(_10377_));
 sky130_fd_sc_hd__o211a_1 _18921_ (.A1(_10238_),
    .A2(_10240_),
    .B1(_10376_),
    .C1(_10377_),
    .X(_10378_));
 sky130_fd_sc_hd__a211oi_1 _18922_ (.A1(_10376_),
    .A2(_10377_),
    .B1(_10238_),
    .C1(_10240_),
    .Y(_10379_));
 sky130_fd_sc_hd__a211oi_2 _18923_ (.A1(_10214_),
    .A2(_10216_),
    .B1(_10378_),
    .C1(_10379_),
    .Y(_10380_));
 sky130_fd_sc_hd__o211a_1 _18924_ (.A1(_10378_),
    .A2(_10379_),
    .B1(_10214_),
    .C1(_10216_),
    .X(_10381_));
 sky130_fd_sc_hd__nand2_1 _18925_ (.A(_10234_),
    .B(_10236_),
    .Y(_10382_));
 sky130_fd_sc_hd__a21o_1 _18926_ (.A1(_10242_),
    .A2(_10249_),
    .B1(_10248_),
    .X(_10383_));
 sky130_fd_sc_hd__nand2_1 _18927_ (.A(net134),
    .B(net238),
    .Y(_10384_));
 sky130_fd_sc_hd__a22o_1 _18928_ (.A1(net138),
    .A2(net233),
    .B1(net228),
    .B2(\mul1.b[11] ),
    .X(_10385_));
 sky130_fd_sc_hd__and3_1 _18929_ (.A(\mul1.b[11] ),
    .B(net140),
    .C(net228),
    .X(_10386_));
 sky130_fd_sc_hd__a21bo_1 _18930_ (.A1(net233),
    .A2(_10386_),
    .B1_N(_10385_),
    .X(_10387_));
 sky130_fd_sc_hd__xor2_1 _18931_ (.A(_10384_),
    .B(_10387_),
    .X(_10388_));
 sky130_fd_sc_hd__and2_1 _18932_ (.A(net149),
    .B(net224),
    .X(_10389_));
 sky130_fd_sc_hd__a22o_1 _18933_ (.A1(net154),
    .A2(net219),
    .B1(net215),
    .B2(net158),
    .X(_10390_));
 sky130_fd_sc_hd__nand4_2 _18934_ (.A(net158),
    .B(net154),
    .C(net219),
    .D(net215),
    .Y(_10391_));
 sky130_fd_sc_hd__a21o_1 _18935_ (.A1(_10390_),
    .A2(_10391_),
    .B1(_10389_),
    .X(_10392_));
 sky130_fd_sc_hd__nand3_1 _18936_ (.A(_10389_),
    .B(_10390_),
    .C(_10391_),
    .Y(_10393_));
 sky130_fd_sc_hd__a21bo_1 _18937_ (.A1(_10229_),
    .A2(_10231_),
    .B1_N(_10230_),
    .X(_10394_));
 sky130_fd_sc_hd__nand3_1 _18938_ (.A(_10392_),
    .B(_10393_),
    .C(_10394_),
    .Y(_10395_));
 sky130_fd_sc_hd__a21o_1 _18939_ (.A1(_10392_),
    .A2(_10393_),
    .B1(_10394_),
    .X(_10396_));
 sky130_fd_sc_hd__nand3_1 _18940_ (.A(_10388_),
    .B(_10395_),
    .C(_10396_),
    .Y(_10397_));
 sky130_fd_sc_hd__a21o_1 _18941_ (.A1(_10395_),
    .A2(_10396_),
    .B1(_10388_),
    .X(_10398_));
 sky130_fd_sc_hd__nand3_2 _18942_ (.A(_10383_),
    .B(_10397_),
    .C(_10398_),
    .Y(_10399_));
 sky130_fd_sc_hd__a21o_1 _18943_ (.A1(_10397_),
    .A2(_10398_),
    .B1(_10383_),
    .X(_10400_));
 sky130_fd_sc_hd__nand3_2 _18944_ (.A(_10382_),
    .B(_10399_),
    .C(_10400_),
    .Y(_10401_));
 sky130_fd_sc_hd__a21o_1 _18945_ (.A1(_10399_),
    .A2(_10400_),
    .B1(_10382_),
    .X(_10402_));
 sky130_fd_sc_hd__nand2_1 _18946_ (.A(_10401_),
    .B(_10402_),
    .Y(_10403_));
 sky130_fd_sc_hd__nand2_1 _18947_ (.A(_10245_),
    .B(_10247_),
    .Y(_10404_));
 sky130_fd_sc_hd__a22o_1 _18948_ (.A1(net167),
    .A2(net209),
    .B1(net206),
    .B2(net173),
    .X(_10405_));
 sky130_fd_sc_hd__nand4_2 _18949_ (.A(net173),
    .B(net167),
    .C(net209),
    .D(net206),
    .Y(_10406_));
 sky130_fd_sc_hd__a22o_1 _18950_ (.A1(net161),
    .A2(net212),
    .B1(_10405_),
    .B2(_10406_),
    .X(_10407_));
 sky130_fd_sc_hd__nand4_2 _18951_ (.A(net163),
    .B(net212),
    .C(_10405_),
    .D(_10406_),
    .Y(_10408_));
 sky130_fd_sc_hd__o211a_1 _18952_ (.A1(_10253_),
    .A2(_10254_),
    .B1(_10407_),
    .C1(_10408_),
    .X(_10409_));
 sky130_fd_sc_hd__a211o_1 _18953_ (.A1(_10407_),
    .A2(_10408_),
    .B1(_10253_),
    .C1(_10254_),
    .X(_10410_));
 sky130_fd_sc_hd__nand2b_1 _18954_ (.A_N(_10409_),
    .B(_10410_),
    .Y(_10411_));
 sky130_fd_sc_hd__xnor2_2 _18955_ (.A(_10404_),
    .B(_10411_),
    .Y(_10412_));
 sky130_fd_sc_hd__nand2_1 _18956_ (.A(net178),
    .B(net202),
    .Y(_10413_));
 sky130_fd_sc_hd__a22o_1 _18957_ (.A1(net183),
    .A2(net199),
    .B1(net197),
    .B2(net187),
    .X(_10414_));
 sky130_fd_sc_hd__and3_1 _18958_ (.A(net187),
    .B(net183),
    .C(net197),
    .X(_10415_));
 sky130_fd_sc_hd__a21bo_1 _18959_ (.A1(net199),
    .A2(_10415_),
    .B1_N(_10414_),
    .X(_10416_));
 sky130_fd_sc_hd__xor2_2 _18960_ (.A(_10413_),
    .B(_10416_),
    .X(_10417_));
 sky130_fd_sc_hd__nand2_1 _18961_ (.A(net190),
    .B(net196),
    .Y(_10418_));
 sky130_fd_sc_hd__a21oi_1 _18962_ (.A1(net623),
    .A2(net193),
    .B1(net62),
    .Y(_10419_));
 sky130_fd_sc_hd__and3_1 _18963_ (.A(net623),
    .B(net193),
    .C(net62),
    .X(_10420_));
 sky130_fd_sc_hd__or3_1 _18964_ (.A(_10418_),
    .B(_10419_),
    .C(_10420_),
    .X(_10421_));
 sky130_fd_sc_hd__o21ai_1 _18965_ (.A1(_10419_),
    .A2(_10420_),
    .B1(_10418_),
    .Y(_10422_));
 sky130_fd_sc_hd__a21bo_1 _18966_ (.A1(_10257_),
    .A2(_10258_),
    .B1_N(_10259_),
    .X(_10423_));
 sky130_fd_sc_hd__nand3_1 _18967_ (.A(_10421_),
    .B(_10422_),
    .C(_10423_),
    .Y(_10424_));
 sky130_fd_sc_hd__a21o_1 _18968_ (.A1(_10421_),
    .A2(_10422_),
    .B1(_10423_),
    .X(_10425_));
 sky130_fd_sc_hd__nand3_2 _18969_ (.A(_10417_),
    .B(_10424_),
    .C(_10425_),
    .Y(_10426_));
 sky130_fd_sc_hd__a21o_1 _18970_ (.A1(_10424_),
    .A2(_10425_),
    .B1(_10417_),
    .X(_10427_));
 sky130_fd_sc_hd__a21bo_1 _18971_ (.A1(_10256_),
    .A2(_10264_),
    .B1_N(_10263_),
    .X(_10428_));
 sky130_fd_sc_hd__nand3_4 _18972_ (.A(_10426_),
    .B(_10427_),
    .C(_10428_),
    .Y(_10429_));
 sky130_fd_sc_hd__a21o_1 _18973_ (.A1(_10426_),
    .A2(_10427_),
    .B1(_10428_),
    .X(_10430_));
 sky130_fd_sc_hd__and3_1 _18974_ (.A(_10412_),
    .B(_10429_),
    .C(_10430_),
    .X(_10431_));
 sky130_fd_sc_hd__nand3_2 _18975_ (.A(_10412_),
    .B(_10429_),
    .C(_10430_),
    .Y(_10432_));
 sky130_fd_sc_hd__a21oi_2 _18976_ (.A1(_10429_),
    .A2(_10430_),
    .B1(_10412_),
    .Y(_10433_));
 sky130_fd_sc_hd__a211oi_4 _18977_ (.A1(_10268_),
    .A2(_10271_),
    .B1(_10431_),
    .C1(_10433_),
    .Y(_10434_));
 sky130_fd_sc_hd__o211a_1 _18978_ (.A1(_10431_),
    .A2(_10433_),
    .B1(_10268_),
    .C1(_10271_),
    .X(_10435_));
 sky130_fd_sc_hd__nor3_2 _18979_ (.A(_10403_),
    .B(_10434_),
    .C(_10435_),
    .Y(_10436_));
 sky130_fd_sc_hd__o21a_1 _18980_ (.A1(_10434_),
    .A2(_10435_),
    .B1(_10403_),
    .X(_10437_));
 sky130_fd_sc_hd__a211o_2 _18981_ (.A1(_10273_),
    .A2(_10275_),
    .B1(_10436_),
    .C1(_10437_),
    .X(_10438_));
 sky130_fd_sc_hd__o211ai_2 _18982_ (.A1(_10436_),
    .A2(_10437_),
    .B1(_10273_),
    .C1(_10275_),
    .Y(_10439_));
 sky130_fd_sc_hd__or4bb_4 _18983_ (.A(_10380_),
    .B(_10381_),
    .C_N(_10438_),
    .D_N(_10439_),
    .X(_10440_));
 sky130_fd_sc_hd__a2bb2o_1 _18984_ (.A1_N(_10380_),
    .A2_N(_10381_),
    .B1(_10438_),
    .B2(_10439_),
    .X(_10441_));
 sky130_fd_sc_hd__o211ai_4 _18985_ (.A1(_10277_),
    .A2(_10279_),
    .B1(_10440_),
    .C1(_10441_),
    .Y(_10442_));
 sky130_fd_sc_hd__a211o_1 _18986_ (.A1(_10440_),
    .A2(_10441_),
    .B1(_10277_),
    .C1(_10279_),
    .X(_10443_));
 sky130_fd_sc_hd__or4bb_2 _18987_ (.A(_10346_),
    .B(_10347_),
    .C_N(_10442_),
    .D_N(_10443_),
    .X(_10444_));
 sky130_fd_sc_hd__a2bb2o_1 _18988_ (.A1_N(_10346_),
    .A2_N(_10347_),
    .B1(_10442_),
    .B2(_10443_),
    .X(_10445_));
 sky130_fd_sc_hd__o211a_1 _18989_ (.A1(_10282_),
    .A2(_10284_),
    .B1(_10444_),
    .C1(_10445_),
    .X(_10446_));
 sky130_fd_sc_hd__a211oi_1 _18990_ (.A1(_10444_),
    .A2(_10445_),
    .B1(_10282_),
    .C1(_10284_),
    .Y(_10447_));
 sky130_fd_sc_hd__or3_1 _18991_ (.A(_10303_),
    .B(_10446_),
    .C(_10447_),
    .X(_10448_));
 sky130_fd_sc_hd__o21ai_1 _18992_ (.A1(_10446_),
    .A2(_10447_),
    .B1(_10303_),
    .Y(_10449_));
 sky130_fd_sc_hd__o211a_1 _18993_ (.A1(_10286_),
    .A2(_10288_),
    .B1(_10448_),
    .C1(_10449_),
    .X(_10450_));
 sky130_fd_sc_hd__a211oi_1 _18994_ (.A1(_10448_),
    .A2(_10449_),
    .B1(_10286_),
    .C1(_10288_),
    .Y(_10451_));
 sky130_fd_sc_hd__or3b_2 _18995_ (.A(_10450_),
    .B(_10451_),
    .C_N(_10164_),
    .X(_10452_));
 sky130_fd_sc_hd__o21bai_2 _18996_ (.A1(_10450_),
    .A2(_10451_),
    .B1_N(_10164_),
    .Y(_10453_));
 sky130_fd_sc_hd__nand2_1 _18997_ (.A(_10452_),
    .B(_10453_),
    .Y(_10454_));
 sky130_fd_sc_hd__a21oi_2 _18998_ (.A1(_10452_),
    .A2(_10453_),
    .B1(_10291_),
    .Y(_10455_));
 sky130_fd_sc_hd__and3_1 _18999_ (.A(_10291_),
    .B(_10452_),
    .C(_10453_),
    .X(_10456_));
 sky130_fd_sc_hd__nor2_2 _19000_ (.A(_10455_),
    .B(_10456_),
    .Y(_10457_));
 sky130_fd_sc_hd__xnor2_4 _19001_ (.A(_10302_),
    .B(_10457_),
    .Y(_10458_));
 sky130_fd_sc_hd__nor2_1 _19002_ (.A(_03049_),
    .B(_10458_),
    .Y(_10459_));
 sky130_fd_sc_hd__a221o_1 _19003_ (.A1(\temp[14] ),
    .A2(net7),
    .B1(_05615_),
    .B2(_03052_),
    .C1(_10459_),
    .X(_10460_));
 sky130_fd_sc_hd__mux2_1 _19004_ (.A0(net743),
    .A1(_10460_),
    .S(net4),
    .X(_00313_));
 sky130_fd_sc_hd__a21bo_1 _19005_ (.A1(_10304_),
    .A2(_10345_),
    .B1_N(_10344_),
    .X(_10461_));
 sky130_fd_sc_hd__nor2_1 _19006_ (.A(_10340_),
    .B(_10342_),
    .Y(_10462_));
 sky130_fd_sc_hd__nor2_2 _19007_ (.A(_10378_),
    .B(_10380_),
    .Y(_10463_));
 sky130_fd_sc_hd__and4b_1 _19008_ (.A_N(net321),
    .B(net65),
    .C(net62),
    .D(net316),
    .X(_10464_));
 sky130_fd_sc_hd__o2bb2a_1 _19009_ (.A1_N(net316),
    .A2_N(net65),
    .B1(net56),
    .B2(net321),
    .X(_10465_));
 sky130_fd_sc_hd__nor2_1 _19010_ (.A(_10464_),
    .B(_10465_),
    .Y(_10466_));
 sky130_fd_sc_hd__inv_2 _19011_ (.A(_10466_),
    .Y(_10467_));
 sky130_fd_sc_hd__a22o_1 _19012_ (.A1(net302),
    .A2(net74),
    .B1(net71),
    .B2(net307),
    .X(_10468_));
 sky130_fd_sc_hd__and3_1 _19013_ (.A(net302),
    .B(net307),
    .C(net74),
    .X(_10469_));
 sky130_fd_sc_hd__a21bo_1 _19014_ (.A1(net71),
    .A2(_10469_),
    .B1_N(_10468_),
    .X(_10470_));
 sky130_fd_sc_hd__nand2_1 _19015_ (.A(net311),
    .B(net68),
    .Y(_10471_));
 sky130_fd_sc_hd__xnor2_2 _19016_ (.A(_10470_),
    .B(_10471_),
    .Y(_10472_));
 sky130_fd_sc_hd__or2_1 _19017_ (.A(_10306_),
    .B(_10308_),
    .X(_10473_));
 sky130_fd_sc_hd__and2b_1 _19018_ (.A_N(_10472_),
    .B(_10473_),
    .X(_10474_));
 sky130_fd_sc_hd__xor2_2 _19019_ (.A(_10472_),
    .B(_10473_),
    .X(_10475_));
 sky130_fd_sc_hd__nor2_1 _19020_ (.A(_10467_),
    .B(_10475_),
    .Y(_10476_));
 sky130_fd_sc_hd__xnor2_2 _19021_ (.A(_10467_),
    .B(_10475_),
    .Y(_10477_));
 sky130_fd_sc_hd__a21oi_1 _19022_ (.A1(_10311_),
    .A2(_10319_),
    .B1(_10477_),
    .Y(_10478_));
 sky130_fd_sc_hd__a21o_1 _19023_ (.A1(_10311_),
    .A2(_10319_),
    .B1(_10477_),
    .X(_10479_));
 sky130_fd_sc_hd__nand3_1 _19024_ (.A(_10311_),
    .B(_10319_),
    .C(_10477_),
    .Y(_10480_));
 sky130_fd_sc_hd__o211a_1 _19025_ (.A1(_10314_),
    .A2(_10316_),
    .B1(_10479_),
    .C1(_10480_),
    .X(_10481_));
 sky130_fd_sc_hd__a211oi_2 _19026_ (.A1(_10479_),
    .A2(_10480_),
    .B1(_10314_),
    .C1(_10316_),
    .Y(_10482_));
 sky130_fd_sc_hd__a21o_1 _19027_ (.A1(_10352_),
    .A2(_10360_),
    .B1(_10359_),
    .X(_10483_));
 sky130_fd_sc_hd__nand2_1 _19028_ (.A(_10328_),
    .B(_10330_),
    .Y(_10484_));
 sky130_fd_sc_hd__a22o_1 _19029_ (.A1(net285),
    .A2(net81),
    .B1(net78),
    .B2(net291),
    .X(_10485_));
 sky130_fd_sc_hd__nand4_1 _19030_ (.A(net285),
    .B(net291),
    .C(net82),
    .D(\mul1.b[25] ),
    .Y(_10486_));
 sky130_fd_sc_hd__a22oi_2 _19031_ (.A1(net297),
    .A2(net75),
    .B1(_10485_),
    .B2(_10486_),
    .Y(_10487_));
 sky130_fd_sc_hd__and4_1 _19032_ (.A(net297),
    .B(net75),
    .C(_10485_),
    .D(_10486_),
    .X(_10488_));
 sky130_fd_sc_hd__a211o_1 _19033_ (.A1(_10349_),
    .A2(_10351_),
    .B1(_10487_),
    .C1(_10488_),
    .X(_10489_));
 sky130_fd_sc_hd__o211ai_2 _19034_ (.A1(_10487_),
    .A2(_10488_),
    .B1(_10349_),
    .C1(_10351_),
    .Y(_10490_));
 sky130_fd_sc_hd__nand3_2 _19035_ (.A(_10484_),
    .B(_10489_),
    .C(_10490_),
    .Y(_10491_));
 sky130_fd_sc_hd__a21o_1 _19036_ (.A1(_10489_),
    .A2(_10490_),
    .B1(_10484_),
    .X(_10492_));
 sky130_fd_sc_hd__and3_1 _19037_ (.A(_10483_),
    .B(_10491_),
    .C(_10492_),
    .X(_10493_));
 sky130_fd_sc_hd__a21oi_1 _19038_ (.A1(_10491_),
    .A2(_10492_),
    .B1(_10483_),
    .Y(_10494_));
 sky130_fd_sc_hd__a211o_1 _19039_ (.A1(_10331_),
    .A2(_10333_),
    .B1(_10493_),
    .C1(_10494_),
    .X(_10495_));
 sky130_fd_sc_hd__o211ai_2 _19040_ (.A1(_10493_),
    .A2(_10494_),
    .B1(_10331_),
    .C1(_10333_),
    .Y(_10496_));
 sky130_fd_sc_hd__o211a_1 _19041_ (.A1(_10335_),
    .A2(_10337_),
    .B1(_10495_),
    .C1(_10496_),
    .X(_10497_));
 sky130_fd_sc_hd__a211oi_2 _19042_ (.A1(_10495_),
    .A2(_10496_),
    .B1(_10335_),
    .C1(_10337_),
    .Y(_10498_));
 sky130_fd_sc_hd__nor4_2 _19043_ (.A(_10481_),
    .B(_10482_),
    .C(_10497_),
    .D(_10498_),
    .Y(_10499_));
 sky130_fd_sc_hd__o22a_1 _19044_ (.A1(_10481_),
    .A2(_10482_),
    .B1(_10497_),
    .B2(_10498_),
    .X(_10500_));
 sky130_fd_sc_hd__nor2_1 _19045_ (.A(_10499_),
    .B(_10500_),
    .Y(_10501_));
 sky130_fd_sc_hd__xnor2_2 _19046_ (.A(_10463_),
    .B(_10501_),
    .Y(_10502_));
 sky130_fd_sc_hd__nand2b_1 _19047_ (.A_N(_10462_),
    .B(_10502_),
    .Y(_10503_));
 sky130_fd_sc_hd__xnor2_2 _19048_ (.A(_10462_),
    .B(_10502_),
    .Y(_10504_));
 sky130_fd_sc_hd__and2b_1 _19049_ (.A_N(_10374_),
    .B(_10376_),
    .X(_10505_));
 sky130_fd_sc_hd__a22o_1 _19050_ (.A1(net270),
    .A2(net94),
    .B1(net89),
    .B2(net275),
    .X(_10506_));
 sky130_fd_sc_hd__and3_1 _19051_ (.A(net270),
    .B(net275),
    .C(net94),
    .X(_10507_));
 sky130_fd_sc_hd__a21bo_1 _19052_ (.A1(net89),
    .A2(_10507_),
    .B1_N(_10506_),
    .X(_10508_));
 sky130_fd_sc_hd__nand2_1 _19053_ (.A(net280),
    .B(net88),
    .Y(_10509_));
 sky130_fd_sc_hd__xor2_1 _19054_ (.A(_10508_),
    .B(_10509_),
    .X(_10510_));
 sky130_fd_sc_hd__a22o_1 _19055_ (.A1(net254),
    .A2(net109),
    .B1(net104),
    .B2(net259),
    .X(_10511_));
 sky130_fd_sc_hd__and4_1 _19056_ (.A(net253),
    .B(net259),
    .C(net108),
    .D(net103),
    .X(_10512_));
 sky130_fd_sc_hd__nand4_1 _19057_ (.A(net253),
    .B(net259),
    .C(net109),
    .D(net104),
    .Y(_10513_));
 sky130_fd_sc_hd__a22o_1 _19058_ (.A1(net264),
    .A2(net100),
    .B1(_10511_),
    .B2(_10513_),
    .X(_10514_));
 sky130_fd_sc_hd__and4_1 _19059_ (.A(net264),
    .B(net100),
    .C(_10511_),
    .D(_10513_),
    .X(_10515_));
 sky130_fd_sc_hd__nand4_1 _19060_ (.A(net264),
    .B(net100),
    .C(_10511_),
    .D(_10513_),
    .Y(_10516_));
 sky130_fd_sc_hd__o211a_1 _19061_ (.A1(_10354_),
    .A2(_10357_),
    .B1(_10514_),
    .C1(_10516_),
    .X(_10517_));
 sky130_fd_sc_hd__a211o_1 _19062_ (.A1(_10514_),
    .A2(_10516_),
    .B1(_10354_),
    .C1(_10357_),
    .X(_10518_));
 sky130_fd_sc_hd__nand2b_1 _19063_ (.A_N(_10517_),
    .B(_10518_),
    .Y(_10519_));
 sky130_fd_sc_hd__xnor2_1 _19064_ (.A(_10510_),
    .B(_10519_),
    .Y(_10520_));
 sky130_fd_sc_hd__nand2_1 _19065_ (.A(_10366_),
    .B(_10368_),
    .Y(_10521_));
 sky130_fd_sc_hd__a32o_1 _19066_ (.A1(net135),
    .A2(net238),
    .A3(_10385_),
    .B1(_10386_),
    .B2(net233),
    .X(_10522_));
 sky130_fd_sc_hd__a22o_1 _19067_ (.A1(net244),
    .A2(net124),
    .B1(net120),
    .B2(net627),
    .X(_10523_));
 sky130_fd_sc_hd__nand4_2 _19068_ (.A(net244),
    .B(net627),
    .C(net124),
    .D(net119),
    .Y(_10524_));
 sky130_fd_sc_hd__a22o_1 _19069_ (.A1(net249),
    .A2(net115),
    .B1(_10523_),
    .B2(_10524_),
    .X(_10525_));
 sky130_fd_sc_hd__nand4_2 _19070_ (.A(net249),
    .B(net115),
    .C(_10523_),
    .D(_10524_),
    .Y(_10526_));
 sky130_fd_sc_hd__nand3_1 _19071_ (.A(_10522_),
    .B(_10525_),
    .C(_10526_),
    .Y(_10527_));
 sky130_fd_sc_hd__a21o_1 _19072_ (.A1(_10525_),
    .A2(_10526_),
    .B1(_10522_),
    .X(_10528_));
 sky130_fd_sc_hd__nand3_1 _19073_ (.A(_10521_),
    .B(_10527_),
    .C(_10528_),
    .Y(_10529_));
 sky130_fd_sc_hd__a21o_1 _19074_ (.A1(_10527_),
    .A2(_10528_),
    .B1(_10521_),
    .X(_10530_));
 sky130_fd_sc_hd__a21bo_1 _19075_ (.A1(_10363_),
    .A2(_10370_),
    .B1_N(_10369_),
    .X(_10531_));
 sky130_fd_sc_hd__nand3_1 _19076_ (.A(_10529_),
    .B(_10530_),
    .C(_10531_),
    .Y(_10532_));
 sky130_fd_sc_hd__a21o_1 _19077_ (.A1(_10529_),
    .A2(_10530_),
    .B1(_10531_),
    .X(_10533_));
 sky130_fd_sc_hd__and3_1 _19078_ (.A(_10520_),
    .B(_10532_),
    .C(_10533_),
    .X(_10534_));
 sky130_fd_sc_hd__a21oi_1 _19079_ (.A1(_10532_),
    .A2(_10533_),
    .B1(_10520_),
    .Y(_10535_));
 sky130_fd_sc_hd__a211o_1 _19080_ (.A1(_10399_),
    .A2(_10401_),
    .B1(_10534_),
    .C1(_10535_),
    .X(_10536_));
 sky130_fd_sc_hd__o211ai_1 _19081_ (.A1(_10534_),
    .A2(_10535_),
    .B1(_10399_),
    .C1(_10401_),
    .Y(_10537_));
 sky130_fd_sc_hd__nand2_1 _19082_ (.A(_10536_),
    .B(_10537_),
    .Y(_10538_));
 sky130_fd_sc_hd__xor2_1 _19083_ (.A(_10505_),
    .B(_10538_),
    .X(_10539_));
 sky130_fd_sc_hd__nand2_1 _19084_ (.A(_10395_),
    .B(_10397_),
    .Y(_10540_));
 sky130_fd_sc_hd__a21o_1 _19085_ (.A1(_10404_),
    .A2(_10410_),
    .B1(_10409_),
    .X(_10541_));
 sky130_fd_sc_hd__a22o_1 _19086_ (.A1(net134),
    .A2(net234),
    .B1(net228),
    .B2(net139),
    .X(_10542_));
 sky130_fd_sc_hd__nand4_1 _19087_ (.A(net139),
    .B(net135),
    .C(net234),
    .D(net229),
    .Y(_10543_));
 sky130_fd_sc_hd__nand2_1 _19088_ (.A(_10542_),
    .B(_10543_),
    .Y(_10544_));
 sky130_fd_sc_hd__and2_1 _19089_ (.A(net130),
    .B(net238),
    .X(_10545_));
 sky130_fd_sc_hd__xnor2_1 _19090_ (.A(_10544_),
    .B(_10545_),
    .Y(_10546_));
 sky130_fd_sc_hd__a22o_1 _19091_ (.A1(net149),
    .A2(net219),
    .B1(net215),
    .B2(net154),
    .X(_10547_));
 sky130_fd_sc_hd__nand4_1 _19092_ (.A(net154),
    .B(net149),
    .C(net219),
    .D(net215),
    .Y(_10548_));
 sky130_fd_sc_hd__and2_1 _19093_ (.A(net143),
    .B(net224),
    .X(_10549_));
 sky130_fd_sc_hd__a21o_1 _19094_ (.A1(_10547_),
    .A2(_10548_),
    .B1(_10549_),
    .X(_10550_));
 sky130_fd_sc_hd__nand3_1 _19095_ (.A(_10547_),
    .B(_10548_),
    .C(_10549_),
    .Y(_10551_));
 sky130_fd_sc_hd__a21bo_1 _19096_ (.A1(_10389_),
    .A2(_10390_),
    .B1_N(_10391_),
    .X(_10552_));
 sky130_fd_sc_hd__nand3_2 _19097_ (.A(_10550_),
    .B(_10551_),
    .C(_10552_),
    .Y(_10553_));
 sky130_fd_sc_hd__a21o_1 _19098_ (.A1(_10550_),
    .A2(_10551_),
    .B1(_10552_),
    .X(_10554_));
 sky130_fd_sc_hd__nand3_2 _19099_ (.A(_10546_),
    .B(_10553_),
    .C(_10554_),
    .Y(_10555_));
 sky130_fd_sc_hd__a21o_1 _19100_ (.A1(_10553_),
    .A2(_10554_),
    .B1(_10546_),
    .X(_10556_));
 sky130_fd_sc_hd__nand3_2 _19101_ (.A(_10541_),
    .B(_10555_),
    .C(_10556_),
    .Y(_10557_));
 sky130_fd_sc_hd__a21o_1 _19102_ (.A1(_10555_),
    .A2(_10556_),
    .B1(_10541_),
    .X(_10558_));
 sky130_fd_sc_hd__nand3_2 _19103_ (.A(_10540_),
    .B(_10557_),
    .C(_10558_),
    .Y(_10559_));
 sky130_fd_sc_hd__a21o_1 _19104_ (.A1(_10557_),
    .A2(_10558_),
    .B1(_10540_),
    .X(_10560_));
 sky130_fd_sc_hd__and2_1 _19105_ (.A(_10559_),
    .B(_10560_),
    .X(_10561_));
 sky130_fd_sc_hd__nand2_1 _19106_ (.A(_10406_),
    .B(_10408_),
    .Y(_10562_));
 sky130_fd_sc_hd__a32o_1 _19107_ (.A1(net178),
    .A2(net202),
    .A3(_10414_),
    .B1(_10415_),
    .B2(net199),
    .X(_10563_));
 sky130_fd_sc_hd__a22o_1 _19108_ (.A1(net161),
    .A2(net209),
    .B1(net206),
    .B2(net167),
    .X(_10564_));
 sky130_fd_sc_hd__nand4_2 _19109_ (.A(net168),
    .B(net161),
    .C(net209),
    .D(net206),
    .Y(_10565_));
 sky130_fd_sc_hd__a22o_1 _19110_ (.A1(net156),
    .A2(net212),
    .B1(_10564_),
    .B2(_10565_),
    .X(_10566_));
 sky130_fd_sc_hd__nand4_1 _19111_ (.A(net156),
    .B(net212),
    .C(_10564_),
    .D(_10565_),
    .Y(_10567_));
 sky130_fd_sc_hd__and3_1 _19112_ (.A(_10563_),
    .B(_10566_),
    .C(_10567_),
    .X(_10568_));
 sky130_fd_sc_hd__a21o_1 _19113_ (.A1(_10566_),
    .A2(_10567_),
    .B1(_10563_),
    .X(_10569_));
 sky130_fd_sc_hd__and2b_1 _19114_ (.A_N(_10568_),
    .B(_10569_),
    .X(_10570_));
 sky130_fd_sc_hd__xor2_2 _19115_ (.A(_10562_),
    .B(_10570_),
    .X(_10571_));
 sky130_fd_sc_hd__a22o_1 _19116_ (.A1(net178),
    .A2(net199),
    .B1(net197),
    .B2(net183),
    .X(_10572_));
 sky130_fd_sc_hd__and3_1 _19117_ (.A(net183),
    .B(net178),
    .C(net197),
    .X(_10573_));
 sky130_fd_sc_hd__a21bo_1 _19118_ (.A1(net199),
    .A2(_10573_),
    .B1_N(_10572_),
    .X(_10574_));
 sky130_fd_sc_hd__nand2_1 _19119_ (.A(net173),
    .B(net202),
    .Y(_10575_));
 sky130_fd_sc_hd__xor2_1 _19120_ (.A(_10574_),
    .B(_10575_),
    .X(_10576_));
 sky130_fd_sc_hd__o21bai_1 _19121_ (.A1(_10418_),
    .A2(_10419_),
    .B1_N(_10420_),
    .Y(_10577_));
 sky130_fd_sc_hd__or2_1 _19122_ (.A(net623),
    .B(net190),
    .X(_10578_));
 sky130_fd_sc_hd__and3_1 _19123_ (.A(net623),
    .B(net190),
    .C(net193),
    .X(_10579_));
 sky130_fd_sc_hd__a21boi_1 _19124_ (.A1(net623),
    .A2(net190),
    .B1_N(net193),
    .Y(_10580_));
 sky130_fd_sc_hd__nand2_1 _19125_ (.A(\mul1.b[2] ),
    .B(net196),
    .Y(_10581_));
 sky130_fd_sc_hd__and3_4 _19126_ (.A(_10578_),
    .B(_10580_),
    .C(_10581_),
    .X(_10582_));
 sky130_fd_sc_hd__a21oi_1 _19127_ (.A1(_10578_),
    .A2(_10580_),
    .B1(_10581_),
    .Y(_10583_));
 sky130_fd_sc_hd__o21ai_1 _19128_ (.A1(_10582_),
    .A2(_10583_),
    .B1(_10577_),
    .Y(_10584_));
 sky130_fd_sc_hd__or3_1 _19129_ (.A(_10577_),
    .B(_10582_),
    .C(_10583_),
    .X(_10585_));
 sky130_fd_sc_hd__nand3_1 _19130_ (.A(_10576_),
    .B(_10584_),
    .C(_10585_),
    .Y(_10586_));
 sky130_fd_sc_hd__a21o_1 _19131_ (.A1(_10584_),
    .A2(_10585_),
    .B1(_10576_),
    .X(_10587_));
 sky130_fd_sc_hd__a21bo_1 _19132_ (.A1(_10417_),
    .A2(_10425_),
    .B1_N(_10424_),
    .X(_10588_));
 sky130_fd_sc_hd__nand3_1 _19133_ (.A(_10586_),
    .B(_10587_),
    .C(_10588_),
    .Y(_10589_));
 sky130_fd_sc_hd__a21o_1 _19134_ (.A1(_10586_),
    .A2(_10587_),
    .B1(_10588_),
    .X(_10590_));
 sky130_fd_sc_hd__and3_1 _19135_ (.A(_10571_),
    .B(_10589_),
    .C(_10590_),
    .X(_10591_));
 sky130_fd_sc_hd__a21oi_2 _19136_ (.A1(_10589_),
    .A2(_10590_),
    .B1(_10571_),
    .Y(_10592_));
 sky130_fd_sc_hd__a211o_2 _19137_ (.A1(_10429_),
    .A2(_10432_),
    .B1(_10591_),
    .C1(_10592_),
    .X(_10593_));
 sky130_fd_sc_hd__o211ai_4 _19138_ (.A1(_10591_),
    .A2(_10592_),
    .B1(_10429_),
    .C1(_10432_),
    .Y(_10594_));
 sky130_fd_sc_hd__nand3_2 _19139_ (.A(_10561_),
    .B(_10593_),
    .C(_10594_),
    .Y(_10595_));
 sky130_fd_sc_hd__a21o_1 _19140_ (.A1(_10593_),
    .A2(_10594_),
    .B1(_10561_),
    .X(_10596_));
 sky130_fd_sc_hd__o211ai_4 _19141_ (.A1(_10434_),
    .A2(_10436_),
    .B1(_10595_),
    .C1(_10596_),
    .Y(_10597_));
 sky130_fd_sc_hd__a211o_1 _19142_ (.A1(_10595_),
    .A2(_10596_),
    .B1(_10434_),
    .C1(_10436_),
    .X(_10598_));
 sky130_fd_sc_hd__and3_1 _19143_ (.A(_10539_),
    .B(_10597_),
    .C(_10598_),
    .X(_10599_));
 sky130_fd_sc_hd__a21oi_2 _19144_ (.A1(_10597_),
    .A2(_10598_),
    .B1(_10539_),
    .Y(_10600_));
 sky130_fd_sc_hd__a211oi_1 _19145_ (.A1(_10438_),
    .A2(_10440_),
    .B1(_10599_),
    .C1(_10600_),
    .Y(_10601_));
 sky130_fd_sc_hd__a211o_1 _19146_ (.A1(_10438_),
    .A2(_10440_),
    .B1(_10599_),
    .C1(_10600_),
    .X(_10602_));
 sky130_fd_sc_hd__o211ai_2 _19147_ (.A1(_10599_),
    .A2(_10600_),
    .B1(_10438_),
    .C1(_10440_),
    .Y(_10603_));
 sky130_fd_sc_hd__and3_1 _19148_ (.A(_10504_),
    .B(_10602_),
    .C(_10603_),
    .X(_10604_));
 sky130_fd_sc_hd__a21oi_1 _19149_ (.A1(_10602_),
    .A2(_10603_),
    .B1(_10504_),
    .Y(_10605_));
 sky130_fd_sc_hd__a211o_1 _19150_ (.A1(_10442_),
    .A2(_10444_),
    .B1(_10604_),
    .C1(_10605_),
    .X(_10606_));
 sky130_fd_sc_hd__o211ai_2 _19151_ (.A1(_10604_),
    .A2(_10605_),
    .B1(_10442_),
    .C1(_10444_),
    .Y(_10607_));
 sky130_fd_sc_hd__and3_1 _19152_ (.A(_10461_),
    .B(_10606_),
    .C(_10607_),
    .X(_10608_));
 sky130_fd_sc_hd__a21oi_1 _19153_ (.A1(_10606_),
    .A2(_10607_),
    .B1(_10461_),
    .Y(_10609_));
 sky130_fd_sc_hd__or2_1 _19154_ (.A(_10608_),
    .B(_10609_),
    .X(_10610_));
 sky130_fd_sc_hd__and2b_1 _19155_ (.A_N(_10446_),
    .B(_10448_),
    .X(_10611_));
 sky130_fd_sc_hd__nor2_1 _19156_ (.A(_10610_),
    .B(_10611_),
    .Y(_10612_));
 sky130_fd_sc_hd__xor2_2 _19157_ (.A(_10610_),
    .B(_10611_),
    .X(_10613_));
 sky130_fd_sc_hd__and2_1 _19158_ (.A(_10322_),
    .B(_10613_),
    .X(_10614_));
 sky130_fd_sc_hd__xnor2_1 _19159_ (.A(_10322_),
    .B(_10613_),
    .Y(_10615_));
 sky130_fd_sc_hd__and2b_1 _19160_ (.A_N(_10450_),
    .B(_10452_),
    .X(_10616_));
 sky130_fd_sc_hd__nor2_1 _19161_ (.A(_10615_),
    .B(_10616_),
    .Y(_10617_));
 sky130_fd_sc_hd__nand2_1 _19162_ (.A(_10615_),
    .B(_10616_),
    .Y(_10618_));
 sky130_fd_sc_hd__nand2b_2 _19163_ (.A_N(_10617_),
    .B(_10618_),
    .Y(_10619_));
 sky130_fd_sc_hd__o2111a_1 _19164_ (.A1(_10455_),
    .A2(_10456_),
    .B1(_09996_),
    .C1(_10146_),
    .D1(_10294_),
    .X(_10620_));
 sky130_fd_sc_hd__a21oi_1 _19165_ (.A1(_10291_),
    .A2(_10293_),
    .B1(_10454_),
    .Y(_10621_));
 sky130_fd_sc_hd__o211a_1 _19166_ (.A1(_10455_),
    .A2(_10456_),
    .B1(_10294_),
    .C1(_10296_),
    .X(_10622_));
 sky130_fd_sc_hd__a211o_1 _19167_ (.A1(_09856_),
    .A2(_10620_),
    .B1(_10621_),
    .C1(_10622_),
    .X(_10623_));
 sky130_fd_sc_hd__a31o_2 _19168_ (.A1(_09305_),
    .A2(_09854_),
    .A3(_10620_),
    .B1(_10623_),
    .X(_10624_));
 sky130_fd_sc_hd__xnor2_2 _19169_ (.A(_10619_),
    .B(_10624_),
    .Y(_10625_));
 sky130_fd_sc_hd__a22o_1 _19170_ (.A1(net764),
    .A2(net7),
    .B1(_05784_),
    .B2(_03052_),
    .X(_10626_));
 sky130_fd_sc_hd__a21o_1 _19171_ (.A1(net10),
    .A2(_10625_),
    .B1(_10626_),
    .X(_10627_));
 sky130_fd_sc_hd__mux2_1 _19172_ (.A0(net834),
    .A1(_10627_),
    .S(net4),
    .X(_00314_));
 sky130_fd_sc_hd__a21oi_1 _19173_ (.A1(_10618_),
    .A2(_10624_),
    .B1(_10617_),
    .Y(_10628_));
 sky130_fd_sc_hd__or2_1 _19174_ (.A(_10478_),
    .B(_10481_),
    .X(_10629_));
 sky130_fd_sc_hd__o31ai_2 _19175_ (.A1(_10463_),
    .A2(_10499_),
    .A3(_10500_),
    .B1(_10503_),
    .Y(_10630_));
 sky130_fd_sc_hd__nor2_1 _19176_ (.A(_10497_),
    .B(_10499_),
    .Y(_10631_));
 sky130_fd_sc_hd__o21ai_2 _19177_ (.A1(_10505_),
    .A2(_10538_),
    .B1(_10536_),
    .Y(_10632_));
 sky130_fd_sc_hd__a22o_1 _19178_ (.A1(net297),
    .A2(net74),
    .B1(net71),
    .B2(net302),
    .X(_10633_));
 sky130_fd_sc_hd__and3_1 _19179_ (.A(net297),
    .B(net302),
    .C(net71),
    .X(_10634_));
 sky130_fd_sc_hd__a21bo_2 _19180_ (.A1(net74),
    .A2(_10634_),
    .B1_N(_10633_),
    .X(_10635_));
 sky130_fd_sc_hd__nand2_2 _19181_ (.A(net307),
    .B(net68),
    .Y(_10636_));
 sky130_fd_sc_hd__xnor2_4 _19182_ (.A(_10635_),
    .B(_10636_),
    .Y(_10637_));
 sky130_fd_sc_hd__o2bb2a_2 _19183_ (.A1_N(net71),
    .A2_N(_10469_),
    .B1(_10470_),
    .B2(_10471_),
    .X(_10638_));
 sky130_fd_sc_hd__xnor2_2 _19184_ (.A(_10637_),
    .B(_10638_),
    .Y(_10639_));
 sky130_fd_sc_hd__and4b_2 _19185_ (.A_N(net317),
    .B(net65),
    .C(net62),
    .D(net311),
    .X(_10640_));
 sky130_fd_sc_hd__inv_2 _19186_ (.A(_10640_),
    .Y(_10641_));
 sky130_fd_sc_hd__o2bb2a_1 _19187_ (.A1_N(net311),
    .A2_N(net65),
    .B1(net56),
    .B2(net317),
    .X(_10642_));
 sky130_fd_sc_hd__nor2_1 _19188_ (.A(_10640_),
    .B(_10642_),
    .Y(_10643_));
 sky130_fd_sc_hd__xnor2_1 _19189_ (.A(_10639_),
    .B(_10643_),
    .Y(_10644_));
 sky130_fd_sc_hd__nor3_1 _19190_ (.A(_10474_),
    .B(_10476_),
    .C(_10644_),
    .Y(_10645_));
 sky130_fd_sc_hd__o21a_1 _19191_ (.A1(_10474_),
    .A2(_10476_),
    .B1(_10644_),
    .X(_10646_));
 sky130_fd_sc_hd__or2_1 _19192_ (.A(_10645_),
    .B(_10646_),
    .X(_10647_));
 sky130_fd_sc_hd__inv_2 _19193_ (.A(_10647_),
    .Y(_10648_));
 sky130_fd_sc_hd__xor2_1 _19194_ (.A(_10464_),
    .B(_10647_),
    .X(_10649_));
 sky130_fd_sc_hd__a21oi_1 _19195_ (.A1(_10510_),
    .A2(_10518_),
    .B1(_10517_),
    .Y(_10650_));
 sky130_fd_sc_hd__a41o_1 _19196_ (.A1(net285),
    .A2(net291),
    .A3(net81),
    .A4(\mul1.b[25] ),
    .B1(_10488_),
    .X(_10651_));
 sky130_fd_sc_hd__a32o_1 _19197_ (.A1(net280),
    .A2(net88),
    .A3(_10506_),
    .B1(_10507_),
    .B2(net90),
    .X(_10652_));
 sky130_fd_sc_hd__a22o_1 _19198_ (.A1(net280),
    .A2(net82),
    .B1(net78),
    .B2(net285),
    .X(_10653_));
 sky130_fd_sc_hd__nand4_2 _19199_ (.A(net280),
    .B(net285),
    .C(net81),
    .D(net78),
    .Y(_10654_));
 sky130_fd_sc_hd__a22o_1 _19200_ (.A1(net291),
    .A2(net75),
    .B1(_10653_),
    .B2(_10654_),
    .X(_10655_));
 sky130_fd_sc_hd__nand4_2 _19201_ (.A(net291),
    .B(net75),
    .C(_10653_),
    .D(_10654_),
    .Y(_10656_));
 sky130_fd_sc_hd__nand3_2 _19202_ (.A(_10652_),
    .B(_10655_),
    .C(_10656_),
    .Y(_10657_));
 sky130_fd_sc_hd__a21o_1 _19203_ (.A1(_10655_),
    .A2(_10656_),
    .B1(_10652_),
    .X(_10658_));
 sky130_fd_sc_hd__nand3_1 _19204_ (.A(_10651_),
    .B(_10657_),
    .C(_10658_),
    .Y(_10659_));
 sky130_fd_sc_hd__a21o_1 _19205_ (.A1(_10657_),
    .A2(_10658_),
    .B1(_10651_),
    .X(_10660_));
 sky130_fd_sc_hd__and3b_1 _19206_ (.A_N(_10650_),
    .B(_10659_),
    .C(_10660_),
    .X(_10661_));
 sky130_fd_sc_hd__a21boi_1 _19207_ (.A1(_10659_),
    .A2(_10660_),
    .B1_N(_10650_),
    .Y(_10662_));
 sky130_fd_sc_hd__a211oi_1 _19208_ (.A1(_10489_),
    .A2(_10491_),
    .B1(_10661_),
    .C1(_10662_),
    .Y(_10663_));
 sky130_fd_sc_hd__o211ai_1 _19209_ (.A1(_10661_),
    .A2(_10662_),
    .B1(_10489_),
    .C1(_10491_),
    .Y(_10664_));
 sky130_fd_sc_hd__nand2b_1 _19210_ (.A_N(_10663_),
    .B(_10664_),
    .Y(_10665_));
 sky130_fd_sc_hd__and2b_1 _19211_ (.A_N(_10493_),
    .B(_10495_),
    .X(_10666_));
 sky130_fd_sc_hd__nor2_1 _19212_ (.A(_10665_),
    .B(_10666_),
    .Y(_10667_));
 sky130_fd_sc_hd__xnor2_1 _19213_ (.A(_10665_),
    .B(_10666_),
    .Y(_10668_));
 sky130_fd_sc_hd__xnor2_1 _19214_ (.A(_10649_),
    .B(_10668_),
    .Y(_10669_));
 sky130_fd_sc_hd__and2b_1 _19215_ (.A_N(_10669_),
    .B(_10632_),
    .X(_10670_));
 sky130_fd_sc_hd__xnor2_1 _19216_ (.A(_10632_),
    .B(_10669_),
    .Y(_10671_));
 sky130_fd_sc_hd__and2b_1 _19217_ (.A_N(_10631_),
    .B(_10671_),
    .X(_10672_));
 sky130_fd_sc_hd__xnor2_1 _19218_ (.A(_10631_),
    .B(_10671_),
    .Y(_10673_));
 sky130_fd_sc_hd__a31o_1 _19219_ (.A1(_10529_),
    .A2(_10530_),
    .A3(_10531_),
    .B1(_10534_),
    .X(_10674_));
 sky130_fd_sc_hd__a22o_1 _19220_ (.A1(net264),
    .A2(net93),
    .B1(net89),
    .B2(net269),
    .X(_10675_));
 sky130_fd_sc_hd__and3_1 _19221_ (.A(net264),
    .B(net269),
    .C(net89),
    .X(_10676_));
 sky130_fd_sc_hd__a21bo_1 _19222_ (.A1(net93),
    .A2(_10676_),
    .B1_N(_10675_),
    .X(_10677_));
 sky130_fd_sc_hd__nand2_1 _19223_ (.A(net275),
    .B(net85),
    .Y(_10678_));
 sky130_fd_sc_hd__xor2_1 _19224_ (.A(_10677_),
    .B(_10678_),
    .X(_10679_));
 sky130_fd_sc_hd__a22o_1 _19225_ (.A1(net249),
    .A2(net108),
    .B1(net103),
    .B2(net254),
    .X(_10680_));
 sky130_fd_sc_hd__and4_1 _19226_ (.A(net248),
    .B(net254),
    .C(net108),
    .D(net103),
    .X(_10681_));
 sky130_fd_sc_hd__nand4_1 _19227_ (.A(net249),
    .B(net254),
    .C(net108),
    .D(net103),
    .Y(_10682_));
 sky130_fd_sc_hd__a22o_1 _19228_ (.A1(net260),
    .A2(net99),
    .B1(_10680_),
    .B2(_10682_),
    .X(_10683_));
 sky130_fd_sc_hd__and4_1 _19229_ (.A(net260),
    .B(net99),
    .C(_10680_),
    .D(_10682_),
    .X(_10684_));
 sky130_fd_sc_hd__nand4_1 _19230_ (.A(net260),
    .B(net99),
    .C(_10680_),
    .D(_10682_),
    .Y(_10685_));
 sky130_fd_sc_hd__o211a_1 _19231_ (.A1(_10512_),
    .A2(_10515_),
    .B1(_10683_),
    .C1(_10685_),
    .X(_10686_));
 sky130_fd_sc_hd__a211o_1 _19232_ (.A1(_10683_),
    .A2(_10685_),
    .B1(_10512_),
    .C1(_10515_),
    .X(_10687_));
 sky130_fd_sc_hd__nand2b_1 _19233_ (.A_N(_10686_),
    .B(_10687_),
    .Y(_10688_));
 sky130_fd_sc_hd__xnor2_1 _19234_ (.A(_10679_),
    .B(_10688_),
    .Y(_10689_));
 sky130_fd_sc_hd__nand2_1 _19235_ (.A(_10524_),
    .B(_10526_),
    .Y(_10690_));
 sky130_fd_sc_hd__a21bo_1 _19236_ (.A1(_10542_),
    .A2(_10545_),
    .B1_N(_10543_),
    .X(_10691_));
 sky130_fd_sc_hd__a22o_1 _19237_ (.A1(net244),
    .A2(net119),
    .B1(net239),
    .B2(net124),
    .X(_10692_));
 sky130_fd_sc_hd__nand4_2 _19238_ (.A(net244),
    .B(net125),
    .C(net119),
    .D(net239),
    .Y(_10693_));
 sky130_fd_sc_hd__a22o_1 _19239_ (.A1(net627),
    .A2(net116),
    .B1(_10692_),
    .B2(_10693_),
    .X(_10694_));
 sky130_fd_sc_hd__nand4_2 _19240_ (.A(net627),
    .B(net115),
    .C(_10692_),
    .D(_10693_),
    .Y(_10695_));
 sky130_fd_sc_hd__nand3_1 _19241_ (.A(_10691_),
    .B(_10694_),
    .C(_10695_),
    .Y(_10696_));
 sky130_fd_sc_hd__a21o_1 _19242_ (.A1(_10694_),
    .A2(_10695_),
    .B1(_10691_),
    .X(_10697_));
 sky130_fd_sc_hd__nand3_1 _19243_ (.A(_10690_),
    .B(_10696_),
    .C(_10697_),
    .Y(_10698_));
 sky130_fd_sc_hd__a21o_1 _19244_ (.A1(_10696_),
    .A2(_10697_),
    .B1(_10690_),
    .X(_10699_));
 sky130_fd_sc_hd__a21bo_1 _19245_ (.A1(_10521_),
    .A2(_10528_),
    .B1_N(_10527_),
    .X(_10700_));
 sky130_fd_sc_hd__nand3_1 _19246_ (.A(_10698_),
    .B(_10699_),
    .C(_10700_),
    .Y(_10701_));
 sky130_fd_sc_hd__a21o_1 _19247_ (.A1(_10698_),
    .A2(_10699_),
    .B1(_10700_),
    .X(_10702_));
 sky130_fd_sc_hd__and3_1 _19248_ (.A(_10689_),
    .B(_10701_),
    .C(_10702_),
    .X(_10703_));
 sky130_fd_sc_hd__a21oi_1 _19249_ (.A1(_10701_),
    .A2(_10702_),
    .B1(_10689_),
    .Y(_10704_));
 sky130_fd_sc_hd__a211o_1 _19250_ (.A1(_10557_),
    .A2(_10559_),
    .B1(_10703_),
    .C1(_10704_),
    .X(_10705_));
 sky130_fd_sc_hd__o211ai_2 _19251_ (.A1(_10703_),
    .A2(_10704_),
    .B1(_10557_),
    .C1(_10559_),
    .Y(_10706_));
 sky130_fd_sc_hd__and3_1 _19252_ (.A(_10674_),
    .B(_10705_),
    .C(_10706_),
    .X(_10707_));
 sky130_fd_sc_hd__a21oi_1 _19253_ (.A1(_10705_),
    .A2(_10706_),
    .B1(_10674_),
    .Y(_10708_));
 sky130_fd_sc_hd__nor2_1 _19254_ (.A(_10707_),
    .B(_10708_),
    .Y(_10709_));
 sky130_fd_sc_hd__a21o_1 _19255_ (.A1(_10562_),
    .A2(_10569_),
    .B1(_10568_),
    .X(_10710_));
 sky130_fd_sc_hd__a22o_1 _19256_ (.A1(net134),
    .A2(net229),
    .B1(net225),
    .B2(net139),
    .X(_10711_));
 sky130_fd_sc_hd__nand4_1 _19257_ (.A(net139),
    .B(net134),
    .C(net229),
    .D(net224),
    .Y(_10712_));
 sky130_fd_sc_hd__nand2_1 _19258_ (.A(_10711_),
    .B(_10712_),
    .Y(_10713_));
 sky130_fd_sc_hd__and2_1 _19259_ (.A(net130),
    .B(net234),
    .X(_10714_));
 sky130_fd_sc_hd__xnor2_1 _19260_ (.A(_10713_),
    .B(_10714_),
    .Y(_10715_));
 sky130_fd_sc_hd__a22o_1 _19261_ (.A1(net148),
    .A2(net215),
    .B1(net211),
    .B2(net153),
    .X(_10716_));
 sky130_fd_sc_hd__nand4_4 _19262_ (.A(net153),
    .B(net148),
    .C(net215),
    .D(net211),
    .Y(_10717_));
 sky130_fd_sc_hd__a22o_1 _19263_ (.A1(net143),
    .A2(net220),
    .B1(_10716_),
    .B2(_10717_),
    .X(_10718_));
 sky130_fd_sc_hd__nand4_2 _19264_ (.A(net143),
    .B(net220),
    .C(_10716_),
    .D(_10717_),
    .Y(_10719_));
 sky130_fd_sc_hd__a21bo_1 _19265_ (.A1(_10547_),
    .A2(_10549_),
    .B1_N(_10548_),
    .X(_10720_));
 sky130_fd_sc_hd__nand3_1 _19266_ (.A(_10718_),
    .B(_10719_),
    .C(_10720_),
    .Y(_10721_));
 sky130_fd_sc_hd__a21o_1 _19267_ (.A1(_10718_),
    .A2(_10719_),
    .B1(_10720_),
    .X(_10722_));
 sky130_fd_sc_hd__nand3_1 _19268_ (.A(_10715_),
    .B(_10721_),
    .C(_10722_),
    .Y(_10723_));
 sky130_fd_sc_hd__a21o_1 _19269_ (.A1(_10721_),
    .A2(_10722_),
    .B1(_10715_),
    .X(_10724_));
 sky130_fd_sc_hd__and3_1 _19270_ (.A(_10710_),
    .B(_10723_),
    .C(_10724_),
    .X(_10725_));
 sky130_fd_sc_hd__nand3_1 _19271_ (.A(_10710_),
    .B(_10723_),
    .C(_10724_),
    .Y(_10726_));
 sky130_fd_sc_hd__a21oi_1 _19272_ (.A1(_10723_),
    .A2(_10724_),
    .B1(_10710_),
    .Y(_10727_));
 sky130_fd_sc_hd__a211o_1 _19273_ (.A1(_10553_),
    .A2(_10555_),
    .B1(_10725_),
    .C1(_10727_),
    .X(_10728_));
 sky130_fd_sc_hd__o211ai_1 _19274_ (.A1(_10725_),
    .A2(_10727_),
    .B1(_10553_),
    .C1(_10555_),
    .Y(_10729_));
 sky130_fd_sc_hd__and2_1 _19275_ (.A(_10728_),
    .B(_10729_),
    .X(_10730_));
 sky130_fd_sc_hd__nand2_1 _19276_ (.A(_10565_),
    .B(_10567_),
    .Y(_10731_));
 sky130_fd_sc_hd__a32o_1 _19277_ (.A1(net173),
    .A2(net202),
    .A3(_10572_),
    .B1(_10573_),
    .B2(net199),
    .X(_10732_));
 sky130_fd_sc_hd__a22o_1 _19278_ (.A1(net161),
    .A2(net206),
    .B1(net202),
    .B2(net168),
    .X(_10733_));
 sky130_fd_sc_hd__nand4_2 _19279_ (.A(net168),
    .B(net161),
    .C(net206),
    .D(net202),
    .Y(_10734_));
 sky130_fd_sc_hd__a22o_1 _19280_ (.A1(net156),
    .A2(net209),
    .B1(_10733_),
    .B2(_10734_),
    .X(_10735_));
 sky130_fd_sc_hd__nand4_2 _19281_ (.A(net156),
    .B(net209),
    .C(_10733_),
    .D(_10734_),
    .Y(_10736_));
 sky130_fd_sc_hd__and3_1 _19282_ (.A(_10732_),
    .B(_10735_),
    .C(_10736_),
    .X(_10737_));
 sky130_fd_sc_hd__a21o_1 _19283_ (.A1(_10735_),
    .A2(_10736_),
    .B1(_10732_),
    .X(_10738_));
 sky130_fd_sc_hd__and2b_1 _19284_ (.A_N(_10737_),
    .B(_10738_),
    .X(_10739_));
 sky130_fd_sc_hd__xnor2_2 _19285_ (.A(_10731_),
    .B(_10739_),
    .Y(_10740_));
 sky130_fd_sc_hd__a22o_1 _19286_ (.A1(net178),
    .A2(net197),
    .B1(net195),
    .B2(net183),
    .X(_10741_));
 sky130_fd_sc_hd__a21bo_1 _19287_ (.A1(net195),
    .A2(_10573_),
    .B1_N(_10741_),
    .X(_10742_));
 sky130_fd_sc_hd__nand2_1 _19288_ (.A(net173),
    .B(net199),
    .Y(_10743_));
 sky130_fd_sc_hd__xor2_2 _19289_ (.A(_10742_),
    .B(_10743_),
    .X(_10744_));
 sky130_fd_sc_hd__mux2_4 _19290_ (.A0(_10579_),
    .A1(_10580_),
    .S(net187),
    .X(_10745_));
 sky130_fd_sc_hd__xor2_2 _19291_ (.A(_10582_),
    .B(_10745_),
    .X(_10746_));
 sky130_fd_sc_hd__xnor2_2 _19292_ (.A(_10744_),
    .B(_10746_),
    .Y(_10747_));
 sky130_fd_sc_hd__a21bo_1 _19293_ (.A1(_10576_),
    .A2(_10585_),
    .B1_N(_10584_),
    .X(_10748_));
 sky130_fd_sc_hd__nand2b_1 _19294_ (.A_N(_10747_),
    .B(_10748_),
    .Y(_10749_));
 sky130_fd_sc_hd__xor2_2 _19295_ (.A(_10747_),
    .B(_10748_),
    .X(_10750_));
 sky130_fd_sc_hd__xnor2_2 _19296_ (.A(_10740_),
    .B(_10750_),
    .Y(_10751_));
 sky130_fd_sc_hd__a21bo_1 _19297_ (.A1(_10571_),
    .A2(_10590_),
    .B1_N(_10589_),
    .X(_10752_));
 sky130_fd_sc_hd__and2b_1 _19298_ (.A_N(_10751_),
    .B(_10752_),
    .X(_10753_));
 sky130_fd_sc_hd__xnor2_2 _19299_ (.A(_10751_),
    .B(_10752_),
    .Y(_10754_));
 sky130_fd_sc_hd__xnor2_2 _19300_ (.A(_10730_),
    .B(_10754_),
    .Y(_10755_));
 sky130_fd_sc_hd__a21bo_1 _19301_ (.A1(_10561_),
    .A2(_10594_),
    .B1_N(_10593_),
    .X(_10756_));
 sky130_fd_sc_hd__and2b_1 _19302_ (.A_N(_10755_),
    .B(_10756_),
    .X(_10757_));
 sky130_fd_sc_hd__xnor2_2 _19303_ (.A(_10755_),
    .B(_10756_),
    .Y(_10758_));
 sky130_fd_sc_hd__xnor2_2 _19304_ (.A(_10709_),
    .B(_10758_),
    .Y(_10759_));
 sky130_fd_sc_hd__a21bo_1 _19305_ (.A1(_10539_),
    .A2(_10598_),
    .B1_N(_10597_),
    .X(_10760_));
 sky130_fd_sc_hd__and2b_1 _19306_ (.A_N(_10759_),
    .B(_10760_),
    .X(_10761_));
 sky130_fd_sc_hd__xnor2_2 _19307_ (.A(_10759_),
    .B(_10760_),
    .Y(_10762_));
 sky130_fd_sc_hd__xor2_1 _19308_ (.A(_10673_),
    .B(_10762_),
    .X(_10763_));
 sky130_fd_sc_hd__a21oi_2 _19309_ (.A1(_10504_),
    .A2(_10603_),
    .B1(_10601_),
    .Y(_10764_));
 sky130_fd_sc_hd__nand2b_1 _19310_ (.A_N(_10764_),
    .B(_10763_),
    .Y(_10765_));
 sky130_fd_sc_hd__xnor2_1 _19311_ (.A(_10763_),
    .B(_10764_),
    .Y(_10766_));
 sky130_fd_sc_hd__nand2_1 _19312_ (.A(_10630_),
    .B(_10766_),
    .Y(_10767_));
 sky130_fd_sc_hd__xnor2_1 _19313_ (.A(_10630_),
    .B(_10766_),
    .Y(_10768_));
 sky130_fd_sc_hd__a21boi_1 _19314_ (.A1(_10461_),
    .A2(_10607_),
    .B1_N(_10606_),
    .Y(_10769_));
 sky130_fd_sc_hd__nor2_1 _19315_ (.A(_10768_),
    .B(_10769_),
    .Y(_10770_));
 sky130_fd_sc_hd__and2_1 _19316_ (.A(_10768_),
    .B(_10769_),
    .X(_10771_));
 sky130_fd_sc_hd__nor2_1 _19317_ (.A(_10770_),
    .B(_10771_),
    .Y(_10772_));
 sky130_fd_sc_hd__xor2_1 _19318_ (.A(_10629_),
    .B(_10772_),
    .X(_10773_));
 sky130_fd_sc_hd__o21a_1 _19319_ (.A1(_10612_),
    .A2(_10614_),
    .B1(_10773_),
    .X(_10774_));
 sky130_fd_sc_hd__or3_1 _19320_ (.A(_10612_),
    .B(_10614_),
    .C(_10773_),
    .X(_10775_));
 sky130_fd_sc_hd__nand2b_2 _19321_ (.A_N(_10774_),
    .B(_10775_),
    .Y(_10776_));
 sky130_fd_sc_hd__xnor2_2 _19322_ (.A(_10628_),
    .B(_10776_),
    .Y(_10777_));
 sky130_fd_sc_hd__o2bb2a_1 _19323_ (.A1_N(\temp[16] ),
    .A2_N(net7),
    .B1(_05935_),
    .B2(net44),
    .X(_10778_));
 sky130_fd_sc_hd__o21ai_1 _19324_ (.A1(_03049_),
    .A2(_10777_),
    .B1(_10778_),
    .Y(_10779_));
 sky130_fd_sc_hd__mux2_1 _19325_ (.A0(net898),
    .A1(_10779_),
    .S(net3),
    .X(_00315_));
 sky130_fd_sc_hd__a21o_1 _19326_ (.A1(_10464_),
    .A2(_10648_),
    .B1(_10646_),
    .X(_10780_));
 sky130_fd_sc_hd__or2_1 _19327_ (.A(_10670_),
    .B(_10672_),
    .X(_10781_));
 sky130_fd_sc_hd__o21ba_1 _19328_ (.A1(_10649_),
    .A2(_10668_),
    .B1_N(_10667_),
    .X(_10782_));
 sky130_fd_sc_hd__a21bo_1 _19329_ (.A1(_10674_),
    .A2(_10706_),
    .B1_N(_10705_),
    .X(_10783_));
 sky130_fd_sc_hd__a22o_1 _19330_ (.A1(net291),
    .A2(net73),
    .B1(net70),
    .B2(net297),
    .X(_10784_));
 sky130_fd_sc_hd__and3_1 _19331_ (.A(net290),
    .B(net297),
    .C(net70),
    .X(_10785_));
 sky130_fd_sc_hd__a21bo_1 _19332_ (.A1(net73),
    .A2(_10785_),
    .B1_N(_10784_),
    .X(_10786_));
 sky130_fd_sc_hd__nand2_1 _19333_ (.A(net302),
    .B(net67),
    .Y(_10787_));
 sky130_fd_sc_hd__xnor2_2 _19334_ (.A(_10786_),
    .B(_10787_),
    .Y(_10788_));
 sky130_fd_sc_hd__o2bb2a_2 _19335_ (.A1_N(net74),
    .A2_N(_10634_),
    .B1(_10635_),
    .B2(_10636_),
    .X(_10789_));
 sky130_fd_sc_hd__xnor2_2 _19336_ (.A(_10788_),
    .B(_10789_),
    .Y(_00520_));
 sky130_fd_sc_hd__and4b_2 _19337_ (.A_N(net311),
    .B(net64),
    .C(net62),
    .D(net307),
    .X(_00521_));
 sky130_fd_sc_hd__inv_2 _19338_ (.A(_00521_),
    .Y(_00522_));
 sky130_fd_sc_hd__o2bb2a_1 _19339_ (.A1_N(net306),
    .A2_N(net64),
    .B1(net56),
    .B2(net312),
    .X(_00523_));
 sky130_fd_sc_hd__nor2_1 _19340_ (.A(_00521_),
    .B(_00523_),
    .Y(_00524_));
 sky130_fd_sc_hd__xnor2_1 _19341_ (.A(_00520_),
    .B(_00524_),
    .Y(_00525_));
 sky130_fd_sc_hd__o32ai_4 _19342_ (.A1(_10639_),
    .A2(_10640_),
    .A3(_10642_),
    .B1(_10638_),
    .B2(_10637_),
    .Y(_00526_));
 sky130_fd_sc_hd__xnor2_1 _19343_ (.A(_00525_),
    .B(_00526_),
    .Y(_00527_));
 sky130_fd_sc_hd__nor2_1 _19344_ (.A(_10641_),
    .B(_00527_),
    .Y(_00528_));
 sky130_fd_sc_hd__and2_1 _19345_ (.A(_10641_),
    .B(_00527_),
    .X(_00529_));
 sky130_fd_sc_hd__or2_1 _19346_ (.A(_00528_),
    .B(_00529_),
    .X(_00530_));
 sky130_fd_sc_hd__a21oi_1 _19347_ (.A1(_10679_),
    .A2(_10687_),
    .B1(_10686_),
    .Y(_00531_));
 sky130_fd_sc_hd__nand2_1 _19348_ (.A(_10654_),
    .B(_10656_),
    .Y(_00532_));
 sky130_fd_sc_hd__a32o_1 _19349_ (.A1(net275),
    .A2(net85),
    .A3(_10675_),
    .B1(_10676_),
    .B2(net96),
    .X(_00533_));
 sky130_fd_sc_hd__a22o_1 _19350_ (.A1(net275),
    .A2(net84),
    .B1(net80),
    .B2(net280),
    .X(_00534_));
 sky130_fd_sc_hd__nand4_2 _19351_ (.A(net275),
    .B(net280),
    .C(net84),
    .D(net80),
    .Y(_00535_));
 sky130_fd_sc_hd__a22o_1 _19352_ (.A1(net285),
    .A2(net77),
    .B1(_00534_),
    .B2(_00535_),
    .X(_00536_));
 sky130_fd_sc_hd__nand4_2 _19353_ (.A(net285),
    .B(net77),
    .C(_00534_),
    .D(_00535_),
    .Y(_00537_));
 sky130_fd_sc_hd__nand3_2 _19354_ (.A(_00533_),
    .B(_00536_),
    .C(_00537_),
    .Y(_00538_));
 sky130_fd_sc_hd__a21o_1 _19355_ (.A1(_00536_),
    .A2(_00537_),
    .B1(_00533_),
    .X(_00539_));
 sky130_fd_sc_hd__nand3_1 _19356_ (.A(_00532_),
    .B(_00538_),
    .C(_00539_),
    .Y(_00540_));
 sky130_fd_sc_hd__a21o_1 _19357_ (.A1(_00538_),
    .A2(_00539_),
    .B1(_00532_),
    .X(_00541_));
 sky130_fd_sc_hd__and3b_1 _19358_ (.A_N(_00531_),
    .B(_00540_),
    .C(_00541_),
    .X(_00542_));
 sky130_fd_sc_hd__a21boi_1 _19359_ (.A1(_00540_),
    .A2(_00541_),
    .B1_N(_00531_),
    .Y(_00543_));
 sky130_fd_sc_hd__a211oi_1 _19360_ (.A1(_10657_),
    .A2(_10659_),
    .B1(_00542_),
    .C1(_00543_),
    .Y(_00544_));
 sky130_fd_sc_hd__o211ai_1 _19361_ (.A1(_00542_),
    .A2(_00543_),
    .B1(_10657_),
    .C1(_10659_),
    .Y(_00545_));
 sky130_fd_sc_hd__nand2b_1 _19362_ (.A_N(_00544_),
    .B(_00545_),
    .Y(_00546_));
 sky130_fd_sc_hd__nor2_1 _19363_ (.A(_10661_),
    .B(_10663_),
    .Y(_00547_));
 sky130_fd_sc_hd__nor2_1 _19364_ (.A(_00546_),
    .B(_00547_),
    .Y(_00548_));
 sky130_fd_sc_hd__xnor2_1 _19365_ (.A(_00546_),
    .B(_00547_),
    .Y(_00549_));
 sky130_fd_sc_hd__xnor2_1 _19366_ (.A(_00530_),
    .B(_00549_),
    .Y(_00550_));
 sky130_fd_sc_hd__and2b_1 _19367_ (.A_N(_00550_),
    .B(_10783_),
    .X(_00551_));
 sky130_fd_sc_hd__xnor2_1 _19368_ (.A(_10783_),
    .B(_00550_),
    .Y(_00552_));
 sky130_fd_sc_hd__and2b_1 _19369_ (.A_N(_10782_),
    .B(_00552_),
    .X(_00553_));
 sky130_fd_sc_hd__xnor2_1 _19370_ (.A(_10782_),
    .B(_00552_),
    .Y(_00554_));
 sky130_fd_sc_hd__a31o_1 _19371_ (.A1(_10698_),
    .A2(_10699_),
    .A3(_10700_),
    .B1(_10703_),
    .X(_00555_));
 sky130_fd_sc_hd__a22o_1 _19372_ (.A1(net259),
    .A2(net95),
    .B1(net92),
    .B2(net266),
    .X(_00556_));
 sky130_fd_sc_hd__and3_1 _19373_ (.A(net259),
    .B(net264),
    .C(net92),
    .X(_00557_));
 sky130_fd_sc_hd__a21bo_1 _19374_ (.A1(net95),
    .A2(_00557_),
    .B1_N(_00556_),
    .X(_00558_));
 sky130_fd_sc_hd__nand2_1 _19375_ (.A(net271),
    .B(net87),
    .Y(_00559_));
 sky130_fd_sc_hd__xor2_1 _19376_ (.A(_00558_),
    .B(_00559_),
    .X(_00560_));
 sky130_fd_sc_hd__a22o_1 _19377_ (.A1(net627),
    .A2(net110),
    .B1(net105),
    .B2(net248),
    .X(_00561_));
 sky130_fd_sc_hd__and4_1 _19378_ (.A(net627),
    .B(net249),
    .C(net110),
    .D(net106),
    .X(_00562_));
 sky130_fd_sc_hd__nand4_1 _19379_ (.A(net627),
    .B(net249),
    .C(net110),
    .D(net105),
    .Y(_00563_));
 sky130_fd_sc_hd__a22o_1 _19380_ (.A1(net254),
    .A2(net99),
    .B1(_00561_),
    .B2(_00563_),
    .X(_00564_));
 sky130_fd_sc_hd__and4_1 _19381_ (.A(net254),
    .B(net101),
    .C(_00561_),
    .D(_00563_),
    .X(_00565_));
 sky130_fd_sc_hd__nand4_1 _19382_ (.A(net254),
    .B(net99),
    .C(_00561_),
    .D(_00563_),
    .Y(_00566_));
 sky130_fd_sc_hd__o211a_1 _19383_ (.A1(_10681_),
    .A2(_10684_),
    .B1(_00564_),
    .C1(_00566_),
    .X(_00567_));
 sky130_fd_sc_hd__a211o_1 _19384_ (.A1(_00564_),
    .A2(_00566_),
    .B1(_10681_),
    .C1(_10684_),
    .X(_00568_));
 sky130_fd_sc_hd__nand2b_1 _19385_ (.A_N(_00567_),
    .B(_00568_),
    .Y(_00569_));
 sky130_fd_sc_hd__xnor2_1 _19386_ (.A(_00560_),
    .B(_00569_),
    .Y(_00570_));
 sky130_fd_sc_hd__nand2_1 _19387_ (.A(_10693_),
    .B(_10695_),
    .Y(_00571_));
 sky130_fd_sc_hd__a21bo_1 _19388_ (.A1(_10711_),
    .A2(_10714_),
    .B1_N(_10712_),
    .X(_00572_));
 sky130_fd_sc_hd__a22o_1 _19389_ (.A1(net120),
    .A2(net239),
    .B1(net234),
    .B2(net125),
    .X(_00573_));
 sky130_fd_sc_hd__nand4_2 _19390_ (.A(net125),
    .B(net120),
    .C(net239),
    .D(net234),
    .Y(_00574_));
 sky130_fd_sc_hd__a22o_1 _19391_ (.A1(net244),
    .A2(net116),
    .B1(_00573_),
    .B2(_00574_),
    .X(_00575_));
 sky130_fd_sc_hd__nand4_2 _19392_ (.A(net244),
    .B(net116),
    .C(_00573_),
    .D(_00574_),
    .Y(_00576_));
 sky130_fd_sc_hd__nand3_1 _19393_ (.A(_00572_),
    .B(_00575_),
    .C(_00576_),
    .Y(_00577_));
 sky130_fd_sc_hd__a21o_1 _19394_ (.A1(_00575_),
    .A2(_00576_),
    .B1(_00572_),
    .X(_00578_));
 sky130_fd_sc_hd__nand3_1 _19395_ (.A(_00571_),
    .B(_00577_),
    .C(_00578_),
    .Y(_00579_));
 sky130_fd_sc_hd__a21o_1 _19396_ (.A1(_00577_),
    .A2(_00578_),
    .B1(_00571_),
    .X(_00580_));
 sky130_fd_sc_hd__a21bo_1 _19397_ (.A1(_10690_),
    .A2(_10697_),
    .B1_N(_10696_),
    .X(_00581_));
 sky130_fd_sc_hd__nand3_1 _19398_ (.A(_00579_),
    .B(_00580_),
    .C(_00581_),
    .Y(_00582_));
 sky130_fd_sc_hd__a21o_1 _19399_ (.A1(_00579_),
    .A2(_00580_),
    .B1(_00581_),
    .X(_00583_));
 sky130_fd_sc_hd__and3_1 _19400_ (.A(_00570_),
    .B(_00582_),
    .C(_00583_),
    .X(_00584_));
 sky130_fd_sc_hd__a21oi_1 _19401_ (.A1(_00582_),
    .A2(_00583_),
    .B1(_00570_),
    .Y(_00585_));
 sky130_fd_sc_hd__a211oi_1 _19402_ (.A1(_10726_),
    .A2(_10728_),
    .B1(_00584_),
    .C1(_00585_),
    .Y(_00586_));
 sky130_fd_sc_hd__o211a_1 _19403_ (.A1(_00584_),
    .A2(_00585_),
    .B1(_10726_),
    .C1(_10728_),
    .X(_00587_));
 sky130_fd_sc_hd__nor2_1 _19404_ (.A(_00586_),
    .B(_00587_),
    .Y(_00588_));
 sky130_fd_sc_hd__xor2_2 _19405_ (.A(_00555_),
    .B(_00588_),
    .X(_00589_));
 sky130_fd_sc_hd__and2_1 _19406_ (.A(_10721_),
    .B(_10723_),
    .X(_00590_));
 sky130_fd_sc_hd__a21o_1 _19407_ (.A1(_10731_),
    .A2(_10738_),
    .B1(_10737_),
    .X(_00591_));
 sky130_fd_sc_hd__a22o_1 _19408_ (.A1(net134),
    .A2(net224),
    .B1(net220),
    .B2(net139),
    .X(_00592_));
 sky130_fd_sc_hd__and3_1 _19409_ (.A(net139),
    .B(net134),
    .C(net224),
    .X(_00593_));
 sky130_fd_sc_hd__a21bo_1 _19410_ (.A1(net220),
    .A2(_00593_),
    .B1_N(_00592_),
    .X(_00594_));
 sky130_fd_sc_hd__nand2_1 _19411_ (.A(net130),
    .B(net228),
    .Y(_00595_));
 sky130_fd_sc_hd__xor2_1 _19412_ (.A(_00594_),
    .B(_00595_),
    .X(_00596_));
 sky130_fd_sc_hd__a22o_1 _19413_ (.A1(net148),
    .A2(net211),
    .B1(net208),
    .B2(net153),
    .X(_00597_));
 sky130_fd_sc_hd__nand4_2 _19414_ (.A(net153),
    .B(net148),
    .C(net211),
    .D(net208),
    .Y(_00598_));
 sky130_fd_sc_hd__inv_2 _19415_ (.A(_00598_),
    .Y(_00599_));
 sky130_fd_sc_hd__a22oi_2 _19416_ (.A1(net143),
    .A2(net216),
    .B1(_00597_),
    .B2(_00598_),
    .Y(_00600_));
 sky130_fd_sc_hd__and4_2 _19417_ (.A(net143),
    .B(net216),
    .C(_00597_),
    .D(_00598_),
    .X(_00601_));
 sky130_fd_sc_hd__a211o_1 _19418_ (.A1(_10717_),
    .A2(_10719_),
    .B1(_00600_),
    .C1(_00601_),
    .X(_00602_));
 sky130_fd_sc_hd__o211ai_2 _19419_ (.A1(_00600_),
    .A2(_00601_),
    .B1(_10717_),
    .C1(_10719_),
    .Y(_00603_));
 sky130_fd_sc_hd__nand3_1 _19420_ (.A(_00596_),
    .B(_00602_),
    .C(_00603_),
    .Y(_00604_));
 sky130_fd_sc_hd__a21o_1 _19421_ (.A1(_00602_),
    .A2(_00603_),
    .B1(_00596_),
    .X(_00605_));
 sky130_fd_sc_hd__nand3_2 _19422_ (.A(_00591_),
    .B(_00604_),
    .C(_00605_),
    .Y(_00606_));
 sky130_fd_sc_hd__a21o_1 _19423_ (.A1(_00604_),
    .A2(_00605_),
    .B1(_00591_),
    .X(_00607_));
 sky130_fd_sc_hd__nand3b_2 _19424_ (.A_N(_00590_),
    .B(_00606_),
    .C(_00607_),
    .Y(_00608_));
 sky130_fd_sc_hd__a21bo_1 _19425_ (.A1(_00606_),
    .A2(_00607_),
    .B1_N(_00590_),
    .X(_00609_));
 sky130_fd_sc_hd__and2_2 _19426_ (.A(_00608_),
    .B(_00609_),
    .X(_00610_));
 sky130_fd_sc_hd__nand2_2 _19427_ (.A(_10734_),
    .B(_10736_),
    .Y(_00611_));
 sky130_fd_sc_hd__a32o_1 _19428_ (.A1(net173),
    .A2(net199),
    .A3(_10741_),
    .B1(_10573_),
    .B2(net195),
    .X(_00612_));
 sky130_fd_sc_hd__a22o_1 _19429_ (.A1(net164),
    .A2(net202),
    .B1(net199),
    .B2(net168),
    .X(_00613_));
 sky130_fd_sc_hd__nand4_2 _19430_ (.A(net168),
    .B(net161),
    .C(net202),
    .D(net199),
    .Y(_00614_));
 sky130_fd_sc_hd__a22o_1 _19431_ (.A1(net156),
    .A2(net206),
    .B1(_00613_),
    .B2(_00614_),
    .X(_00615_));
 sky130_fd_sc_hd__nand4_2 _19432_ (.A(net156),
    .B(net206),
    .C(_00613_),
    .D(_00614_),
    .Y(_00616_));
 sky130_fd_sc_hd__and3_1 _19433_ (.A(_00612_),
    .B(_00615_),
    .C(_00616_),
    .X(_00617_));
 sky130_fd_sc_hd__a21o_1 _19434_ (.A1(_00615_),
    .A2(_00616_),
    .B1(_00612_),
    .X(_00618_));
 sky130_fd_sc_hd__and2b_1 _19435_ (.A_N(_00617_),
    .B(_00618_),
    .X(_00619_));
 sky130_fd_sc_hd__xor2_4 _19436_ (.A(_00611_),
    .B(_00619_),
    .X(_00620_));
 sky130_fd_sc_hd__a22o_1 _19437_ (.A1(net179),
    .A2(net195),
    .B1(net193),
    .B2(net184),
    .X(_00621_));
 sky130_fd_sc_hd__nand4_1 _19438_ (.A(net184),
    .B(net179),
    .C(net196),
    .D(net194),
    .Y(_00622_));
 sky130_fd_sc_hd__and2_1 _19439_ (.A(net173),
    .B(net197),
    .X(_00623_));
 sky130_fd_sc_hd__a21o_1 _19440_ (.A1(_00621_),
    .A2(_00622_),
    .B1(_00623_),
    .X(_00624_));
 sky130_fd_sc_hd__nand3_1 _19441_ (.A(_00621_),
    .B(_00622_),
    .C(_00623_),
    .Y(_00625_));
 sky130_fd_sc_hd__o211a_1 _19442_ (.A1(_10582_),
    .A2(_10745_),
    .B1(_00624_),
    .C1(_00625_),
    .X(_00626_));
 sky130_fd_sc_hd__a211oi_1 _19443_ (.A1(_00624_),
    .A2(_00625_),
    .B1(_10582_),
    .C1(_10745_),
    .Y(_00627_));
 sky130_fd_sc_hd__nor2_2 _19444_ (.A(_00626_),
    .B(_00627_),
    .Y(_00628_));
 sky130_fd_sc_hd__and2_2 _19445_ (.A(net187),
    .B(_10579_),
    .X(_00629_));
 sky130_fd_sc_hd__a21oi_2 _19446_ (.A1(_10744_),
    .A2(_10746_),
    .B1(_00629_),
    .Y(_00630_));
 sky130_fd_sc_hd__and2b_1 _19447_ (.A_N(_00630_),
    .B(_00628_),
    .X(_00631_));
 sky130_fd_sc_hd__xnor2_4 _19448_ (.A(_00628_),
    .B(_00630_),
    .Y(_00632_));
 sky130_fd_sc_hd__xor2_4 _19449_ (.A(_00620_),
    .B(_00632_),
    .X(_00633_));
 sky130_fd_sc_hd__o21a_2 _19450_ (.A1(_10740_),
    .A2(_10750_),
    .B1(_10749_),
    .X(_00634_));
 sky130_fd_sc_hd__and2b_1 _19451_ (.A_N(_00634_),
    .B(_00633_),
    .X(_00635_));
 sky130_fd_sc_hd__xnor2_4 _19452_ (.A(_00633_),
    .B(_00634_),
    .Y(_00636_));
 sky130_fd_sc_hd__xor2_4 _19453_ (.A(_00610_),
    .B(_00636_),
    .X(_00637_));
 sky130_fd_sc_hd__a21o_1 _19454_ (.A1(_10730_),
    .A2(_10754_),
    .B1(_10753_),
    .X(_00638_));
 sky130_fd_sc_hd__nand2_1 _19455_ (.A(_00637_),
    .B(_00638_),
    .Y(_00639_));
 sky130_fd_sc_hd__xor2_4 _19456_ (.A(_00637_),
    .B(_00638_),
    .X(_00640_));
 sky130_fd_sc_hd__xnor2_2 _19457_ (.A(_00589_),
    .B(_00640_),
    .Y(_00641_));
 sky130_fd_sc_hd__a21oi_2 _19458_ (.A1(_10709_),
    .A2(_10758_),
    .B1(_10757_),
    .Y(_00642_));
 sky130_fd_sc_hd__nor2_1 _19459_ (.A(_00641_),
    .B(_00642_),
    .Y(_00643_));
 sky130_fd_sc_hd__xor2_2 _19460_ (.A(_00641_),
    .B(_00642_),
    .X(_00644_));
 sky130_fd_sc_hd__xor2_1 _19461_ (.A(_00554_),
    .B(_00644_),
    .X(_00645_));
 sky130_fd_sc_hd__a21oi_1 _19462_ (.A1(_10673_),
    .A2(_10762_),
    .B1(_10761_),
    .Y(_00646_));
 sky130_fd_sc_hd__nand2b_1 _19463_ (.A_N(_00646_),
    .B(_00645_),
    .Y(_00647_));
 sky130_fd_sc_hd__xnor2_1 _19464_ (.A(_00645_),
    .B(_00646_),
    .Y(_00648_));
 sky130_fd_sc_hd__xnor2_1 _19465_ (.A(_10781_),
    .B(_00648_),
    .Y(_00649_));
 sky130_fd_sc_hd__a21o_1 _19466_ (.A1(_10765_),
    .A2(_10767_),
    .B1(_00649_),
    .X(_00650_));
 sky130_fd_sc_hd__nand3_1 _19467_ (.A(_10765_),
    .B(_10767_),
    .C(_00649_),
    .Y(_00651_));
 sky130_fd_sc_hd__and2_1 _19468_ (.A(_00650_),
    .B(_00651_),
    .X(_00652_));
 sky130_fd_sc_hd__xnor2_2 _19469_ (.A(_10780_),
    .B(_00652_),
    .Y(_00653_));
 sky130_fd_sc_hd__a21oi_2 _19470_ (.A1(_10629_),
    .A2(_10772_),
    .B1(_10770_),
    .Y(_00654_));
 sky130_fd_sc_hd__or2_1 _19471_ (.A(_00653_),
    .B(_00654_),
    .X(_00655_));
 sky130_fd_sc_hd__xnor2_2 _19472_ (.A(_00653_),
    .B(_00654_),
    .Y(_00656_));
 sky130_fd_sc_hd__o21ai_2 _19473_ (.A1(_10617_),
    .A2(_10774_),
    .B1(_10775_),
    .Y(_00657_));
 sky130_fd_sc_hd__or3b_1 _19474_ (.A(_10619_),
    .B(_10776_),
    .C_N(_10624_),
    .X(_00658_));
 sky130_fd_sc_hd__and2_1 _19475_ (.A(_00657_),
    .B(_00658_),
    .X(_00659_));
 sky130_fd_sc_hd__xnor2_2 _19476_ (.A(_00656_),
    .B(_00659_),
    .Y(_00660_));
 sky130_fd_sc_hd__o2bb2a_1 _19477_ (.A1_N(\temp[17] ),
    .A2_N(net7),
    .B1(_06090_),
    .B2(net44),
    .X(_00661_));
 sky130_fd_sc_hd__o21ai_1 _19478_ (.A1(_03049_),
    .A2(_00660_),
    .B1(_00661_),
    .Y(_00662_));
 sky130_fd_sc_hd__mux2_1 _19479_ (.A0(net863),
    .A1(_00662_),
    .S(net4),
    .X(_00316_));
 sky130_fd_sc_hd__o21a_1 _19480_ (.A1(_00656_),
    .A2(_00659_),
    .B1(_00655_),
    .X(_00663_));
 sky130_fd_sc_hd__a21bo_1 _19481_ (.A1(_10780_),
    .A2(_00652_),
    .B1_N(_00650_),
    .X(_00664_));
 sky130_fd_sc_hd__a21o_1 _19482_ (.A1(_00525_),
    .A2(_00526_),
    .B1(_00528_),
    .X(_00665_));
 sky130_fd_sc_hd__or2_1 _19483_ (.A(_00551_),
    .B(_00553_),
    .X(_00666_));
 sky130_fd_sc_hd__o21ba_1 _19484_ (.A1(_00530_),
    .A2(_00549_),
    .B1_N(_00548_),
    .X(_00667_));
 sky130_fd_sc_hd__a21o_1 _19485_ (.A1(_00555_),
    .A2(_00588_),
    .B1(_00586_),
    .X(_00668_));
 sky130_fd_sc_hd__a22o_1 _19486_ (.A1(net286),
    .A2(net73),
    .B1(net70),
    .B2(net290),
    .X(_00669_));
 sky130_fd_sc_hd__and3_1 _19487_ (.A(net286),
    .B(net290),
    .C(net70),
    .X(_00670_));
 sky130_fd_sc_hd__a21bo_2 _19488_ (.A1(net73),
    .A2(_00670_),
    .B1_N(_00669_),
    .X(_00671_));
 sky130_fd_sc_hd__nand2_2 _19489_ (.A(net297),
    .B(net67),
    .Y(_00672_));
 sky130_fd_sc_hd__xnor2_4 _19490_ (.A(_00671_),
    .B(_00672_),
    .Y(_00673_));
 sky130_fd_sc_hd__o2bb2a_2 _19491_ (.A1_N(net73),
    .A2_N(_10785_),
    .B1(_10786_),
    .B2(_10787_),
    .X(_00674_));
 sky130_fd_sc_hd__xnor2_2 _19492_ (.A(_00673_),
    .B(_00674_),
    .Y(_00675_));
 sky130_fd_sc_hd__and4b_2 _19493_ (.A_N(net306),
    .B(net64),
    .C(net62),
    .D(net302),
    .X(_00676_));
 sky130_fd_sc_hd__inv_2 _19494_ (.A(_00676_),
    .Y(_00677_));
 sky130_fd_sc_hd__o2bb2a_1 _19495_ (.A1_N(net301),
    .A2_N(net64),
    .B1(net56),
    .B2(net306),
    .X(_00678_));
 sky130_fd_sc_hd__nor2_1 _19496_ (.A(_00676_),
    .B(_00678_),
    .Y(_00679_));
 sky130_fd_sc_hd__xnor2_1 _19497_ (.A(_00675_),
    .B(_00679_),
    .Y(_00680_));
 sky130_fd_sc_hd__o32ai_4 _19498_ (.A1(_00520_),
    .A2(_00521_),
    .A3(_00523_),
    .B1(_10789_),
    .B2(_10788_),
    .Y(_00681_));
 sky130_fd_sc_hd__xnor2_1 _19499_ (.A(_00680_),
    .B(_00681_),
    .Y(_00682_));
 sky130_fd_sc_hd__nor2_1 _19500_ (.A(_00522_),
    .B(_00682_),
    .Y(_00683_));
 sky130_fd_sc_hd__and2_1 _19501_ (.A(_00522_),
    .B(_00682_),
    .X(_00684_));
 sky130_fd_sc_hd__or2_1 _19502_ (.A(_00683_),
    .B(_00684_),
    .X(_00685_));
 sky130_fd_sc_hd__a21oi_1 _19503_ (.A1(_00560_),
    .A2(_00568_),
    .B1(_00567_),
    .Y(_00686_));
 sky130_fd_sc_hd__nand2_1 _19504_ (.A(_00535_),
    .B(_00537_),
    .Y(_00687_));
 sky130_fd_sc_hd__a32o_1 _19505_ (.A1(net271),
    .A2(net87),
    .A3(_00556_),
    .B1(_00557_),
    .B2(net96),
    .X(_00688_));
 sky130_fd_sc_hd__a22o_1 _19506_ (.A1(net269),
    .A2(net84),
    .B1(net80),
    .B2(net275),
    .X(_00689_));
 sky130_fd_sc_hd__nand4_2 _19507_ (.A(net269),
    .B(net275),
    .C(net84),
    .D(net80),
    .Y(_00690_));
 sky130_fd_sc_hd__a22o_1 _19508_ (.A1(net280),
    .A2(net77),
    .B1(_00689_),
    .B2(_00690_),
    .X(_00691_));
 sky130_fd_sc_hd__nand4_2 _19509_ (.A(net280),
    .B(net77),
    .C(_00689_),
    .D(_00690_),
    .Y(_00692_));
 sky130_fd_sc_hd__nand3_2 _19510_ (.A(_00688_),
    .B(_00691_),
    .C(_00692_),
    .Y(_00693_));
 sky130_fd_sc_hd__a21o_1 _19511_ (.A1(_00691_),
    .A2(_00692_),
    .B1(_00688_),
    .X(_00694_));
 sky130_fd_sc_hd__nand3_2 _19512_ (.A(_00687_),
    .B(_00693_),
    .C(_00694_),
    .Y(_00695_));
 sky130_fd_sc_hd__a21o_1 _19513_ (.A1(_00693_),
    .A2(_00694_),
    .B1(_00687_),
    .X(_00696_));
 sky130_fd_sc_hd__and3b_1 _19514_ (.A_N(_00686_),
    .B(_00695_),
    .C(_00696_),
    .X(_00697_));
 sky130_fd_sc_hd__a21boi_1 _19515_ (.A1(_00695_),
    .A2(_00696_),
    .B1_N(_00686_),
    .Y(_00698_));
 sky130_fd_sc_hd__a211oi_1 _19516_ (.A1(_00538_),
    .A2(_00540_),
    .B1(_00697_),
    .C1(_00698_),
    .Y(_00699_));
 sky130_fd_sc_hd__o211ai_1 _19517_ (.A1(_00697_),
    .A2(_00698_),
    .B1(_00538_),
    .C1(_00540_),
    .Y(_00700_));
 sky130_fd_sc_hd__nand2b_1 _19518_ (.A_N(_00699_),
    .B(_00700_),
    .Y(_00701_));
 sky130_fd_sc_hd__nor2_1 _19519_ (.A(_00542_),
    .B(_00544_),
    .Y(_00702_));
 sky130_fd_sc_hd__nor2_1 _19520_ (.A(_00701_),
    .B(_00702_),
    .Y(_00703_));
 sky130_fd_sc_hd__xnor2_1 _19521_ (.A(_00701_),
    .B(_00702_),
    .Y(_00704_));
 sky130_fd_sc_hd__xnor2_1 _19522_ (.A(_00685_),
    .B(_00704_),
    .Y(_00705_));
 sky130_fd_sc_hd__and2b_1 _19523_ (.A_N(_00705_),
    .B(_00668_),
    .X(_00706_));
 sky130_fd_sc_hd__xnor2_1 _19524_ (.A(_00668_),
    .B(_00705_),
    .Y(_00707_));
 sky130_fd_sc_hd__and2b_1 _19525_ (.A_N(_00667_),
    .B(_00707_),
    .X(_00708_));
 sky130_fd_sc_hd__xnor2_1 _19526_ (.A(_00667_),
    .B(_00707_),
    .Y(_00709_));
 sky130_fd_sc_hd__a31o_1 _19527_ (.A1(_00579_),
    .A2(_00580_),
    .A3(_00581_),
    .B1(_00584_),
    .X(_00710_));
 sky130_fd_sc_hd__a22o_1 _19528_ (.A1(net253),
    .A2(net95),
    .B1(net92),
    .B2(net261),
    .X(_00711_));
 sky130_fd_sc_hd__and3_1 _19529_ (.A(net253),
    .B(net259),
    .C(net92),
    .X(_00712_));
 sky130_fd_sc_hd__a21bo_1 _19530_ (.A1(net95),
    .A2(_00712_),
    .B1_N(_00711_),
    .X(_00713_));
 sky130_fd_sc_hd__nand2_1 _19531_ (.A(net266),
    .B(net87),
    .Y(_00714_));
 sky130_fd_sc_hd__xor2_1 _19532_ (.A(_00713_),
    .B(_00714_),
    .X(_00715_));
 sky130_fd_sc_hd__a22o_1 _19533_ (.A1(net243),
    .A2(net110),
    .B1(net105),
    .B2(net626),
    .X(_00716_));
 sky130_fd_sc_hd__and4_1 _19534_ (.A(net243),
    .B(net626),
    .C(net110),
    .D(net106),
    .X(_00717_));
 sky130_fd_sc_hd__nand4_2 _19535_ (.A(net243),
    .B(net627),
    .C(net111),
    .D(net105),
    .Y(_00718_));
 sky130_fd_sc_hd__a22o_1 _19536_ (.A1(net248),
    .A2(net101),
    .B1(_00716_),
    .B2(_00718_),
    .X(_00719_));
 sky130_fd_sc_hd__and4_1 _19537_ (.A(net248),
    .B(net101),
    .C(_00716_),
    .D(_00718_),
    .X(_00720_));
 sky130_fd_sc_hd__nand4_1 _19538_ (.A(net248),
    .B(net101),
    .C(_00716_),
    .D(_00718_),
    .Y(_00721_));
 sky130_fd_sc_hd__o211a_1 _19539_ (.A1(_00562_),
    .A2(_00565_),
    .B1(_00719_),
    .C1(_00721_),
    .X(_00722_));
 sky130_fd_sc_hd__a211o_1 _19540_ (.A1(_00719_),
    .A2(_00721_),
    .B1(_00562_),
    .C1(_00565_),
    .X(_00723_));
 sky130_fd_sc_hd__nand2b_1 _19541_ (.A_N(_00722_),
    .B(_00723_),
    .Y(_00724_));
 sky130_fd_sc_hd__xnor2_1 _19542_ (.A(_00715_),
    .B(_00724_),
    .Y(_00725_));
 sky130_fd_sc_hd__nand2_1 _19543_ (.A(_00574_),
    .B(_00576_),
    .Y(_00726_));
 sky130_fd_sc_hd__a32o_1 _19544_ (.A1(net130),
    .A2(net228),
    .A3(_00592_),
    .B1(_00593_),
    .B2(net220),
    .X(_00727_));
 sky130_fd_sc_hd__a22o_1 _19545_ (.A1(net120),
    .A2(net233),
    .B1(net228),
    .B2(net125),
    .X(_00728_));
 sky130_fd_sc_hd__nand4_2 _19546_ (.A(net125),
    .B(net120),
    .C(net234),
    .D(net228),
    .Y(_00729_));
 sky130_fd_sc_hd__a22o_1 _19547_ (.A1(\mul1.b[17] ),
    .A2(net239),
    .B1(_00728_),
    .B2(_00729_),
    .X(_00730_));
 sky130_fd_sc_hd__nand4_2 _19548_ (.A(\mul1.b[17] ),
    .B(net239),
    .C(_00728_),
    .D(_00729_),
    .Y(_00731_));
 sky130_fd_sc_hd__nand3_1 _19549_ (.A(_00727_),
    .B(_00730_),
    .C(_00731_),
    .Y(_00732_));
 sky130_fd_sc_hd__a21o_1 _19550_ (.A1(_00730_),
    .A2(_00731_),
    .B1(_00727_),
    .X(_00733_));
 sky130_fd_sc_hd__nand3_1 _19551_ (.A(_00726_),
    .B(_00732_),
    .C(_00733_),
    .Y(_00734_));
 sky130_fd_sc_hd__a21o_1 _19552_ (.A1(_00732_),
    .A2(_00733_),
    .B1(_00726_),
    .X(_00735_));
 sky130_fd_sc_hd__a21bo_1 _19553_ (.A1(_00571_),
    .A2(_00578_),
    .B1_N(_00577_),
    .X(_00736_));
 sky130_fd_sc_hd__nand3_1 _19554_ (.A(_00734_),
    .B(_00735_),
    .C(_00736_),
    .Y(_00737_));
 sky130_fd_sc_hd__a21o_1 _19555_ (.A1(_00734_),
    .A2(_00735_),
    .B1(_00736_),
    .X(_00738_));
 sky130_fd_sc_hd__and3_1 _19556_ (.A(_00725_),
    .B(_00737_),
    .C(_00738_),
    .X(_00739_));
 sky130_fd_sc_hd__a21oi_1 _19557_ (.A1(_00737_),
    .A2(_00738_),
    .B1(_00725_),
    .Y(_00740_));
 sky130_fd_sc_hd__a211o_1 _19558_ (.A1(_00606_),
    .A2(_00608_),
    .B1(_00739_),
    .C1(_00740_),
    .X(_00741_));
 sky130_fd_sc_hd__o211ai_2 _19559_ (.A1(_00739_),
    .A2(_00740_),
    .B1(_00606_),
    .C1(_00608_),
    .Y(_00742_));
 sky130_fd_sc_hd__and3_1 _19560_ (.A(_00710_),
    .B(_00741_),
    .C(_00742_),
    .X(_00743_));
 sky130_fd_sc_hd__a21oi_1 _19561_ (.A1(_00741_),
    .A2(_00742_),
    .B1(_00710_),
    .Y(_00744_));
 sky130_fd_sc_hd__nor2_1 _19562_ (.A(_00743_),
    .B(_00744_),
    .Y(_00745_));
 sky130_fd_sc_hd__nand2_1 _19563_ (.A(_00602_),
    .B(_00604_),
    .Y(_00746_));
 sky130_fd_sc_hd__a21o_1 _19564_ (.A1(_00611_),
    .A2(_00618_),
    .B1(_00617_),
    .X(_00747_));
 sky130_fd_sc_hd__a22o_1 _19565_ (.A1(net134),
    .A2(net220),
    .B1(net216),
    .B2(net139),
    .X(_00748_));
 sky130_fd_sc_hd__and3_1 _19566_ (.A(net139),
    .B(net134),
    .C(net220),
    .X(_00749_));
 sky130_fd_sc_hd__a21bo_1 _19567_ (.A1(net216),
    .A2(_00749_),
    .B1_N(_00748_),
    .X(_00750_));
 sky130_fd_sc_hd__nand2_1 _19568_ (.A(net130),
    .B(net224),
    .Y(_00751_));
 sky130_fd_sc_hd__xor2_1 _19569_ (.A(_00750_),
    .B(_00751_),
    .X(_00752_));
 sky130_fd_sc_hd__a22o_1 _19570_ (.A1(net148),
    .A2(net208),
    .B1(net205),
    .B2(net153),
    .X(_00753_));
 sky130_fd_sc_hd__nand4_4 _19571_ (.A(net153),
    .B(net148),
    .C(net208),
    .D(net205),
    .Y(_00754_));
 sky130_fd_sc_hd__inv_2 _19572_ (.A(_00754_),
    .Y(_00755_));
 sky130_fd_sc_hd__a22o_1 _19573_ (.A1(net143),
    .A2(net211),
    .B1(_00753_),
    .B2(_00754_),
    .X(_00756_));
 sky130_fd_sc_hd__and4_1 _19574_ (.A(net143),
    .B(net212),
    .C(_00753_),
    .D(_00754_),
    .X(_00757_));
 sky130_fd_sc_hd__nand4_2 _19575_ (.A(net143),
    .B(net212),
    .C(_00753_),
    .D(_00754_),
    .Y(_00758_));
 sky130_fd_sc_hd__o211ai_4 _19576_ (.A1(_00599_),
    .A2(_00601_),
    .B1(_00756_),
    .C1(_00758_),
    .Y(_00759_));
 sky130_fd_sc_hd__a211o_1 _19577_ (.A1(_00756_),
    .A2(_00758_),
    .B1(_00599_),
    .C1(_00601_),
    .X(_00760_));
 sky130_fd_sc_hd__nand3_2 _19578_ (.A(_00752_),
    .B(_00759_),
    .C(_00760_),
    .Y(_00761_));
 sky130_fd_sc_hd__a21o_1 _19579_ (.A1(_00759_),
    .A2(_00760_),
    .B1(_00752_),
    .X(_00762_));
 sky130_fd_sc_hd__and3_1 _19580_ (.A(_00747_),
    .B(_00761_),
    .C(_00762_),
    .X(_00763_));
 sky130_fd_sc_hd__nand3_1 _19581_ (.A(_00747_),
    .B(_00761_),
    .C(_00762_),
    .Y(_00764_));
 sky130_fd_sc_hd__a21o_1 _19582_ (.A1(_00761_),
    .A2(_00762_),
    .B1(_00747_),
    .X(_00765_));
 sky130_fd_sc_hd__and3_1 _19583_ (.A(_00746_),
    .B(_00764_),
    .C(_00765_),
    .X(_00766_));
 sky130_fd_sc_hd__a21oi_1 _19584_ (.A1(_00764_),
    .A2(_00765_),
    .B1(_00746_),
    .Y(_00767_));
 sky130_fd_sc_hd__nor2_2 _19585_ (.A(_00766_),
    .B(_00767_),
    .Y(_00768_));
 sky130_fd_sc_hd__and3_1 _19586_ (.A(net183),
    .B(net178),
    .C(net193),
    .X(_00769_));
 sky130_fd_sc_hd__nand3_2 _19587_ (.A(net183),
    .B(net178),
    .C(net194),
    .Y(_00770_));
 sky130_fd_sc_hd__o21a_2 _19588_ (.A1(net183),
    .A2(net178),
    .B1(net193),
    .X(_00771_));
 sky130_fd_sc_hd__a22o_1 _19589_ (.A1(net173),
    .A2(net195),
    .B1(_00770_),
    .B2(_00771_),
    .X(_00772_));
 sky130_fd_sc_hd__nand4_2 _19590_ (.A(net174),
    .B(net196),
    .C(_00770_),
    .D(_00771_),
    .Y(_00773_));
 sky130_fd_sc_hd__a211o_1 _19591_ (.A1(_00772_),
    .A2(_00773_),
    .B1(_10582_),
    .C1(_10745_),
    .X(_00774_));
 sky130_fd_sc_hd__o211a_1 _19592_ (.A1(_10582_),
    .A2(_10745_),
    .B1(_00772_),
    .C1(_00773_),
    .X(_00775_));
 sky130_fd_sc_hd__o211ai_2 _19593_ (.A1(_10582_),
    .A2(_10745_),
    .B1(_00772_),
    .C1(_00773_),
    .Y(_00776_));
 sky130_fd_sc_hd__a211oi_1 _19594_ (.A1(_00774_),
    .A2(_00776_),
    .B1(_00626_),
    .C1(_00629_),
    .Y(_00777_));
 sky130_fd_sc_hd__a211o_1 _19595_ (.A1(_00774_),
    .A2(_00776_),
    .B1(_00626_),
    .C1(_00629_),
    .X(_00778_));
 sky130_fd_sc_hd__o211a_1 _19596_ (.A1(_00626_),
    .A2(_00629_),
    .B1(_00774_),
    .C1(_00776_),
    .X(_00779_));
 sky130_fd_sc_hd__nor2_2 _19597_ (.A(_00777_),
    .B(_00779_),
    .Y(_00780_));
 sky130_fd_sc_hd__nand2_1 _19598_ (.A(_00614_),
    .B(_00616_),
    .Y(_00781_));
 sky130_fd_sc_hd__a21bo_1 _19599_ (.A1(_00621_),
    .A2(_00623_),
    .B1_N(_00622_),
    .X(_00782_));
 sky130_fd_sc_hd__a22o_1 _19600_ (.A1(net163),
    .A2(net200),
    .B1(net197),
    .B2(net170),
    .X(_00783_));
 sky130_fd_sc_hd__nand4_2 _19601_ (.A(net170),
    .B(net163),
    .C(net200),
    .D(net198),
    .Y(_00784_));
 sky130_fd_sc_hd__a22o_1 _19602_ (.A1(net157),
    .A2(net202),
    .B1(_00783_),
    .B2(_00784_),
    .X(_00785_));
 sky130_fd_sc_hd__nand4_2 _19603_ (.A(net158),
    .B(net203),
    .C(_00783_),
    .D(_00784_),
    .Y(_00786_));
 sky130_fd_sc_hd__nand3_1 _19604_ (.A(_00782_),
    .B(_00785_),
    .C(_00786_),
    .Y(_00787_));
 sky130_fd_sc_hd__a21o_1 _19605_ (.A1(_00785_),
    .A2(_00786_),
    .B1(_00782_),
    .X(_00788_));
 sky130_fd_sc_hd__nand3_1 _19606_ (.A(_00781_),
    .B(_00787_),
    .C(_00788_),
    .Y(_00789_));
 sky130_fd_sc_hd__a21o_1 _19607_ (.A1(_00787_),
    .A2(_00788_),
    .B1(_00781_),
    .X(_00790_));
 sky130_fd_sc_hd__and2_1 _19608_ (.A(_00789_),
    .B(_00790_),
    .X(_00791_));
 sky130_fd_sc_hd__xnor2_4 _19609_ (.A(_00780_),
    .B(_00791_),
    .Y(_00792_));
 sky130_fd_sc_hd__a21oi_4 _19610_ (.A1(_00620_),
    .A2(_00632_),
    .B1(_00631_),
    .Y(_00793_));
 sky130_fd_sc_hd__nor2_1 _19611_ (.A(_00792_),
    .B(_00793_),
    .Y(_00794_));
 sky130_fd_sc_hd__xor2_4 _19612_ (.A(_00792_),
    .B(_00793_),
    .X(_00795_));
 sky130_fd_sc_hd__xor2_4 _19613_ (.A(_00768_),
    .B(_00795_),
    .X(_00796_));
 sky130_fd_sc_hd__a21oi_2 _19614_ (.A1(_00610_),
    .A2(_00636_),
    .B1(_00635_),
    .Y(_00797_));
 sky130_fd_sc_hd__and2b_1 _19615_ (.A_N(_00797_),
    .B(_00796_),
    .X(_00798_));
 sky130_fd_sc_hd__xnor2_4 _19616_ (.A(_00796_),
    .B(_00797_),
    .Y(_00799_));
 sky130_fd_sc_hd__xnor2_2 _19617_ (.A(_00745_),
    .B(_00799_),
    .Y(_00800_));
 sky130_fd_sc_hd__a21boi_2 _19618_ (.A1(_00589_),
    .A2(_00640_),
    .B1_N(_00639_),
    .Y(_00801_));
 sky130_fd_sc_hd__nor2_1 _19619_ (.A(_00800_),
    .B(_00801_),
    .Y(_00802_));
 sky130_fd_sc_hd__xor2_2 _19620_ (.A(_00800_),
    .B(_00801_),
    .X(_00803_));
 sky130_fd_sc_hd__xor2_1 _19621_ (.A(_00709_),
    .B(_00803_),
    .X(_00804_));
 sky130_fd_sc_hd__a21oi_1 _19622_ (.A1(_00554_),
    .A2(_00644_),
    .B1(_00643_),
    .Y(_00805_));
 sky130_fd_sc_hd__nand2b_1 _19623_ (.A_N(_00805_),
    .B(_00804_),
    .Y(_00806_));
 sky130_fd_sc_hd__xnor2_1 _19624_ (.A(_00804_),
    .B(_00805_),
    .Y(_00807_));
 sky130_fd_sc_hd__nand2_1 _19625_ (.A(_00666_),
    .B(_00807_),
    .Y(_00808_));
 sky130_fd_sc_hd__xnor2_1 _19626_ (.A(_00666_),
    .B(_00807_),
    .Y(_00809_));
 sky130_fd_sc_hd__a21boi_1 _19627_ (.A1(_10781_),
    .A2(_00648_),
    .B1_N(_00647_),
    .Y(_00810_));
 sky130_fd_sc_hd__nor2_1 _19628_ (.A(_00809_),
    .B(_00810_),
    .Y(_00811_));
 sky130_fd_sc_hd__nand2_1 _19629_ (.A(_00809_),
    .B(_00810_),
    .Y(_00812_));
 sky130_fd_sc_hd__and2b_1 _19630_ (.A_N(_00811_),
    .B(_00812_),
    .X(_00813_));
 sky130_fd_sc_hd__xnor2_2 _19631_ (.A(_00665_),
    .B(_00813_),
    .Y(_00814_));
 sky130_fd_sc_hd__nand2b_1 _19632_ (.A_N(_00814_),
    .B(_00664_),
    .Y(_00815_));
 sky130_fd_sc_hd__and2b_1 _19633_ (.A_N(_00664_),
    .B(_00814_),
    .X(_00816_));
 sky130_fd_sc_hd__xnor2_2 _19634_ (.A(_00664_),
    .B(_00814_),
    .Y(_00817_));
 sky130_fd_sc_hd__xnor2_2 _19635_ (.A(_00663_),
    .B(_00817_),
    .Y(_00818_));
 sky130_fd_sc_hd__nor2_1 _19636_ (.A(net44),
    .B(_06244_),
    .Y(_00819_));
 sky130_fd_sc_hd__a221o_1 _19637_ (.A1(\temp[18] ),
    .A2(net7),
    .B1(_00818_),
    .B2(net10),
    .C1(_00819_),
    .X(_00820_));
 sky130_fd_sc_hd__mux2_1 _19638_ (.A0(net783),
    .A1(_00820_),
    .S(_03055_),
    .X(_00317_));
 sky130_fd_sc_hd__a21o_1 _19639_ (.A1(_00680_),
    .A2(_00681_),
    .B1(_00683_),
    .X(_00821_));
 sky130_fd_sc_hd__or2_1 _19640_ (.A(_00706_),
    .B(_00708_),
    .X(_00822_));
 sky130_fd_sc_hd__o21ba_1 _19641_ (.A1(_00685_),
    .A2(_00704_),
    .B1_N(_00703_),
    .X(_00823_));
 sky130_fd_sc_hd__a21bo_1 _19642_ (.A1(_00710_),
    .A2(_00742_),
    .B1_N(_00741_),
    .X(_00824_));
 sky130_fd_sc_hd__a22o_1 _19643_ (.A1(net281),
    .A2(net73),
    .B1(net70),
    .B2(net286),
    .X(_00825_));
 sky130_fd_sc_hd__nand4_1 _19644_ (.A(net281),
    .B(net285),
    .C(net73),
    .D(net70),
    .Y(_00826_));
 sky130_fd_sc_hd__nand2_1 _19645_ (.A(_00825_),
    .B(_00826_),
    .Y(_00827_));
 sky130_fd_sc_hd__nand2_1 _19646_ (.A(net291),
    .B(net67),
    .Y(_00828_));
 sky130_fd_sc_hd__xnor2_2 _19647_ (.A(_00827_),
    .B(_00828_),
    .Y(_00829_));
 sky130_fd_sc_hd__o2bb2a_2 _19648_ (.A1_N(net73),
    .A2_N(_00670_),
    .B1(_00671_),
    .B2(_00672_),
    .X(_00830_));
 sky130_fd_sc_hd__xnor2_2 _19649_ (.A(_00829_),
    .B(_00830_),
    .Y(_00831_));
 sky130_fd_sc_hd__and4b_2 _19650_ (.A_N(net301),
    .B(net64),
    .C(net62),
    .D(net297),
    .X(_00832_));
 sky130_fd_sc_hd__inv_2 _19651_ (.A(_00832_),
    .Y(_00833_));
 sky130_fd_sc_hd__o2bb2a_1 _19652_ (.A1_N(net297),
    .A2_N(net64),
    .B1(net56),
    .B2(net302),
    .X(_00834_));
 sky130_fd_sc_hd__nor2_1 _19653_ (.A(_00832_),
    .B(_00834_),
    .Y(_00835_));
 sky130_fd_sc_hd__xnor2_1 _19654_ (.A(_00831_),
    .B(_00835_),
    .Y(_00836_));
 sky130_fd_sc_hd__o32ai_4 _19655_ (.A1(_00675_),
    .A2(_00676_),
    .A3(_00678_),
    .B1(_00674_),
    .B2(_00673_),
    .Y(_00837_));
 sky130_fd_sc_hd__xnor2_1 _19656_ (.A(_00836_),
    .B(_00837_),
    .Y(_00838_));
 sky130_fd_sc_hd__nor2_1 _19657_ (.A(_00677_),
    .B(_00838_),
    .Y(_00839_));
 sky130_fd_sc_hd__and2_1 _19658_ (.A(_00677_),
    .B(_00838_),
    .X(_00840_));
 sky130_fd_sc_hd__or2_1 _19659_ (.A(_00839_),
    .B(_00840_),
    .X(_00841_));
 sky130_fd_sc_hd__a21oi_1 _19660_ (.A1(_00715_),
    .A2(_00723_),
    .B1(_00722_),
    .Y(_00842_));
 sky130_fd_sc_hd__nand2_1 _19661_ (.A(_00690_),
    .B(_00692_),
    .Y(_00843_));
 sky130_fd_sc_hd__a32o_1 _19662_ (.A1(net266),
    .A2(net87),
    .A3(_00711_),
    .B1(_00712_),
    .B2(net95),
    .X(_00844_));
 sky130_fd_sc_hd__a22o_1 _19663_ (.A1(net265),
    .A2(net84),
    .B1(net80),
    .B2(net271),
    .X(_00845_));
 sky130_fd_sc_hd__nand4_2 _19664_ (.A(net265),
    .B(net271),
    .C(net84),
    .D(net80),
    .Y(_00846_));
 sky130_fd_sc_hd__a22o_1 _19665_ (.A1(net275),
    .A2(net77),
    .B1(_00845_),
    .B2(_00846_),
    .X(_00847_));
 sky130_fd_sc_hd__nand4_2 _19666_ (.A(net275),
    .B(net77),
    .C(_00845_),
    .D(_00846_),
    .Y(_00848_));
 sky130_fd_sc_hd__nand3_2 _19667_ (.A(_00844_),
    .B(_00847_),
    .C(_00848_),
    .Y(_00849_));
 sky130_fd_sc_hd__a21o_1 _19668_ (.A1(_00847_),
    .A2(_00848_),
    .B1(_00844_),
    .X(_00850_));
 sky130_fd_sc_hd__nand3_2 _19669_ (.A(_00843_),
    .B(_00849_),
    .C(_00850_),
    .Y(_00851_));
 sky130_fd_sc_hd__a21o_1 _19670_ (.A1(_00849_),
    .A2(_00850_),
    .B1(_00843_),
    .X(_00852_));
 sky130_fd_sc_hd__and3b_1 _19671_ (.A_N(_00842_),
    .B(_00851_),
    .C(_00852_),
    .X(_00853_));
 sky130_fd_sc_hd__a21boi_1 _19672_ (.A1(_00851_),
    .A2(_00852_),
    .B1_N(_00842_),
    .Y(_00854_));
 sky130_fd_sc_hd__a211oi_2 _19673_ (.A1(_00693_),
    .A2(_00695_),
    .B1(_00853_),
    .C1(_00854_),
    .Y(_00855_));
 sky130_fd_sc_hd__o211ai_1 _19674_ (.A1(_00853_),
    .A2(_00854_),
    .B1(_00693_),
    .C1(_00695_),
    .Y(_00856_));
 sky130_fd_sc_hd__nand2b_1 _19675_ (.A_N(_00855_),
    .B(_00856_),
    .Y(_00857_));
 sky130_fd_sc_hd__nor2_1 _19676_ (.A(_00697_),
    .B(_00699_),
    .Y(_00858_));
 sky130_fd_sc_hd__nor2_1 _19677_ (.A(_00857_),
    .B(_00858_),
    .Y(_00859_));
 sky130_fd_sc_hd__xnor2_1 _19678_ (.A(_00857_),
    .B(_00858_),
    .Y(_00860_));
 sky130_fd_sc_hd__xnor2_1 _19679_ (.A(_00841_),
    .B(_00860_),
    .Y(_00861_));
 sky130_fd_sc_hd__and2b_1 _19680_ (.A_N(_00861_),
    .B(_00824_),
    .X(_00862_));
 sky130_fd_sc_hd__xnor2_1 _19681_ (.A(_00824_),
    .B(_00861_),
    .Y(_00863_));
 sky130_fd_sc_hd__and2b_1 _19682_ (.A_N(_00823_),
    .B(_00863_),
    .X(_00864_));
 sky130_fd_sc_hd__xnor2_1 _19683_ (.A(_00823_),
    .B(_00863_),
    .Y(_00865_));
 sky130_fd_sc_hd__a31o_1 _19684_ (.A1(_00734_),
    .A2(_00735_),
    .A3(_00736_),
    .B1(_00739_),
    .X(_00866_));
 sky130_fd_sc_hd__a22o_1 _19685_ (.A1(net248),
    .A2(net95),
    .B1(net92),
    .B2(net256),
    .X(_00867_));
 sky130_fd_sc_hd__and3_1 _19686_ (.A(net248),
    .B(net253),
    .C(net92),
    .X(_00868_));
 sky130_fd_sc_hd__a21bo_1 _19687_ (.A1(net96),
    .A2(_00868_),
    .B1_N(_00867_),
    .X(_00869_));
 sky130_fd_sc_hd__nand2_1 _19688_ (.A(net262),
    .B(net87),
    .Y(_00870_));
 sky130_fd_sc_hd__xor2_1 _19689_ (.A(_00869_),
    .B(_00870_),
    .X(_00871_));
 sky130_fd_sc_hd__a22o_1 _19690_ (.A1(net239),
    .A2(net111),
    .B1(net105),
    .B2(net243),
    .X(_00872_));
 sky130_fd_sc_hd__and4_1 _19691_ (.A(net245),
    .B(net239),
    .C(net110),
    .D(net106),
    .X(_00873_));
 sky130_fd_sc_hd__nand4_1 _19692_ (.A(net244),
    .B(net239),
    .C(net111),
    .D(net105),
    .Y(_00874_));
 sky130_fd_sc_hd__a22o_1 _19693_ (.A1(net626),
    .A2(net101),
    .B1(_00872_),
    .B2(_00874_),
    .X(_00875_));
 sky130_fd_sc_hd__and4_1 _19694_ (.A(net626),
    .B(net101),
    .C(_00872_),
    .D(_00874_),
    .X(_00876_));
 sky130_fd_sc_hd__nand4_1 _19695_ (.A(net626),
    .B(net101),
    .C(_00872_),
    .D(_00874_),
    .Y(_00877_));
 sky130_fd_sc_hd__o211a_1 _19696_ (.A1(_00717_),
    .A2(_00720_),
    .B1(_00875_),
    .C1(_00877_),
    .X(_00878_));
 sky130_fd_sc_hd__a211o_1 _19697_ (.A1(_00875_),
    .A2(_00877_),
    .B1(_00717_),
    .C1(_00720_),
    .X(_00879_));
 sky130_fd_sc_hd__nand2b_1 _19698_ (.A_N(_00878_),
    .B(_00879_),
    .Y(_00880_));
 sky130_fd_sc_hd__xnor2_1 _19699_ (.A(_00871_),
    .B(_00880_),
    .Y(_00881_));
 sky130_fd_sc_hd__nand2_1 _19700_ (.A(_00729_),
    .B(_00731_),
    .Y(_00882_));
 sky130_fd_sc_hd__a32o_1 _19701_ (.A1(net130),
    .A2(net224),
    .A3(_00748_),
    .B1(_00749_),
    .B2(net216),
    .X(_00883_));
 sky130_fd_sc_hd__a22o_1 _19702_ (.A1(net120),
    .A2(net229),
    .B1(net224),
    .B2(net125),
    .X(_00884_));
 sky130_fd_sc_hd__nand4_2 _19703_ (.A(net125),
    .B(net120),
    .C(net229),
    .D(net224),
    .Y(_00885_));
 sky130_fd_sc_hd__a22o_1 _19704_ (.A1(net116),
    .A2(net234),
    .B1(_00884_),
    .B2(_00885_),
    .X(_00886_));
 sky130_fd_sc_hd__nand4_2 _19705_ (.A(net116),
    .B(net234),
    .C(_00884_),
    .D(_00885_),
    .Y(_00887_));
 sky130_fd_sc_hd__nand3_1 _19706_ (.A(_00883_),
    .B(_00886_),
    .C(_00887_),
    .Y(_00888_));
 sky130_fd_sc_hd__a21o_1 _19707_ (.A1(_00886_),
    .A2(_00887_),
    .B1(_00883_),
    .X(_00889_));
 sky130_fd_sc_hd__nand3_1 _19708_ (.A(_00882_),
    .B(_00888_),
    .C(_00889_),
    .Y(_00890_));
 sky130_fd_sc_hd__a21o_1 _19709_ (.A1(_00888_),
    .A2(_00889_),
    .B1(_00882_),
    .X(_00891_));
 sky130_fd_sc_hd__a21bo_1 _19710_ (.A1(_00726_),
    .A2(_00733_),
    .B1_N(_00732_),
    .X(_00892_));
 sky130_fd_sc_hd__nand3_2 _19711_ (.A(_00890_),
    .B(_00891_),
    .C(_00892_),
    .Y(_00893_));
 sky130_fd_sc_hd__inv_2 _19712_ (.A(_00893_),
    .Y(_00894_));
 sky130_fd_sc_hd__a21o_1 _19713_ (.A1(_00890_),
    .A2(_00891_),
    .B1(_00892_),
    .X(_00895_));
 sky130_fd_sc_hd__and3_1 _19714_ (.A(_00881_),
    .B(_00893_),
    .C(_00895_),
    .X(_00896_));
 sky130_fd_sc_hd__nand3_1 _19715_ (.A(_00881_),
    .B(_00893_),
    .C(_00895_),
    .Y(_00897_));
 sky130_fd_sc_hd__a21o_1 _19716_ (.A1(_00893_),
    .A2(_00895_),
    .B1(_00881_),
    .X(_00898_));
 sky130_fd_sc_hd__o211ai_2 _19717_ (.A1(_00763_),
    .A2(_00766_),
    .B1(_00897_),
    .C1(_00898_),
    .Y(_00899_));
 sky130_fd_sc_hd__a211o_1 _19718_ (.A1(_00897_),
    .A2(_00898_),
    .B1(_00763_),
    .C1(_00766_),
    .X(_00900_));
 sky130_fd_sc_hd__and3_1 _19719_ (.A(_00866_),
    .B(_00899_),
    .C(_00900_),
    .X(_00901_));
 sky130_fd_sc_hd__a21oi_1 _19720_ (.A1(_00899_),
    .A2(_00900_),
    .B1(_00866_),
    .Y(_00902_));
 sky130_fd_sc_hd__nor2_2 _19721_ (.A(_00901_),
    .B(_00902_),
    .Y(_00903_));
 sky130_fd_sc_hd__a22o_1 _19722_ (.A1(net174),
    .A2(net193),
    .B1(_00770_),
    .B2(_00771_),
    .X(_00904_));
 sky130_fd_sc_hd__nand3_1 _19723_ (.A(net174),
    .B(_00770_),
    .C(_00771_),
    .Y(_00905_));
 sky130_fd_sc_hd__a211o_1 _19724_ (.A1(_00904_),
    .A2(_00905_),
    .B1(_10582_),
    .C1(_10745_),
    .X(_00906_));
 sky130_fd_sc_hd__o211ai_2 _19725_ (.A1(_10582_),
    .A2(_10745_),
    .B1(_00904_),
    .C1(_00905_),
    .Y(_00907_));
 sky130_fd_sc_hd__o211a_1 _19726_ (.A1(_00629_),
    .A2(_00775_),
    .B1(_00906_),
    .C1(_00907_),
    .X(_00908_));
 sky130_fd_sc_hd__o211ai_1 _19727_ (.A1(_00629_),
    .A2(_00775_),
    .B1(_00906_),
    .C1(_00907_),
    .Y(_00909_));
 sky130_fd_sc_hd__a211o_1 _19728_ (.A1(_00906_),
    .A2(_00907_),
    .B1(_00629_),
    .C1(_00775_),
    .X(_00910_));
 sky130_fd_sc_hd__nand2_1 _19729_ (.A(_00784_),
    .B(_00786_),
    .Y(_00911_));
 sky130_fd_sc_hd__a31o_1 _19730_ (.A1(net174),
    .A2(net196),
    .A3(_00771_),
    .B1(_00769_),
    .X(_00912_));
 sky130_fd_sc_hd__a22o_1 _19731_ (.A1(net163),
    .A2(net197),
    .B1(net196),
    .B2(net170),
    .X(_00913_));
 sky130_fd_sc_hd__nand4_2 _19732_ (.A(net170),
    .B(net163),
    .C(net197),
    .D(net195),
    .Y(_00914_));
 sky130_fd_sc_hd__a22o_1 _19733_ (.A1(net158),
    .A2(net199),
    .B1(_00913_),
    .B2(_00914_),
    .X(_00915_));
 sky130_fd_sc_hd__nand4_1 _19734_ (.A(net158),
    .B(net199),
    .C(_00913_),
    .D(_00914_),
    .Y(_00916_));
 sky130_fd_sc_hd__nand3_1 _19735_ (.A(_00912_),
    .B(_00915_),
    .C(_00916_),
    .Y(_00917_));
 sky130_fd_sc_hd__a21o_1 _19736_ (.A1(_00915_),
    .A2(_00916_),
    .B1(_00912_),
    .X(_00918_));
 sky130_fd_sc_hd__nand3_1 _19737_ (.A(_00911_),
    .B(_00917_),
    .C(_00918_),
    .Y(_00919_));
 sky130_fd_sc_hd__a21o_1 _19738_ (.A1(_00917_),
    .A2(_00918_),
    .B1(_00911_),
    .X(_00920_));
 sky130_fd_sc_hd__a22o_1 _19739_ (.A1(_00909_),
    .A2(_00910_),
    .B1(_00919_),
    .B2(_00920_),
    .X(_00921_));
 sky130_fd_sc_hd__nand4_1 _19740_ (.A(_00909_),
    .B(_00910_),
    .C(_00919_),
    .D(_00920_),
    .Y(_00922_));
 sky130_fd_sc_hd__a31o_1 _19741_ (.A1(_00778_),
    .A2(_00789_),
    .A3(_00790_),
    .B1(_00779_),
    .X(_00923_));
 sky130_fd_sc_hd__a21oi_1 _19742_ (.A1(_00921_),
    .A2(_00922_),
    .B1(_00923_),
    .Y(_00924_));
 sky130_fd_sc_hd__and3_1 _19743_ (.A(_00921_),
    .B(_00922_),
    .C(_00923_),
    .X(_00925_));
 sky130_fd_sc_hd__a21bo_1 _19744_ (.A1(_00781_),
    .A2(_00788_),
    .B1_N(_00787_),
    .X(_00926_));
 sky130_fd_sc_hd__a22o_1 _19745_ (.A1(net134),
    .A2(net216),
    .B1(net212),
    .B2(net139),
    .X(_00927_));
 sky130_fd_sc_hd__and3_1 _19746_ (.A(net139),
    .B(net134),
    .C(net216),
    .X(_00928_));
 sky130_fd_sc_hd__a21bo_1 _19747_ (.A1(net212),
    .A2(_00928_),
    .B1_N(_00927_),
    .X(_00929_));
 sky130_fd_sc_hd__nand2_1 _19748_ (.A(net130),
    .B(net220),
    .Y(_00930_));
 sky130_fd_sc_hd__xor2_1 _19749_ (.A(_00929_),
    .B(_00930_),
    .X(_00931_));
 sky130_fd_sc_hd__a22o_1 _19750_ (.A1(net148),
    .A2(net205),
    .B1(net203),
    .B2(net153),
    .X(_00932_));
 sky130_fd_sc_hd__nand4_4 _19751_ (.A(net153),
    .B(net148),
    .C(net206),
    .D(net203),
    .Y(_00933_));
 sky130_fd_sc_hd__a22o_1 _19752_ (.A1(\mul1.b[11] ),
    .A2(net209),
    .B1(_00932_),
    .B2(_00933_),
    .X(_00934_));
 sky130_fd_sc_hd__nand4_4 _19753_ (.A(net143),
    .B(net209),
    .C(_00932_),
    .D(_00933_),
    .Y(_00935_));
 sky130_fd_sc_hd__o211ai_4 _19754_ (.A1(_00755_),
    .A2(_00757_),
    .B1(_00934_),
    .C1(_00935_),
    .Y(_00936_));
 sky130_fd_sc_hd__a211o_1 _19755_ (.A1(_00934_),
    .A2(_00935_),
    .B1(_00755_),
    .C1(_00757_),
    .X(_00937_));
 sky130_fd_sc_hd__nand3_2 _19756_ (.A(_00931_),
    .B(_00936_),
    .C(_00937_),
    .Y(_00938_));
 sky130_fd_sc_hd__a21o_1 _19757_ (.A1(_00936_),
    .A2(_00937_),
    .B1(_00931_),
    .X(_00939_));
 sky130_fd_sc_hd__and3_1 _19758_ (.A(_00926_),
    .B(_00938_),
    .C(_00939_),
    .X(_00940_));
 sky130_fd_sc_hd__inv_2 _19759_ (.A(_00940_),
    .Y(_00941_));
 sky130_fd_sc_hd__a21oi_1 _19760_ (.A1(_00938_),
    .A2(_00939_),
    .B1(_00926_),
    .Y(_00942_));
 sky130_fd_sc_hd__a211o_2 _19761_ (.A1(_00759_),
    .A2(_00761_),
    .B1(_00940_),
    .C1(_00942_),
    .X(_00943_));
 sky130_fd_sc_hd__o211ai_1 _19762_ (.A1(_00940_),
    .A2(_00942_),
    .B1(_00759_),
    .C1(_00761_),
    .Y(_00944_));
 sky130_fd_sc_hd__and4bb_1 _19763_ (.A_N(_00924_),
    .B_N(_00925_),
    .C(_00943_),
    .D(_00944_),
    .X(_00945_));
 sky130_fd_sc_hd__a2bb2o_1 _19764_ (.A1_N(_00924_),
    .A2_N(_00925_),
    .B1(_00943_),
    .B2(_00944_),
    .X(_00946_));
 sky130_fd_sc_hd__and2b_1 _19765_ (.A_N(_00945_),
    .B(_00946_),
    .X(_00947_));
 sky130_fd_sc_hd__a21oi_2 _19766_ (.A1(_00768_),
    .A2(_00795_),
    .B1(_00794_),
    .Y(_00948_));
 sky130_fd_sc_hd__and2b_1 _19767_ (.A_N(_00948_),
    .B(_00947_),
    .X(_00949_));
 sky130_fd_sc_hd__xnor2_2 _19768_ (.A(_00947_),
    .B(_00948_),
    .Y(_00950_));
 sky130_fd_sc_hd__xnor2_2 _19769_ (.A(_00903_),
    .B(_00950_),
    .Y(_00951_));
 sky130_fd_sc_hd__a21oi_2 _19770_ (.A1(_00745_),
    .A2(_00799_),
    .B1(_00798_),
    .Y(_00952_));
 sky130_fd_sc_hd__nor2_1 _19771_ (.A(_00951_),
    .B(_00952_),
    .Y(_00953_));
 sky130_fd_sc_hd__xor2_2 _19772_ (.A(_00951_),
    .B(_00952_),
    .X(_00954_));
 sky130_fd_sc_hd__xor2_1 _19773_ (.A(_00865_),
    .B(_00954_),
    .X(_00955_));
 sky130_fd_sc_hd__a21oi_1 _19774_ (.A1(_00709_),
    .A2(_00803_),
    .B1(_00802_),
    .Y(_00956_));
 sky130_fd_sc_hd__nand2b_1 _19775_ (.A_N(_00956_),
    .B(_00955_),
    .Y(_00957_));
 sky130_fd_sc_hd__xnor2_1 _19776_ (.A(_00955_),
    .B(_00956_),
    .Y(_00958_));
 sky130_fd_sc_hd__xnor2_1 _19777_ (.A(_00822_),
    .B(_00958_),
    .Y(_00959_));
 sky130_fd_sc_hd__a21o_1 _19778_ (.A1(_00806_),
    .A2(_00808_),
    .B1(_00959_),
    .X(_00960_));
 sky130_fd_sc_hd__nand3_1 _19779_ (.A(_00806_),
    .B(_00808_),
    .C(_00959_),
    .Y(_00961_));
 sky130_fd_sc_hd__and2_1 _19780_ (.A(_00960_),
    .B(_00961_),
    .X(_00962_));
 sky130_fd_sc_hd__nand2_1 _19781_ (.A(_00821_),
    .B(_00962_),
    .Y(_00963_));
 sky130_fd_sc_hd__xnor2_1 _19782_ (.A(_00821_),
    .B(_00962_),
    .Y(_00964_));
 sky130_fd_sc_hd__a21oi_1 _19783_ (.A1(_00665_),
    .A2(_00812_),
    .B1(_00811_),
    .Y(_00965_));
 sky130_fd_sc_hd__or2_1 _19784_ (.A(_00964_),
    .B(_00965_),
    .X(_00966_));
 sky130_fd_sc_hd__nand2_1 _19785_ (.A(_00964_),
    .B(_00965_),
    .Y(_00967_));
 sky130_fd_sc_hd__and2_1 _19786_ (.A(_00966_),
    .B(_00967_),
    .X(_00968_));
 sky130_fd_sc_hd__nand2b_1 _19787_ (.A_N(_00656_),
    .B(_00817_),
    .Y(_00969_));
 sky130_fd_sc_hd__nor3_1 _19788_ (.A(_10619_),
    .B(_10776_),
    .C(_00969_),
    .Y(_00970_));
 sky130_fd_sc_hd__o221ai_4 _19789_ (.A1(_00655_),
    .A2(_00816_),
    .B1(_00969_),
    .B2(_00657_),
    .C1(_00815_),
    .Y(_00971_));
 sky130_fd_sc_hd__a21oi_4 _19790_ (.A1(_10624_),
    .A2(_00970_),
    .B1(_00971_),
    .Y(_00972_));
 sky130_fd_sc_hd__nand2b_1 _19791_ (.A_N(_00972_),
    .B(_00968_),
    .Y(_00973_));
 sky130_fd_sc_hd__xor2_2 _19792_ (.A(_00968_),
    .B(_00972_),
    .X(_00974_));
 sky130_fd_sc_hd__nor2_1 _19793_ (.A(_03049_),
    .B(_00974_),
    .Y(_00975_));
 sky130_fd_sc_hd__a221o_1 _19794_ (.A1(\temp[19] ),
    .A2(net8),
    .B1(_06402_),
    .B2(_03052_),
    .C1(_00975_),
    .X(_00976_));
 sky130_fd_sc_hd__mux2_1 _19795_ (.A0(net772),
    .A1(_00976_),
    .S(net4),
    .X(_00318_));
 sky130_fd_sc_hd__nand2_1 _19796_ (.A(_00966_),
    .B(_00973_),
    .Y(_00977_));
 sky130_fd_sc_hd__a21o_1 _19797_ (.A1(_00836_),
    .A2(_00837_),
    .B1(_00839_),
    .X(_00978_));
 sky130_fd_sc_hd__or2_1 _19798_ (.A(_00862_),
    .B(_00864_),
    .X(_00979_));
 sky130_fd_sc_hd__o21ba_1 _19799_ (.A1(_00841_),
    .A2(_00860_),
    .B1_N(_00859_),
    .X(_00980_));
 sky130_fd_sc_hd__a21bo_1 _19800_ (.A1(_00866_),
    .A2(_00900_),
    .B1_N(_00899_),
    .X(_00981_));
 sky130_fd_sc_hd__a22o_1 _19801_ (.A1(net275),
    .A2(net73),
    .B1(net70),
    .B2(net280),
    .X(_00982_));
 sky130_fd_sc_hd__nand4_2 _19802_ (.A(net275),
    .B(net280),
    .C(net73),
    .D(net70),
    .Y(_00983_));
 sky130_fd_sc_hd__a22o_1 _19803_ (.A1(net285),
    .A2(net67),
    .B1(_00982_),
    .B2(_00983_),
    .X(_00984_));
 sky130_fd_sc_hd__nand4_2 _19804_ (.A(net285),
    .B(net67),
    .C(_00982_),
    .D(_00983_),
    .Y(_00985_));
 sky130_fd_sc_hd__o21ai_1 _19805_ (.A1(_00827_),
    .A2(_00828_),
    .B1(_00826_),
    .Y(_00986_));
 sky130_fd_sc_hd__a21oi_1 _19806_ (.A1(_00984_),
    .A2(_00985_),
    .B1(_00986_),
    .Y(_00987_));
 sky130_fd_sc_hd__a21o_1 _19807_ (.A1(_00984_),
    .A2(_00985_),
    .B1(_00986_),
    .X(_00988_));
 sky130_fd_sc_hd__and3_1 _19808_ (.A(_00984_),
    .B(_00985_),
    .C(_00986_),
    .X(_00989_));
 sky130_fd_sc_hd__or2_1 _19809_ (.A(_00987_),
    .B(_00989_),
    .X(_00990_));
 sky130_fd_sc_hd__and4b_1 _19810_ (.A_N(net297),
    .B(net64),
    .C(net62),
    .D(net291),
    .X(_00991_));
 sky130_fd_sc_hd__inv_2 _19811_ (.A(_00991_),
    .Y(_00992_));
 sky130_fd_sc_hd__o2bb2a_1 _19812_ (.A1_N(net291),
    .A2_N(net64),
    .B1(_02568_),
    .B2(net297),
    .X(_00993_));
 sky130_fd_sc_hd__nor2_1 _19813_ (.A(_00991_),
    .B(_00993_),
    .Y(_00994_));
 sky130_fd_sc_hd__xnor2_2 _19814_ (.A(_00990_),
    .B(_00994_),
    .Y(_00995_));
 sky130_fd_sc_hd__o32ai_4 _19815_ (.A1(_00831_),
    .A2(_00832_),
    .A3(_00834_),
    .B1(_00830_),
    .B2(_00829_),
    .Y(_00996_));
 sky130_fd_sc_hd__xnor2_2 _19816_ (.A(_00995_),
    .B(_00996_),
    .Y(_00997_));
 sky130_fd_sc_hd__nor2_1 _19817_ (.A(_00833_),
    .B(_00997_),
    .Y(_00998_));
 sky130_fd_sc_hd__xnor2_2 _19818_ (.A(_00833_),
    .B(_00997_),
    .Y(_00999_));
 sky130_fd_sc_hd__a21o_1 _19819_ (.A1(_00871_),
    .A2(_00879_),
    .B1(_00878_),
    .X(_01000_));
 sky130_fd_sc_hd__nand2_1 _19820_ (.A(_00846_),
    .B(_00848_),
    .Y(_01001_));
 sky130_fd_sc_hd__a32o_1 _19821_ (.A1(net261),
    .A2(net87),
    .A3(_00867_),
    .B1(_00868_),
    .B2(net95),
    .X(_01002_));
 sky130_fd_sc_hd__a22o_1 _19822_ (.A1(net262),
    .A2(net84),
    .B1(net80),
    .B2(net265),
    .X(_01003_));
 sky130_fd_sc_hd__nand4_2 _19823_ (.A(net262),
    .B(net265),
    .C(net84),
    .D(net80),
    .Y(_01004_));
 sky130_fd_sc_hd__a22o_1 _19824_ (.A1(net269),
    .A2(net77),
    .B1(_01003_),
    .B2(_01004_),
    .X(_01005_));
 sky130_fd_sc_hd__nand4_2 _19825_ (.A(net269),
    .B(net77),
    .C(_01003_),
    .D(_01004_),
    .Y(_01006_));
 sky130_fd_sc_hd__nand3_2 _19826_ (.A(_01002_),
    .B(_01005_),
    .C(_01006_),
    .Y(_01007_));
 sky130_fd_sc_hd__a21o_1 _19827_ (.A1(_01005_),
    .A2(_01006_),
    .B1(_01002_),
    .X(_01008_));
 sky130_fd_sc_hd__nand3_2 _19828_ (.A(_01001_),
    .B(_01007_),
    .C(_01008_),
    .Y(_01009_));
 sky130_fd_sc_hd__a21o_1 _19829_ (.A1(_01007_),
    .A2(_01008_),
    .B1(_01001_),
    .X(_01010_));
 sky130_fd_sc_hd__and3_1 _19830_ (.A(_01000_),
    .B(_01009_),
    .C(_01010_),
    .X(_01011_));
 sky130_fd_sc_hd__a21oi_2 _19831_ (.A1(_01009_),
    .A2(_01010_),
    .B1(_01000_),
    .Y(_01012_));
 sky130_fd_sc_hd__a211oi_1 _19832_ (.A1(_00849_),
    .A2(_00851_),
    .B1(_01011_),
    .C1(_01012_),
    .Y(_01013_));
 sky130_fd_sc_hd__a211o_1 _19833_ (.A1(_00849_),
    .A2(_00851_),
    .B1(_01011_),
    .C1(_01012_),
    .X(_01014_));
 sky130_fd_sc_hd__o211ai_2 _19834_ (.A1(_01011_),
    .A2(_01012_),
    .B1(_00849_),
    .C1(_00851_),
    .Y(_01015_));
 sky130_fd_sc_hd__o211ai_2 _19835_ (.A1(_00853_),
    .A2(_00855_),
    .B1(_01014_),
    .C1(_01015_),
    .Y(_01016_));
 sky130_fd_sc_hd__a211o_1 _19836_ (.A1(_01014_),
    .A2(_01015_),
    .B1(_00853_),
    .C1(_00855_),
    .X(_01017_));
 sky130_fd_sc_hd__nand2_1 _19837_ (.A(_01016_),
    .B(_01017_),
    .Y(_01018_));
 sky130_fd_sc_hd__or2_1 _19838_ (.A(_00999_),
    .B(_01018_),
    .X(_01019_));
 sky130_fd_sc_hd__nand2_1 _19839_ (.A(_00999_),
    .B(_01018_),
    .Y(_01020_));
 sky130_fd_sc_hd__xnor2_1 _19840_ (.A(_00999_),
    .B(_01018_),
    .Y(_01021_));
 sky130_fd_sc_hd__xnor2_1 _19841_ (.A(_00981_),
    .B(_01021_),
    .Y(_01022_));
 sky130_fd_sc_hd__and2b_1 _19842_ (.A_N(_00980_),
    .B(_01022_),
    .X(_01023_));
 sky130_fd_sc_hd__xnor2_1 _19843_ (.A(_00980_),
    .B(_01022_),
    .Y(_01024_));
 sky130_fd_sc_hd__and3_2 _19844_ (.A(_00629_),
    .B(_00906_),
    .C(_00907_),
    .X(_01025_));
 sky130_fd_sc_hd__inv_2 _19845_ (.A(_01025_),
    .Y(_01026_));
 sky130_fd_sc_hd__nor2_2 _19846_ (.A(_00629_),
    .B(_00906_),
    .Y(_01027_));
 sky130_fd_sc_hd__or2_1 _19847_ (.A(_00629_),
    .B(_00906_),
    .X(_01028_));
 sky130_fd_sc_hd__nor2_2 _19848_ (.A(_01025_),
    .B(_01027_),
    .Y(_01029_));
 sky130_fd_sc_hd__nand2_1 _19849_ (.A(_00914_),
    .B(_00916_),
    .Y(_01030_));
 sky130_fd_sc_hd__a21o_2 _19850_ (.A1(net174),
    .A2(_00771_),
    .B1(_00769_),
    .X(_01031_));
 sky130_fd_sc_hd__a22o_1 _19851_ (.A1(net161),
    .A2(net195),
    .B1(net193),
    .B2(net167),
    .X(_01032_));
 sky130_fd_sc_hd__nand4_2 _19852_ (.A(net167),
    .B(net161),
    .C(net195),
    .D(net193),
    .Y(_01033_));
 sky130_fd_sc_hd__a22o_1 _19853_ (.A1(net156),
    .A2(net197),
    .B1(_01032_),
    .B2(_01033_),
    .X(_01034_));
 sky130_fd_sc_hd__nand4_1 _19854_ (.A(net158),
    .B(net197),
    .C(_01032_),
    .D(_01033_),
    .Y(_01035_));
 sky130_fd_sc_hd__nand3_1 _19855_ (.A(_01031_),
    .B(_01034_),
    .C(_01035_),
    .Y(_01036_));
 sky130_fd_sc_hd__a21o_1 _19856_ (.A1(_01034_),
    .A2(_01035_),
    .B1(_01031_),
    .X(_01037_));
 sky130_fd_sc_hd__nand3_1 _19857_ (.A(_01030_),
    .B(_01036_),
    .C(_01037_),
    .Y(_01038_));
 sky130_fd_sc_hd__a21o_1 _19858_ (.A1(_01036_),
    .A2(_01037_),
    .B1(_01030_),
    .X(_01039_));
 sky130_fd_sc_hd__a2bb2o_1 _19859_ (.A1_N(_01025_),
    .A2_N(_01027_),
    .B1(_01038_),
    .B2(_01039_),
    .X(_01040_));
 sky130_fd_sc_hd__or4bb_1 _19860_ (.A(_01025_),
    .B(_01027_),
    .C_N(_01038_),
    .D_N(_01039_),
    .X(_01041_));
 sky130_fd_sc_hd__a31o_1 _19861_ (.A1(_00910_),
    .A2(_00919_),
    .A3(_00920_),
    .B1(_00908_),
    .X(_01042_));
 sky130_fd_sc_hd__a21oi_2 _19862_ (.A1(_01040_),
    .A2(_01041_),
    .B1(_01042_),
    .Y(_01043_));
 sky130_fd_sc_hd__and3_2 _19863_ (.A(_01040_),
    .B(_01041_),
    .C(_01042_),
    .X(_01044_));
 sky130_fd_sc_hd__a21bo_1 _19864_ (.A1(_00911_),
    .A2(_00918_),
    .B1_N(_00917_),
    .X(_01045_));
 sky130_fd_sc_hd__a22o_1 _19865_ (.A1(net134),
    .A2(net213),
    .B1(net208),
    .B2(net139),
    .X(_01046_));
 sky130_fd_sc_hd__nand4_1 _19866_ (.A(net139),
    .B(net134),
    .C(net212),
    .D(net208),
    .Y(_01047_));
 sky130_fd_sc_hd__nand2_1 _19867_ (.A(_01046_),
    .B(_01047_),
    .Y(_01048_));
 sky130_fd_sc_hd__and2_1 _19868_ (.A(net130),
    .B(net216),
    .X(_01049_));
 sky130_fd_sc_hd__xnor2_1 _19869_ (.A(_01048_),
    .B(_01049_),
    .Y(_01050_));
 sky130_fd_sc_hd__a22o_1 _19870_ (.A1(net148),
    .A2(net203),
    .B1(net200),
    .B2(net153),
    .X(_01051_));
 sky130_fd_sc_hd__and4_1 _19871_ (.A(net153),
    .B(net148),
    .C(net203),
    .D(net200),
    .X(_01052_));
 sky130_fd_sc_hd__nand4_1 _19872_ (.A(net153),
    .B(net148),
    .C(net203),
    .D(net200),
    .Y(_01053_));
 sky130_fd_sc_hd__a22oi_2 _19873_ (.A1(\mul1.b[11] ),
    .A2(net205),
    .B1(_01051_),
    .B2(_01053_),
    .Y(_01054_));
 sky130_fd_sc_hd__and4_2 _19874_ (.A(net143),
    .B(net205),
    .C(_01051_),
    .D(_01053_),
    .X(_01055_));
 sky130_fd_sc_hd__a211o_1 _19875_ (.A1(_00933_),
    .A2(_00935_),
    .B1(_01054_),
    .C1(_01055_),
    .X(_01056_));
 sky130_fd_sc_hd__o211ai_2 _19876_ (.A1(_01054_),
    .A2(_01055_),
    .B1(_00933_),
    .C1(_00935_),
    .Y(_01057_));
 sky130_fd_sc_hd__nand3_2 _19877_ (.A(_01050_),
    .B(_01056_),
    .C(_01057_),
    .Y(_01058_));
 sky130_fd_sc_hd__a21o_1 _19878_ (.A1(_01056_),
    .A2(_01057_),
    .B1(_01050_),
    .X(_01059_));
 sky130_fd_sc_hd__and3_2 _19879_ (.A(_01045_),
    .B(_01058_),
    .C(_01059_),
    .X(_01060_));
 sky130_fd_sc_hd__a21oi_2 _19880_ (.A1(_01058_),
    .A2(_01059_),
    .B1(_01045_),
    .Y(_01061_));
 sky130_fd_sc_hd__a211oi_4 _19881_ (.A1(_00936_),
    .A2(_00938_),
    .B1(_01060_),
    .C1(_01061_),
    .Y(_01062_));
 sky130_fd_sc_hd__o211a_1 _19882_ (.A1(_01060_),
    .A2(_01061_),
    .B1(_00936_),
    .C1(_00938_),
    .X(_01063_));
 sky130_fd_sc_hd__o22ai_1 _19883_ (.A1(_01043_),
    .A2(_01044_),
    .B1(_01062_),
    .B2(_01063_),
    .Y(_01064_));
 sky130_fd_sc_hd__nor4_1 _19884_ (.A(_01043_),
    .B(_01044_),
    .C(_01062_),
    .D(_01063_),
    .Y(_01065_));
 sky130_fd_sc_hd__or4_1 _19885_ (.A(_01043_),
    .B(_01044_),
    .C(_01062_),
    .D(_01063_),
    .X(_01066_));
 sky130_fd_sc_hd__o211a_1 _19886_ (.A1(_00925_),
    .A2(_00945_),
    .B1(_01064_),
    .C1(_01066_),
    .X(_01067_));
 sky130_fd_sc_hd__inv_2 _19887_ (.A(_01067_),
    .Y(_01068_));
 sky130_fd_sc_hd__a211oi_1 _19888_ (.A1(_01064_),
    .A2(_01066_),
    .B1(_00925_),
    .C1(_00945_),
    .Y(_01069_));
 sky130_fd_sc_hd__a22o_1 _19889_ (.A1(net628),
    .A2(net95),
    .B1(net92),
    .B2(net250),
    .X(_01070_));
 sky130_fd_sc_hd__nand4_1 _19890_ (.A(net628),
    .B(net250),
    .C(net95),
    .D(net92),
    .Y(_01071_));
 sky130_fd_sc_hd__nand2_1 _19891_ (.A(_01070_),
    .B(_01071_),
    .Y(_01072_));
 sky130_fd_sc_hd__and2_1 _19892_ (.A(net256),
    .B(net87),
    .X(_01073_));
 sky130_fd_sc_hd__xnor2_1 _19893_ (.A(_01072_),
    .B(_01073_),
    .Y(_01074_));
 sky130_fd_sc_hd__a22o_1 _19894_ (.A1(net110),
    .A2(net233),
    .B1(net105),
    .B2(net241),
    .X(_01075_));
 sky130_fd_sc_hd__nand4_1 _19895_ (.A(net241),
    .B(net110),
    .C(net236),
    .D(net105),
    .Y(_01076_));
 sky130_fd_sc_hd__and2_1 _19896_ (.A(net245),
    .B(net101),
    .X(_01077_));
 sky130_fd_sc_hd__a21o_1 _19897_ (.A1(_01075_),
    .A2(_01076_),
    .B1(_01077_),
    .X(_01078_));
 sky130_fd_sc_hd__nand3_1 _19898_ (.A(_01075_),
    .B(_01076_),
    .C(_01077_),
    .Y(_01079_));
 sky130_fd_sc_hd__o211a_1 _19899_ (.A1(_00873_),
    .A2(_00876_),
    .B1(_01078_),
    .C1(_01079_),
    .X(_01080_));
 sky130_fd_sc_hd__a211o_1 _19900_ (.A1(_01078_),
    .A2(_01079_),
    .B1(_00873_),
    .C1(_00876_),
    .X(_01081_));
 sky130_fd_sc_hd__nand2b_1 _19901_ (.A_N(_01080_),
    .B(_01081_),
    .Y(_01082_));
 sky130_fd_sc_hd__xnor2_1 _19902_ (.A(_01074_),
    .B(_01082_),
    .Y(_01083_));
 sky130_fd_sc_hd__nand2_1 _19903_ (.A(_00885_),
    .B(_00887_),
    .Y(_01084_));
 sky130_fd_sc_hd__a32o_1 _19904_ (.A1(net130),
    .A2(net220),
    .A3(_00927_),
    .B1(_00928_),
    .B2(net212),
    .X(_01085_));
 sky130_fd_sc_hd__a22o_1 _19905_ (.A1(net120),
    .A2(net224),
    .B1(net220),
    .B2(net125),
    .X(_01086_));
 sky130_fd_sc_hd__nand4_2 _19906_ (.A(net125),
    .B(net120),
    .C(net224),
    .D(net220),
    .Y(_01087_));
 sky130_fd_sc_hd__a22o_1 _19907_ (.A1(net116),
    .A2(net231),
    .B1(_01086_),
    .B2(_01087_),
    .X(_01088_));
 sky130_fd_sc_hd__nand4_2 _19908_ (.A(net116),
    .B(net231),
    .C(_01086_),
    .D(_01087_),
    .Y(_01089_));
 sky130_fd_sc_hd__nand3_1 _19909_ (.A(_01085_),
    .B(_01088_),
    .C(_01089_),
    .Y(_01090_));
 sky130_fd_sc_hd__a21o_1 _19910_ (.A1(_01088_),
    .A2(_01089_),
    .B1(_01085_),
    .X(_01091_));
 sky130_fd_sc_hd__nand3_1 _19911_ (.A(_01084_),
    .B(_01090_),
    .C(_01091_),
    .Y(_01092_));
 sky130_fd_sc_hd__a21o_1 _19912_ (.A1(_01090_),
    .A2(_01091_),
    .B1(_01084_),
    .X(_01093_));
 sky130_fd_sc_hd__a21bo_1 _19913_ (.A1(_00882_),
    .A2(_00889_),
    .B1_N(_00888_),
    .X(_01094_));
 sky130_fd_sc_hd__nand3_2 _19914_ (.A(_01092_),
    .B(_01093_),
    .C(_01094_),
    .Y(_01095_));
 sky130_fd_sc_hd__inv_2 _19915_ (.A(_01095_),
    .Y(_01096_));
 sky130_fd_sc_hd__a21o_1 _19916_ (.A1(_01092_),
    .A2(_01093_),
    .B1(_01094_),
    .X(_01097_));
 sky130_fd_sc_hd__and3_2 _19917_ (.A(_01083_),
    .B(_01095_),
    .C(_01097_),
    .X(_01098_));
 sky130_fd_sc_hd__a21oi_2 _19918_ (.A1(_01095_),
    .A2(_01097_),
    .B1(_01083_),
    .Y(_01099_));
 sky130_fd_sc_hd__a211o_2 _19919_ (.A1(_00941_),
    .A2(_00943_),
    .B1(_01098_),
    .C1(_01099_),
    .X(_01100_));
 sky130_fd_sc_hd__o211ai_4 _19920_ (.A1(_01098_),
    .A2(_01099_),
    .B1(_00941_),
    .C1(_00943_),
    .Y(_01101_));
 sky130_fd_sc_hd__o211ai_4 _19921_ (.A1(_00894_),
    .A2(_00896_),
    .B1(_01100_),
    .C1(_01101_),
    .Y(_01102_));
 sky130_fd_sc_hd__a211o_1 _19922_ (.A1(_01100_),
    .A2(_01101_),
    .B1(_00894_),
    .C1(_00896_),
    .X(_01103_));
 sky130_fd_sc_hd__or4bb_1 _19923_ (.A(_01067_),
    .B(_01069_),
    .C_N(_01102_),
    .D_N(_01103_),
    .X(_01104_));
 sky130_fd_sc_hd__a2bb2o_1 _19924_ (.A1_N(_01067_),
    .A2_N(_01069_),
    .B1(_01102_),
    .B2(_01103_),
    .X(_01105_));
 sky130_fd_sc_hd__and2_1 _19925_ (.A(_01104_),
    .B(_01105_),
    .X(_01106_));
 sky130_fd_sc_hd__a21oi_2 _19926_ (.A1(_00903_),
    .A2(_00950_),
    .B1(_00949_),
    .Y(_01107_));
 sky130_fd_sc_hd__and2b_1 _19927_ (.A_N(_01107_),
    .B(_01106_),
    .X(_01108_));
 sky130_fd_sc_hd__xnor2_2 _19928_ (.A(_01106_),
    .B(_01107_),
    .Y(_01109_));
 sky130_fd_sc_hd__xor2_1 _19929_ (.A(_01024_),
    .B(_01109_),
    .X(_01110_));
 sky130_fd_sc_hd__a21oi_1 _19930_ (.A1(_00865_),
    .A2(_00954_),
    .B1(_00953_),
    .Y(_01111_));
 sky130_fd_sc_hd__nand2b_1 _19931_ (.A_N(_01111_),
    .B(_01110_),
    .Y(_01112_));
 sky130_fd_sc_hd__xnor2_1 _19932_ (.A(_01110_),
    .B(_01111_),
    .Y(_01113_));
 sky130_fd_sc_hd__nand2_1 _19933_ (.A(_00979_),
    .B(_01113_),
    .Y(_01114_));
 sky130_fd_sc_hd__xnor2_1 _19934_ (.A(_00979_),
    .B(_01113_),
    .Y(_01115_));
 sky130_fd_sc_hd__a21boi_1 _19935_ (.A1(_00822_),
    .A2(_00958_),
    .B1_N(_00957_),
    .Y(_01116_));
 sky130_fd_sc_hd__nor2_1 _19936_ (.A(_01115_),
    .B(_01116_),
    .Y(_01117_));
 sky130_fd_sc_hd__nand2_1 _19937_ (.A(_01115_),
    .B(_01116_),
    .Y(_01118_));
 sky130_fd_sc_hd__and2b_1 _19938_ (.A_N(_01117_),
    .B(_01118_),
    .X(_01119_));
 sky130_fd_sc_hd__xnor2_1 _19939_ (.A(_00978_),
    .B(_01119_),
    .Y(_01120_));
 sky130_fd_sc_hd__a21o_1 _19940_ (.A1(_00960_),
    .A2(_00963_),
    .B1(_01120_),
    .X(_01121_));
 sky130_fd_sc_hd__inv_2 _19941_ (.A(_01121_),
    .Y(_01122_));
 sky130_fd_sc_hd__and3_1 _19942_ (.A(_00960_),
    .B(_00963_),
    .C(_01120_),
    .X(_01123_));
 sky130_fd_sc_hd__nor2_1 _19943_ (.A(_01122_),
    .B(_01123_),
    .Y(_01124_));
 sky130_fd_sc_hd__xnor2_2 _19944_ (.A(_00977_),
    .B(_01124_),
    .Y(_01125_));
 sky130_fd_sc_hd__nand2_1 _19945_ (.A(net733),
    .B(net8),
    .Y(_01126_));
 sky130_fd_sc_hd__o221ai_1 _19946_ (.A1(net44),
    .A2(_06552_),
    .B1(_01125_),
    .B2(_03049_),
    .C1(_01126_),
    .Y(_01127_));
 sky130_fd_sc_hd__mux2_1 _19947_ (.A0(net735),
    .A1(_01127_),
    .S(net4),
    .X(_00319_));
 sky130_fd_sc_hd__a21o_1 _19948_ (.A1(_00995_),
    .A2(_00996_),
    .B1(_00998_),
    .X(_01128_));
 sky130_fd_sc_hd__a31o_1 _19949_ (.A1(_00981_),
    .A2(_01019_),
    .A3(_01020_),
    .B1(_01023_),
    .X(_01129_));
 sky130_fd_sc_hd__nand2_1 _19950_ (.A(_01033_),
    .B(_01035_),
    .Y(_01130_));
 sky130_fd_sc_hd__nand3_2 _19951_ (.A(net167),
    .B(net161),
    .C(net193),
    .Y(_01131_));
 sky130_fd_sc_hd__o21a_1 _19952_ (.A1(net167),
    .A2(net161),
    .B1(net193),
    .X(_01132_));
 sky130_fd_sc_hd__nand2_1 _19953_ (.A(_01131_),
    .B(_01132_),
    .Y(_01133_));
 sky130_fd_sc_hd__a22o_1 _19954_ (.A1(net158),
    .A2(net195),
    .B1(_01131_),
    .B2(_01132_),
    .X(_01134_));
 sky130_fd_sc_hd__nand4_2 _19955_ (.A(net158),
    .B(net195),
    .C(_01131_),
    .D(_01132_),
    .Y(_01135_));
 sky130_fd_sc_hd__nand3_1 _19956_ (.A(_01031_),
    .B(_01134_),
    .C(_01135_),
    .Y(_01136_));
 sky130_fd_sc_hd__a21o_1 _19957_ (.A1(_01134_),
    .A2(_01135_),
    .B1(_01031_),
    .X(_01137_));
 sky130_fd_sc_hd__and3_1 _19958_ (.A(_01130_),
    .B(_01136_),
    .C(_01137_),
    .X(_01138_));
 sky130_fd_sc_hd__a21oi_1 _19959_ (.A1(_01136_),
    .A2(_01137_),
    .B1(_01130_),
    .Y(_01139_));
 sky130_fd_sc_hd__o22ai_1 _19960_ (.A1(_01025_),
    .A2(_01027_),
    .B1(_01138_),
    .B2(_01139_),
    .Y(_01140_));
 sky130_fd_sc_hd__or4_1 _19961_ (.A(_01025_),
    .B(_01027_),
    .C(_01138_),
    .D(_01139_),
    .X(_01141_));
 sky130_fd_sc_hd__a31o_1 _19962_ (.A1(_01028_),
    .A2(_01038_),
    .A3(_01039_),
    .B1(_01025_),
    .X(_01142_));
 sky130_fd_sc_hd__and3_1 _19963_ (.A(_01140_),
    .B(_01141_),
    .C(_01142_),
    .X(_01143_));
 sky130_fd_sc_hd__a21oi_1 _19964_ (.A1(_01140_),
    .A2(_01141_),
    .B1(_01142_),
    .Y(_01144_));
 sky130_fd_sc_hd__a21bo_1 _19965_ (.A1(_01030_),
    .A2(_01037_),
    .B1_N(_01036_),
    .X(_01145_));
 sky130_fd_sc_hd__a22o_1 _19966_ (.A1(net134),
    .A2(net208),
    .B1(net205),
    .B2(net139),
    .X(_01146_));
 sky130_fd_sc_hd__and3_1 _19967_ (.A(net139),
    .B(net134),
    .C(net210),
    .X(_01147_));
 sky130_fd_sc_hd__a21bo_1 _19968_ (.A1(net205),
    .A2(_01147_),
    .B1_N(_01146_),
    .X(_01148_));
 sky130_fd_sc_hd__nand2_1 _19969_ (.A(net130),
    .B(net213),
    .Y(_01149_));
 sky130_fd_sc_hd__xor2_1 _19970_ (.A(_01148_),
    .B(_01149_),
    .X(_01150_));
 sky130_fd_sc_hd__a22o_1 _19971_ (.A1(net148),
    .A2(net200),
    .B1(net198),
    .B2(net153),
    .X(_01151_));
 sky130_fd_sc_hd__nand4_2 _19972_ (.A(net153),
    .B(net148),
    .C(net200),
    .D(net198),
    .Y(_01152_));
 sky130_fd_sc_hd__a22o_1 _19973_ (.A1(net143),
    .A2(net202),
    .B1(_01151_),
    .B2(_01152_),
    .X(_01153_));
 sky130_fd_sc_hd__nand4_2 _19974_ (.A(net143),
    .B(net202),
    .C(_01151_),
    .D(_01152_),
    .Y(_01154_));
 sky130_fd_sc_hd__o211ai_2 _19975_ (.A1(_01052_),
    .A2(_01055_),
    .B1(_01153_),
    .C1(_01154_),
    .Y(_01155_));
 sky130_fd_sc_hd__a211o_1 _19976_ (.A1(_01153_),
    .A2(_01154_),
    .B1(_01052_),
    .C1(_01055_),
    .X(_01156_));
 sky130_fd_sc_hd__nand3_1 _19977_ (.A(_01150_),
    .B(_01155_),
    .C(_01156_),
    .Y(_01157_));
 sky130_fd_sc_hd__a21o_1 _19978_ (.A1(_01155_),
    .A2(_01156_),
    .B1(_01150_),
    .X(_01158_));
 sky130_fd_sc_hd__and3_1 _19979_ (.A(_01145_),
    .B(_01157_),
    .C(_01158_),
    .X(_01159_));
 sky130_fd_sc_hd__a21oi_1 _19980_ (.A1(_01157_),
    .A2(_01158_),
    .B1(_01145_),
    .Y(_01160_));
 sky130_fd_sc_hd__a211oi_1 _19981_ (.A1(_01056_),
    .A2(_01058_),
    .B1(_01159_),
    .C1(_01160_),
    .Y(_01161_));
 sky130_fd_sc_hd__o211a_1 _19982_ (.A1(_01159_),
    .A2(_01160_),
    .B1(_01056_),
    .C1(_01058_),
    .X(_01162_));
 sky130_fd_sc_hd__o22ai_1 _19983_ (.A1(_01143_),
    .A2(_01144_),
    .B1(_01161_),
    .B2(_01162_),
    .Y(_01163_));
 sky130_fd_sc_hd__or4_1 _19984_ (.A(_01143_),
    .B(_01144_),
    .C(_01161_),
    .D(_01162_),
    .X(_01164_));
 sky130_fd_sc_hd__a211oi_1 _19985_ (.A1(_01163_),
    .A2(_01164_),
    .B1(_01044_),
    .C1(_01065_),
    .Y(_01165_));
 sky130_fd_sc_hd__o211a_1 _19986_ (.A1(_01044_),
    .A2(_01065_),
    .B1(_01163_),
    .C1(_01164_),
    .X(_01166_));
 sky130_fd_sc_hd__a22o_1 _19987_ (.A1(net245),
    .A2(net96),
    .B1(net92),
    .B2(net628),
    .X(_01167_));
 sky130_fd_sc_hd__and3_1 _19988_ (.A(net245),
    .B(net628),
    .C(net92),
    .X(_01168_));
 sky130_fd_sc_hd__a21bo_1 _19989_ (.A1(net96),
    .A2(_01168_),
    .B1_N(_01167_),
    .X(_01169_));
 sky130_fd_sc_hd__nand2_1 _19990_ (.A(net250),
    .B(net87),
    .Y(_01170_));
 sky130_fd_sc_hd__xnor2_1 _19991_ (.A(_01169_),
    .B(_01170_),
    .Y(_01171_));
 sky130_fd_sc_hd__a22o_1 _19992_ (.A1(net236),
    .A2(net105),
    .B1(net230),
    .B2(net110),
    .X(_01172_));
 sky130_fd_sc_hd__nand4_2 _19993_ (.A(net110),
    .B(net236),
    .C(net105),
    .D(net231),
    .Y(_01173_));
 sky130_fd_sc_hd__a22o_1 _19994_ (.A1(net241),
    .A2(net101),
    .B1(_01172_),
    .B2(_01173_),
    .X(_01174_));
 sky130_fd_sc_hd__nand4_2 _19995_ (.A(net241),
    .B(net101),
    .C(_01172_),
    .D(_01173_),
    .Y(_01175_));
 sky130_fd_sc_hd__a21bo_1 _19996_ (.A1(_01075_),
    .A2(_01077_),
    .B1_N(_01076_),
    .X(_01176_));
 sky130_fd_sc_hd__nand3_1 _19997_ (.A(_01174_),
    .B(_01175_),
    .C(_01176_),
    .Y(_01177_));
 sky130_fd_sc_hd__a21o_1 _19998_ (.A1(_01174_),
    .A2(_01175_),
    .B1(_01176_),
    .X(_01178_));
 sky130_fd_sc_hd__nand2_1 _19999_ (.A(_01177_),
    .B(_01178_),
    .Y(_01179_));
 sky130_fd_sc_hd__xor2_1 _20000_ (.A(_01171_),
    .B(_01179_),
    .X(_01180_));
 sky130_fd_sc_hd__nand2_1 _20001_ (.A(_01087_),
    .B(_01089_),
    .Y(_01181_));
 sky130_fd_sc_hd__a21boi_1 _20002_ (.A1(_01046_),
    .A2(_01049_),
    .B1_N(_01047_),
    .Y(_01182_));
 sky130_fd_sc_hd__a22oi_1 _20003_ (.A1(net121),
    .A2(net222),
    .B1(net216),
    .B2(net126),
    .Y(_01183_));
 sky130_fd_sc_hd__and4_1 _20004_ (.A(net126),
    .B(net121),
    .C(net222),
    .D(net217),
    .X(_01184_));
 sky130_fd_sc_hd__o2bb2a_1 _20005_ (.A1_N(net116),
    .A2_N(net226),
    .B1(_01183_),
    .B2(_01184_),
    .X(_01185_));
 sky130_fd_sc_hd__and4bb_1 _20006_ (.A_N(_01183_),
    .B_N(_01184_),
    .C(net116),
    .D(net226),
    .X(_01186_));
 sky130_fd_sc_hd__or3_1 _20007_ (.A(_01182_),
    .B(_01185_),
    .C(_01186_),
    .X(_01187_));
 sky130_fd_sc_hd__o21ai_1 _20008_ (.A1(_01185_),
    .A2(_01186_),
    .B1(_01182_),
    .Y(_01188_));
 sky130_fd_sc_hd__nand3_1 _20009_ (.A(_01181_),
    .B(_01187_),
    .C(_01188_),
    .Y(_01189_));
 sky130_fd_sc_hd__a21o_1 _20010_ (.A1(_01187_),
    .A2(_01188_),
    .B1(_01181_),
    .X(_01190_));
 sky130_fd_sc_hd__a21bo_1 _20011_ (.A1(_01084_),
    .A2(_01091_),
    .B1_N(_01090_),
    .X(_01191_));
 sky130_fd_sc_hd__nand3_1 _20012_ (.A(_01189_),
    .B(_01190_),
    .C(_01191_),
    .Y(_01192_));
 sky130_fd_sc_hd__a21o_1 _20013_ (.A1(_01189_),
    .A2(_01190_),
    .B1(_01191_),
    .X(_01193_));
 sky130_fd_sc_hd__nand3_1 _20014_ (.A(_01180_),
    .B(_01192_),
    .C(_01193_),
    .Y(_01194_));
 sky130_fd_sc_hd__a21o_1 _20015_ (.A1(_01192_),
    .A2(_01193_),
    .B1(_01180_),
    .X(_01195_));
 sky130_fd_sc_hd__o211ai_2 _20016_ (.A1(_01060_),
    .A2(_01062_),
    .B1(_01194_),
    .C1(_01195_),
    .Y(_01196_));
 sky130_fd_sc_hd__a211o_1 _20017_ (.A1(_01194_),
    .A2(_01195_),
    .B1(_01060_),
    .C1(_01062_),
    .X(_01197_));
 sky130_fd_sc_hd__o211ai_2 _20018_ (.A1(_01096_),
    .A2(_01098_),
    .B1(_01196_),
    .C1(_01197_),
    .Y(_01198_));
 sky130_fd_sc_hd__a211o_1 _20019_ (.A1(_01196_),
    .A2(_01197_),
    .B1(_01096_),
    .C1(_01098_),
    .X(_01199_));
 sky130_fd_sc_hd__and4bb_1 _20020_ (.A_N(_01165_),
    .B_N(_01166_),
    .C(_01198_),
    .D(_01199_),
    .X(_01200_));
 sky130_fd_sc_hd__a2bb2oi_1 _20021_ (.A1_N(_01165_),
    .A2_N(_01166_),
    .B1(_01198_),
    .B2(_01199_),
    .Y(_01201_));
 sky130_fd_sc_hd__a211o_1 _20022_ (.A1(_01068_),
    .A2(_01104_),
    .B1(_01200_),
    .C1(_01201_),
    .X(_01202_));
 sky130_fd_sc_hd__o211ai_1 _20023_ (.A1(_01200_),
    .A2(_01201_),
    .B1(_01068_),
    .C1(_01104_),
    .Y(_01203_));
 sky130_fd_sc_hd__nand2_1 _20024_ (.A(_01202_),
    .B(_01203_),
    .Y(_01204_));
 sky130_fd_sc_hd__a22oi_1 _20025_ (.A1(net269),
    .A2(net73),
    .B1(net70),
    .B2(net275),
    .Y(_01205_));
 sky130_fd_sc_hd__and4_1 _20026_ (.A(net269),
    .B(net275),
    .C(net73),
    .D(net70),
    .X(_01206_));
 sky130_fd_sc_hd__o2bb2a_1 _20027_ (.A1_N(net280),
    .A2_N(net67),
    .B1(_01205_),
    .B2(_01206_),
    .X(_01207_));
 sky130_fd_sc_hd__and4bb_1 _20028_ (.A_N(_01205_),
    .B_N(_01206_),
    .C(net280),
    .D(net67),
    .X(_01208_));
 sky130_fd_sc_hd__o211a_1 _20029_ (.A1(_01207_),
    .A2(_01208_),
    .B1(_00983_),
    .C1(_00985_),
    .X(_01209_));
 sky130_fd_sc_hd__a211o_1 _20030_ (.A1(_00983_),
    .A2(_00985_),
    .B1(_01207_),
    .C1(_01208_),
    .X(_01210_));
 sky130_fd_sc_hd__nand2b_1 _20031_ (.A_N(_01209_),
    .B(_01210_),
    .Y(_01211_));
 sky130_fd_sc_hd__and4b_1 _20032_ (.A_N(net291),
    .B(net64),
    .C(net62),
    .D(net285),
    .X(_01212_));
 sky130_fd_sc_hd__inv_2 _20033_ (.A(_01212_),
    .Y(_01213_));
 sky130_fd_sc_hd__o2bb2a_1 _20034_ (.A1_N(net285),
    .A2_N(net64),
    .B1(net56),
    .B2(net290),
    .X(_01214_));
 sky130_fd_sc_hd__nor2_1 _20035_ (.A(_01212_),
    .B(_01214_),
    .Y(_01215_));
 sky130_fd_sc_hd__xnor2_1 _20036_ (.A(_01211_),
    .B(_01215_),
    .Y(_01216_));
 sky130_fd_sc_hd__a21o_1 _20037_ (.A1(_00988_),
    .A2(_00994_),
    .B1(_00989_),
    .X(_01217_));
 sky130_fd_sc_hd__and2_1 _20038_ (.A(_01216_),
    .B(_01217_),
    .X(_01218_));
 sky130_fd_sc_hd__xnor2_1 _20039_ (.A(_01216_),
    .B(_01217_),
    .Y(_01219_));
 sky130_fd_sc_hd__nor2_1 _20040_ (.A(_00992_),
    .B(_01219_),
    .Y(_01220_));
 sky130_fd_sc_hd__xnor2_1 _20041_ (.A(_00992_),
    .B(_01219_),
    .Y(_01221_));
 sky130_fd_sc_hd__a21o_1 _20042_ (.A1(_01074_),
    .A2(_01081_),
    .B1(_01080_),
    .X(_01222_));
 sky130_fd_sc_hd__nand2_1 _20043_ (.A(_01004_),
    .B(_01006_),
    .Y(_01223_));
 sky130_fd_sc_hd__a21boi_1 _20044_ (.A1(_01070_),
    .A2(_01073_),
    .B1_N(_01071_),
    .Y(_01224_));
 sky130_fd_sc_hd__a22oi_1 _20045_ (.A1(net255),
    .A2(net84),
    .B1(net80),
    .B2(net261),
    .Y(_01225_));
 sky130_fd_sc_hd__and4_1 _20046_ (.A(net255),
    .B(net261),
    .C(net84),
    .D(net80),
    .X(_01226_));
 sky130_fd_sc_hd__o2bb2a_1 _20047_ (.A1_N(net265),
    .A2_N(net77),
    .B1(_01225_),
    .B2(_01226_),
    .X(_01227_));
 sky130_fd_sc_hd__and4bb_1 _20048_ (.A_N(_01225_),
    .B_N(_01226_),
    .C(net265),
    .D(net77),
    .X(_01228_));
 sky130_fd_sc_hd__or3_1 _20049_ (.A(_01224_),
    .B(_01227_),
    .C(_01228_),
    .X(_01229_));
 sky130_fd_sc_hd__o21ai_1 _20050_ (.A1(_01227_),
    .A2(_01228_),
    .B1(_01224_),
    .Y(_01230_));
 sky130_fd_sc_hd__nand3_1 _20051_ (.A(_01223_),
    .B(_01229_),
    .C(_01230_),
    .Y(_01231_));
 sky130_fd_sc_hd__a21o_1 _20052_ (.A1(_01229_),
    .A2(_01230_),
    .B1(_01223_),
    .X(_01232_));
 sky130_fd_sc_hd__and3_1 _20053_ (.A(_01222_),
    .B(_01231_),
    .C(_01232_),
    .X(_01233_));
 sky130_fd_sc_hd__a21oi_1 _20054_ (.A1(_01231_),
    .A2(_01232_),
    .B1(_01222_),
    .Y(_01234_));
 sky130_fd_sc_hd__a211o_1 _20055_ (.A1(_01007_),
    .A2(_01009_),
    .B1(_01233_),
    .C1(_01234_),
    .X(_01235_));
 sky130_fd_sc_hd__o211ai_2 _20056_ (.A1(_01233_),
    .A2(_01234_),
    .B1(_01007_),
    .C1(_01009_),
    .Y(_01236_));
 sky130_fd_sc_hd__o211a_1 _20057_ (.A1(_01011_),
    .A2(_01013_),
    .B1(_01235_),
    .C1(_01236_),
    .X(_01237_));
 sky130_fd_sc_hd__a211oi_1 _20058_ (.A1(_01235_),
    .A2(_01236_),
    .B1(_01011_),
    .C1(_01013_),
    .Y(_01238_));
 sky130_fd_sc_hd__nor3_1 _20059_ (.A(_01221_),
    .B(_01237_),
    .C(_01238_),
    .Y(_01239_));
 sky130_fd_sc_hd__o21a_1 _20060_ (.A1(_01237_),
    .A2(_01238_),
    .B1(_01221_),
    .X(_01240_));
 sky130_fd_sc_hd__a211oi_2 _20061_ (.A1(_01100_),
    .A2(_01102_),
    .B1(_01239_),
    .C1(_01240_),
    .Y(_01241_));
 sky130_fd_sc_hd__o211a_1 _20062_ (.A1(_01239_),
    .A2(_01240_),
    .B1(_01100_),
    .C1(_01102_),
    .X(_01242_));
 sky130_fd_sc_hd__a211oi_1 _20063_ (.A1(_01016_),
    .A2(_01019_),
    .B1(_01241_),
    .C1(_01242_),
    .Y(_01243_));
 sky130_fd_sc_hd__o211a_1 _20064_ (.A1(_01241_),
    .A2(_01242_),
    .B1(_01016_),
    .C1(_01019_),
    .X(_01244_));
 sky130_fd_sc_hd__or2_1 _20065_ (.A(_01243_),
    .B(_01244_),
    .X(_01245_));
 sky130_fd_sc_hd__xnor2_1 _20066_ (.A(_01204_),
    .B(_01245_),
    .Y(_01246_));
 sky130_fd_sc_hd__a21o_1 _20067_ (.A1(_01024_),
    .A2(_01109_),
    .B1(_01108_),
    .X(_01247_));
 sky130_fd_sc_hd__and2b_1 _20068_ (.A_N(_01246_),
    .B(_01247_),
    .X(_01248_));
 sky130_fd_sc_hd__xnor2_1 _20069_ (.A(_01246_),
    .B(_01247_),
    .Y(_01249_));
 sky130_fd_sc_hd__xnor2_1 _20070_ (.A(_01129_),
    .B(_01249_),
    .Y(_01250_));
 sky130_fd_sc_hd__a21o_1 _20071_ (.A1(_01112_),
    .A2(_01114_),
    .B1(_01250_),
    .X(_01251_));
 sky130_fd_sc_hd__nand3_1 _20072_ (.A(_01112_),
    .B(_01114_),
    .C(_01250_),
    .Y(_01252_));
 sky130_fd_sc_hd__and2_1 _20073_ (.A(_01251_),
    .B(_01252_),
    .X(_01253_));
 sky130_fd_sc_hd__nand2_1 _20074_ (.A(_01128_),
    .B(_01253_),
    .Y(_01254_));
 sky130_fd_sc_hd__xnor2_1 _20075_ (.A(_01128_),
    .B(_01253_),
    .Y(_01255_));
 sky130_fd_sc_hd__a21oi_1 _20076_ (.A1(_00978_),
    .A2(_01118_),
    .B1(_01117_),
    .Y(_01256_));
 sky130_fd_sc_hd__or2_1 _20077_ (.A(_01255_),
    .B(_01256_),
    .X(_01257_));
 sky130_fd_sc_hd__nand2_1 _20078_ (.A(_01255_),
    .B(_01256_),
    .Y(_01258_));
 sky130_fd_sc_hd__nand2_1 _20079_ (.A(_01257_),
    .B(_01258_),
    .Y(_01259_));
 sky130_fd_sc_hd__a21o_1 _20080_ (.A1(_00966_),
    .A2(_01121_),
    .B1(_01123_),
    .X(_01260_));
 sky130_fd_sc_hd__nand2_1 _20081_ (.A(_00968_),
    .B(_01124_),
    .Y(_01261_));
 sky130_fd_sc_hd__o21a_1 _20082_ (.A1(_00972_),
    .A2(_01261_),
    .B1(_01260_),
    .X(_01262_));
 sky130_fd_sc_hd__xnor2_2 _20083_ (.A(_01259_),
    .B(_01262_),
    .Y(_01263_));
 sky130_fd_sc_hd__o22a_1 _20084_ (.A1(net44),
    .A2(_06691_),
    .B1(_01263_),
    .B2(_03049_),
    .X(_01264_));
 sky130_fd_sc_hd__a21bo_1 _20085_ (.A1(net684),
    .A2(net8),
    .B1_N(_01264_),
    .X(_01265_));
 sky130_fd_sc_hd__mux2_1 _20086_ (.A0(net696),
    .A1(_01265_),
    .S(net4),
    .X(_00320_));
 sky130_fd_sc_hd__nand2_1 _20087_ (.A(_01131_),
    .B(_01135_),
    .Y(_01266_));
 sky130_fd_sc_hd__nand2_1 _20088_ (.A(net158),
    .B(net193),
    .Y(_01267_));
 sky130_fd_sc_hd__xnor2_2 _20089_ (.A(_01133_),
    .B(_01267_),
    .Y(_01268_));
 sky130_fd_sc_hd__and2b_1 _20090_ (.A_N(_01268_),
    .B(_01031_),
    .X(_01269_));
 sky130_fd_sc_hd__xor2_2 _20091_ (.A(_01031_),
    .B(_01268_),
    .X(_01270_));
 sky130_fd_sc_hd__and2b_1 _20092_ (.A_N(_01270_),
    .B(_01266_),
    .X(_01271_));
 sky130_fd_sc_hd__xnor2_2 _20093_ (.A(_01266_),
    .B(_01270_),
    .Y(_01272_));
 sky130_fd_sc_hd__xnor2_2 _20094_ (.A(_01029_),
    .B(_01272_),
    .Y(_01273_));
 sky130_fd_sc_hd__nand2_1 _20095_ (.A(_01026_),
    .B(_01141_),
    .Y(_01274_));
 sky130_fd_sc_hd__nand2b_1 _20096_ (.A_N(_01273_),
    .B(_01274_),
    .Y(_01275_));
 sky130_fd_sc_hd__xnor2_2 _20097_ (.A(_01273_),
    .B(_01274_),
    .Y(_01276_));
 sky130_fd_sc_hd__nand2_1 _20098_ (.A(_01155_),
    .B(_01157_),
    .Y(_01277_));
 sky130_fd_sc_hd__a31o_1 _20099_ (.A1(_01031_),
    .A2(_01134_),
    .A3(_01135_),
    .B1(_01138_),
    .X(_01278_));
 sky130_fd_sc_hd__a22o_1 _20100_ (.A1(net134),
    .A2(\mul1.a[26] ),
    .B1(net202),
    .B2(net139),
    .X(_01279_));
 sky130_fd_sc_hd__nand4_2 _20101_ (.A(net139),
    .B(net134),
    .C(\mul1.a[26] ),
    .D(\mul1.a[27] ),
    .Y(_01280_));
 sky130_fd_sc_hd__a22o_1 _20102_ (.A1(net130),
    .A2(\mul1.a[25] ),
    .B1(_01279_),
    .B2(_01280_),
    .X(_01281_));
 sky130_fd_sc_hd__nand4_1 _20103_ (.A(net130),
    .B(\mul1.a[25] ),
    .C(_01279_),
    .D(_01280_),
    .Y(_01282_));
 sky130_fd_sc_hd__nand2_1 _20104_ (.A(_01281_),
    .B(_01282_),
    .Y(_01283_));
 sky130_fd_sc_hd__a22oi_1 _20105_ (.A1(\mul1.b[10] ),
    .A2(net197),
    .B1(net195),
    .B2(\mul1.b[9] ),
    .Y(_01284_));
 sky130_fd_sc_hd__and4_1 _20106_ (.A(\mul1.b[9] ),
    .B(\mul1.b[10] ),
    .C(net197),
    .D(net195),
    .X(_01285_));
 sky130_fd_sc_hd__o2bb2a_1 _20107_ (.A1_N(net142),
    .A2_N(net199),
    .B1(_01284_),
    .B2(_01285_),
    .X(_01286_));
 sky130_fd_sc_hd__and4bb_1 _20108_ (.A_N(_01284_),
    .B_N(_01285_),
    .C(net142),
    .D(net199),
    .X(_01287_));
 sky130_fd_sc_hd__nor2_1 _20109_ (.A(_01286_),
    .B(_01287_),
    .Y(_01288_));
 sky130_fd_sc_hd__nand2_1 _20110_ (.A(_01152_),
    .B(_01154_),
    .Y(_01289_));
 sky130_fd_sc_hd__nand2_1 _20111_ (.A(_01288_),
    .B(_01289_),
    .Y(_01290_));
 sky130_fd_sc_hd__xnor2_2 _20112_ (.A(_01288_),
    .B(_01289_),
    .Y(_01291_));
 sky130_fd_sc_hd__or2_1 _20113_ (.A(_01283_),
    .B(_01291_),
    .X(_01292_));
 sky130_fd_sc_hd__xor2_2 _20114_ (.A(_01283_),
    .B(_01291_),
    .X(_01293_));
 sky130_fd_sc_hd__and2_1 _20115_ (.A(_01278_),
    .B(_01293_),
    .X(_01294_));
 sky130_fd_sc_hd__xnor2_2 _20116_ (.A(_01278_),
    .B(_01293_),
    .Y(_01295_));
 sky130_fd_sc_hd__nand2b_1 _20117_ (.A_N(_01295_),
    .B(_01277_),
    .Y(_01296_));
 sky130_fd_sc_hd__inv_2 _20118_ (.A(_01296_),
    .Y(_01297_));
 sky130_fd_sc_hd__xnor2_2 _20119_ (.A(_01277_),
    .B(_01295_),
    .Y(_01298_));
 sky130_fd_sc_hd__nand2_1 _20120_ (.A(_01276_),
    .B(_01298_),
    .Y(_01299_));
 sky130_fd_sc_hd__xnor2_2 _20121_ (.A(_01276_),
    .B(_01298_),
    .Y(_01300_));
 sky130_fd_sc_hd__nand2b_1 _20122_ (.A_N(_01143_),
    .B(_01164_),
    .Y(_01301_));
 sky130_fd_sc_hd__nand2b_1 _20123_ (.A_N(_01300_),
    .B(_01301_),
    .Y(_01302_));
 sky130_fd_sc_hd__xnor2_2 _20124_ (.A(_01300_),
    .B(_01301_),
    .Y(_01303_));
 sky130_fd_sc_hd__and2_1 _20125_ (.A(_01192_),
    .B(_01194_),
    .X(_01304_));
 sky130_fd_sc_hd__nor2_1 _20126_ (.A(_01159_),
    .B(_01161_),
    .Y(_01305_));
 sky130_fd_sc_hd__a22o_1 _20127_ (.A1(net241),
    .A2(net95),
    .B1(net92),
    .B2(net245),
    .X(_01306_));
 sky130_fd_sc_hd__nand4_2 _20128_ (.A(net245),
    .B(net241),
    .C(net95),
    .D(net92),
    .Y(_01307_));
 sky130_fd_sc_hd__a22o_1 _20129_ (.A1(net628),
    .A2(net87),
    .B1(_01306_),
    .B2(_01307_),
    .X(_01308_));
 sky130_fd_sc_hd__nand4_1 _20130_ (.A(net628),
    .B(net87),
    .C(_01306_),
    .D(_01307_),
    .Y(_01309_));
 sky130_fd_sc_hd__nand2_1 _20131_ (.A(_01308_),
    .B(_01309_),
    .Y(_01310_));
 sky130_fd_sc_hd__a22o_1 _20132_ (.A1(net105),
    .A2(net231),
    .B1(net227),
    .B2(net110),
    .X(_01311_));
 sky130_fd_sc_hd__and4_1 _20133_ (.A(net110),
    .B(net105),
    .C(net231),
    .D(net227),
    .X(_01312_));
 sky130_fd_sc_hd__inv_2 _20134_ (.A(_01312_),
    .Y(_01313_));
 sky130_fd_sc_hd__a22oi_1 _20135_ (.A1(net236),
    .A2(net101),
    .B1(_01311_),
    .B2(_01313_),
    .Y(_01314_));
 sky130_fd_sc_hd__and4_1 _20136_ (.A(net236),
    .B(net101),
    .C(_01311_),
    .D(_01313_),
    .X(_01315_));
 sky130_fd_sc_hd__or2_1 _20137_ (.A(_01314_),
    .B(_01315_),
    .X(_01316_));
 sky130_fd_sc_hd__nand2_1 _20138_ (.A(_01173_),
    .B(_01175_),
    .Y(_01317_));
 sky130_fd_sc_hd__or3b_1 _20139_ (.A(_01314_),
    .B(_01315_),
    .C_N(_01317_),
    .X(_01318_));
 sky130_fd_sc_hd__xor2_2 _20140_ (.A(_01316_),
    .B(_01317_),
    .X(_01319_));
 sky130_fd_sc_hd__or2_1 _20141_ (.A(_01310_),
    .B(_01319_),
    .X(_01320_));
 sky130_fd_sc_hd__xor2_2 _20142_ (.A(_01310_),
    .B(_01319_),
    .X(_01321_));
 sky130_fd_sc_hd__or2_1 _20143_ (.A(_01184_),
    .B(_01186_),
    .X(_01322_));
 sky130_fd_sc_hd__o2bb2a_1 _20144_ (.A1_N(net205),
    .A2_N(_01147_),
    .B1(_01148_),
    .B2(_01149_),
    .X(_01323_));
 sky130_fd_sc_hd__a22oi_1 _20145_ (.A1(net121),
    .A2(net217),
    .B1(net213),
    .B2(net125),
    .Y(_01324_));
 sky130_fd_sc_hd__and4_1 _20146_ (.A(net126),
    .B(net120),
    .C(net217),
    .D(net213),
    .X(_01325_));
 sky130_fd_sc_hd__o2bb2a_1 _20147_ (.A1_N(net116),
    .A2_N(net222),
    .B1(_01324_),
    .B2(_01325_),
    .X(_01326_));
 sky130_fd_sc_hd__and4bb_1 _20148_ (.A_N(_01324_),
    .B_N(_01325_),
    .C(net116),
    .D(net222),
    .X(_01327_));
 sky130_fd_sc_hd__or2_1 _20149_ (.A(_01326_),
    .B(_01327_),
    .X(_01328_));
 sky130_fd_sc_hd__or2_1 _20150_ (.A(_01323_),
    .B(_01328_),
    .X(_01329_));
 sky130_fd_sc_hd__xor2_2 _20151_ (.A(_01323_),
    .B(_01328_),
    .X(_01330_));
 sky130_fd_sc_hd__nand2_1 _20152_ (.A(_01322_),
    .B(_01330_),
    .Y(_01331_));
 sky130_fd_sc_hd__xnor2_2 _20153_ (.A(_01322_),
    .B(_01330_),
    .Y(_01332_));
 sky130_fd_sc_hd__nand2_1 _20154_ (.A(_01187_),
    .B(_01189_),
    .Y(_01333_));
 sky130_fd_sc_hd__and2b_1 _20155_ (.A_N(_01332_),
    .B(_01333_),
    .X(_01334_));
 sky130_fd_sc_hd__xnor2_2 _20156_ (.A(_01332_),
    .B(_01333_),
    .Y(_01335_));
 sky130_fd_sc_hd__xor2_2 _20157_ (.A(_01321_),
    .B(_01335_),
    .X(_01336_));
 sky130_fd_sc_hd__nand2b_1 _20158_ (.A_N(_01305_),
    .B(_01336_),
    .Y(_01337_));
 sky130_fd_sc_hd__xnor2_2 _20159_ (.A(_01305_),
    .B(_01336_),
    .Y(_01338_));
 sky130_fd_sc_hd__nand2b_1 _20160_ (.A_N(_01304_),
    .B(_01338_),
    .Y(_01339_));
 sky130_fd_sc_hd__xnor2_2 _20161_ (.A(_01304_),
    .B(_01338_),
    .Y(_01340_));
 sky130_fd_sc_hd__nand2_1 _20162_ (.A(_01303_),
    .B(_01340_),
    .Y(_01341_));
 sky130_fd_sc_hd__xnor2_2 _20163_ (.A(_01303_),
    .B(_01340_),
    .Y(_01342_));
 sky130_fd_sc_hd__nor2_1 _20164_ (.A(_01166_),
    .B(_01200_),
    .Y(_01343_));
 sky130_fd_sc_hd__nor2_2 _20165_ (.A(_01342_),
    .B(_01343_),
    .Y(_01344_));
 sky130_fd_sc_hd__xnor2_2 _20166_ (.A(_01342_),
    .B(_01343_),
    .Y(_01345_));
 sky130_fd_sc_hd__or2_1 _20167_ (.A(_01237_),
    .B(_01239_),
    .X(_01346_));
 sky130_fd_sc_hd__nand2_1 _20168_ (.A(_01196_),
    .B(_01198_),
    .Y(_01347_));
 sky130_fd_sc_hd__a22o_1 _20169_ (.A1(net265),
    .A2(net73),
    .B1(net70),
    .B2(net269),
    .X(_01348_));
 sky130_fd_sc_hd__and4_1 _20170_ (.A(net265),
    .B(net269),
    .C(net73),
    .D(net70),
    .X(_01349_));
 sky130_fd_sc_hd__inv_2 _20171_ (.A(_01349_),
    .Y(_01350_));
 sky130_fd_sc_hd__a22oi_1 _20172_ (.A1(net275),
    .A2(net67),
    .B1(_01348_),
    .B2(_01350_),
    .Y(_01351_));
 sky130_fd_sc_hd__and4_1 _20173_ (.A(net276),
    .B(net67),
    .C(_01348_),
    .D(_01350_),
    .X(_01352_));
 sky130_fd_sc_hd__or2_1 _20174_ (.A(_01351_),
    .B(_01352_),
    .X(_01353_));
 sky130_fd_sc_hd__or2_1 _20175_ (.A(_01206_),
    .B(_01208_),
    .X(_01354_));
 sky130_fd_sc_hd__or3b_1 _20176_ (.A(_01351_),
    .B(_01352_),
    .C_N(_01354_),
    .X(_01355_));
 sky130_fd_sc_hd__xor2_2 _20177_ (.A(_01353_),
    .B(_01354_),
    .X(_01356_));
 sky130_fd_sc_hd__and4b_2 _20178_ (.A_N(net285),
    .B(net64),
    .C(net62),
    .D(net280),
    .X(_01357_));
 sky130_fd_sc_hd__o2bb2a_1 _20179_ (.A1_N(net281),
    .A2_N(net64),
    .B1(net56),
    .B2(net285),
    .X(_01358_));
 sky130_fd_sc_hd__nor2_1 _20180_ (.A(_01357_),
    .B(_01358_),
    .Y(_01359_));
 sky130_fd_sc_hd__xnor2_1 _20181_ (.A(_01356_),
    .B(_01359_),
    .Y(_01360_));
 sky130_fd_sc_hd__o31ai_2 _20182_ (.A1(_01209_),
    .A2(_01212_),
    .A3(_01214_),
    .B1(_01210_),
    .Y(_01361_));
 sky130_fd_sc_hd__nand2_1 _20183_ (.A(_01360_),
    .B(_01361_),
    .Y(_01362_));
 sky130_fd_sc_hd__xnor2_1 _20184_ (.A(_01360_),
    .B(_01361_),
    .Y(_01363_));
 sky130_fd_sc_hd__xnor2_1 _20185_ (.A(_01213_),
    .B(_01363_),
    .Y(_01364_));
 sky130_fd_sc_hd__nand2_1 _20186_ (.A(_01229_),
    .B(_01231_),
    .Y(_01365_));
 sky130_fd_sc_hd__o21a_1 _20187_ (.A1(_01171_),
    .A2(_01179_),
    .B1(_01177_),
    .X(_01366_));
 sky130_fd_sc_hd__or2_1 _20188_ (.A(_01226_),
    .B(_01228_),
    .X(_01367_));
 sky130_fd_sc_hd__a32oi_4 _20189_ (.A1(net250),
    .A2(net87),
    .A3(_01167_),
    .B1(_01168_),
    .B2(net96),
    .Y(_01368_));
 sky130_fd_sc_hd__a22oi_1 _20190_ (.A1(net250),
    .A2(net84),
    .B1(net80),
    .B2(net255),
    .Y(_01369_));
 sky130_fd_sc_hd__and4_1 _20191_ (.A(net250),
    .B(net255),
    .C(net84),
    .D(net80),
    .X(_01370_));
 sky130_fd_sc_hd__o2bb2a_1 _20192_ (.A1_N(net261),
    .A2_N(net77),
    .B1(_01369_),
    .B2(_01370_),
    .X(_01371_));
 sky130_fd_sc_hd__and4bb_1 _20193_ (.A_N(_01369_),
    .B_N(_01370_),
    .C(net261),
    .D(net77),
    .X(_01372_));
 sky130_fd_sc_hd__or2_1 _20194_ (.A(_01371_),
    .B(_01372_),
    .X(_01373_));
 sky130_fd_sc_hd__or2_1 _20195_ (.A(_01368_),
    .B(_01373_),
    .X(_01374_));
 sky130_fd_sc_hd__xor2_1 _20196_ (.A(_01368_),
    .B(_01373_),
    .X(_01375_));
 sky130_fd_sc_hd__nand2_1 _20197_ (.A(_01367_),
    .B(_01375_),
    .Y(_01376_));
 sky130_fd_sc_hd__xnor2_1 _20198_ (.A(_01367_),
    .B(_01375_),
    .Y(_01377_));
 sky130_fd_sc_hd__nor2_1 _20199_ (.A(_01366_),
    .B(_01377_),
    .Y(_01378_));
 sky130_fd_sc_hd__xor2_1 _20200_ (.A(_01366_),
    .B(_01377_),
    .X(_01379_));
 sky130_fd_sc_hd__and2_1 _20201_ (.A(_01365_),
    .B(_01379_),
    .X(_01380_));
 sky130_fd_sc_hd__xnor2_1 _20202_ (.A(_01365_),
    .B(_01379_),
    .Y(_01381_));
 sky130_fd_sc_hd__and2b_1 _20203_ (.A_N(_01233_),
    .B(_01235_),
    .X(_01382_));
 sky130_fd_sc_hd__or2_1 _20204_ (.A(_01381_),
    .B(_01382_),
    .X(_01383_));
 sky130_fd_sc_hd__xnor2_1 _20205_ (.A(_01381_),
    .B(_01382_),
    .Y(_01384_));
 sky130_fd_sc_hd__xnor2_1 _20206_ (.A(_01364_),
    .B(_01384_),
    .Y(_01385_));
 sky130_fd_sc_hd__and2b_1 _20207_ (.A_N(_01385_),
    .B(_01347_),
    .X(_01386_));
 sky130_fd_sc_hd__xnor2_1 _20208_ (.A(_01347_),
    .B(_01385_),
    .Y(_01387_));
 sky130_fd_sc_hd__and2_1 _20209_ (.A(_01346_),
    .B(_01387_),
    .X(_01388_));
 sky130_fd_sc_hd__xnor2_1 _20210_ (.A(_01346_),
    .B(_01387_),
    .Y(_01389_));
 sky130_fd_sc_hd__nor2_1 _20211_ (.A(_01345_),
    .B(_01389_),
    .Y(_01390_));
 sky130_fd_sc_hd__xnor2_1 _20212_ (.A(_01345_),
    .B(_01389_),
    .Y(_01391_));
 sky130_fd_sc_hd__o21ai_1 _20213_ (.A1(_01204_),
    .A2(_01245_),
    .B1(_01202_),
    .Y(_01392_));
 sky130_fd_sc_hd__and2b_1 _20214_ (.A_N(_01391_),
    .B(_01392_),
    .X(_01393_));
 sky130_fd_sc_hd__xor2_1 _20215_ (.A(_01391_),
    .B(_01392_),
    .X(_01394_));
 sky130_fd_sc_hd__nor2_1 _20216_ (.A(_01241_),
    .B(_01243_),
    .Y(_01395_));
 sky130_fd_sc_hd__nor2_1 _20217_ (.A(_01394_),
    .B(_01395_),
    .Y(_01396_));
 sky130_fd_sc_hd__xnor2_1 _20218_ (.A(_01394_),
    .B(_01395_),
    .Y(_01397_));
 sky130_fd_sc_hd__a21oi_1 _20219_ (.A1(_01129_),
    .A2(_01249_),
    .B1(_01248_),
    .Y(_01398_));
 sky130_fd_sc_hd__xnor2_1 _20220_ (.A(_01397_),
    .B(_01398_),
    .Y(_01399_));
 sky130_fd_sc_hd__o21ba_1 _20221_ (.A1(_01218_),
    .A2(_01220_),
    .B1_N(_01399_),
    .X(_01400_));
 sky130_fd_sc_hd__or3b_1 _20222_ (.A(_01218_),
    .B(_01220_),
    .C_N(_01399_),
    .X(_01401_));
 sky130_fd_sc_hd__nand2b_1 _20223_ (.A_N(_01400_),
    .B(_01401_),
    .Y(_01402_));
 sky130_fd_sc_hd__and3_1 _20224_ (.A(_01251_),
    .B(_01254_),
    .C(_01402_),
    .X(_01403_));
 sky130_fd_sc_hd__a21o_1 _20225_ (.A1(_01251_),
    .A2(_01254_),
    .B1(_01402_),
    .X(_01404_));
 sky130_fd_sc_hd__nand2b_1 _20226_ (.A_N(_01403_),
    .B(_01404_),
    .Y(_01405_));
 sky130_fd_sc_hd__o21a_1 _20227_ (.A1(_01259_),
    .A2(_01262_),
    .B1(_01257_),
    .X(_01406_));
 sky130_fd_sc_hd__xnor2_2 _20228_ (.A(_01405_),
    .B(_01406_),
    .Y(_01407_));
 sky130_fd_sc_hd__nor2_1 _20229_ (.A(_03049_),
    .B(_01407_),
    .Y(_01408_));
 sky130_fd_sc_hd__a221o_1 _20230_ (.A1(\temp[22] ),
    .A2(net7),
    .B1(_06837_),
    .B2(_03052_),
    .C1(_01408_),
    .X(_01409_));
 sky130_fd_sc_hd__mux2_1 _20231_ (.A0(net804),
    .A1(_01409_),
    .S(net4),
    .X(_00321_));
 sky130_fd_sc_hd__a21o_1 _20232_ (.A1(_01029_),
    .A2(_01272_),
    .B1(_01025_),
    .X(_01410_));
 sky130_fd_sc_hd__o21a_1 _20233_ (.A1(_01133_),
    .A2(_01267_),
    .B1(_01131_),
    .X(_01411_));
 sky130_fd_sc_hd__nor2_1 _20234_ (.A(_01270_),
    .B(_01411_),
    .Y(_01412_));
 sky130_fd_sc_hd__and2_1 _20235_ (.A(_01270_),
    .B(_01411_),
    .X(_01413_));
 sky130_fd_sc_hd__or2_2 _20236_ (.A(_01412_),
    .B(_01413_),
    .X(_01414_));
 sky130_fd_sc_hd__xor2_2 _20237_ (.A(_01029_),
    .B(_01414_),
    .X(_01415_));
 sky130_fd_sc_hd__inv_2 _20238_ (.A(_01415_),
    .Y(_01416_));
 sky130_fd_sc_hd__xnor2_1 _20239_ (.A(_01410_),
    .B(_01415_),
    .Y(_01417_));
 sky130_fd_sc_hd__or2_1 _20240_ (.A(_01269_),
    .B(_01271_),
    .X(_01418_));
 sky130_fd_sc_hd__a22o_1 _20241_ (.A1(net132),
    .A2(net202),
    .B1(net199),
    .B2(net137),
    .X(_01419_));
 sky130_fd_sc_hd__nand4_2 _20242_ (.A(net137),
    .B(net132),
    .C(net202),
    .D(net199),
    .Y(_01420_));
 sky130_fd_sc_hd__a22o_1 _20243_ (.A1(net128),
    .A2(net207),
    .B1(_01419_),
    .B2(_01420_),
    .X(_01421_));
 sky130_fd_sc_hd__nand4_2 _20244_ (.A(net128),
    .B(net207),
    .C(_01419_),
    .D(_01420_),
    .Y(_01422_));
 sky130_fd_sc_hd__nand2_1 _20245_ (.A(_01421_),
    .B(_01422_),
    .Y(_01423_));
 sky130_fd_sc_hd__a22oi_1 _20246_ (.A1(\mul1.b[10] ),
    .A2(net195),
    .B1(net193),
    .B2(\mul1.b[9] ),
    .Y(_01424_));
 sky130_fd_sc_hd__and4_1 _20247_ (.A(\mul1.b[9] ),
    .B(\mul1.b[10] ),
    .C(net195),
    .D(net193),
    .X(_01425_));
 sky130_fd_sc_hd__nor2_1 _20248_ (.A(_01424_),
    .B(_01425_),
    .Y(_01426_));
 sky130_fd_sc_hd__nand2_1 _20249_ (.A(net142),
    .B(net197),
    .Y(_01427_));
 sky130_fd_sc_hd__xor2_1 _20250_ (.A(_01426_),
    .B(_01427_),
    .X(_01428_));
 sky130_fd_sc_hd__nor2_1 _20251_ (.A(_01285_),
    .B(_01287_),
    .Y(_01429_));
 sky130_fd_sc_hd__nor2_1 _20252_ (.A(_01428_),
    .B(_01429_),
    .Y(_01430_));
 sky130_fd_sc_hd__nand2_1 _20253_ (.A(_01428_),
    .B(_01429_),
    .Y(_01431_));
 sky130_fd_sc_hd__nand2b_1 _20254_ (.A_N(_01430_),
    .B(_01431_),
    .Y(_01432_));
 sky130_fd_sc_hd__xor2_1 _20255_ (.A(_01423_),
    .B(_01432_),
    .X(_01433_));
 sky130_fd_sc_hd__xnor2_1 _20256_ (.A(_01418_),
    .B(_01433_),
    .Y(_01434_));
 sky130_fd_sc_hd__a21o_1 _20257_ (.A1(_01290_),
    .A2(_01292_),
    .B1(_01434_),
    .X(_01435_));
 sky130_fd_sc_hd__nand3_1 _20258_ (.A(_01290_),
    .B(_01292_),
    .C(_01434_),
    .Y(_01436_));
 sky130_fd_sc_hd__a21oi_2 _20259_ (.A1(_01435_),
    .A2(_01436_),
    .B1(_01417_),
    .Y(_01437_));
 sky130_fd_sc_hd__and3_1 _20260_ (.A(_01417_),
    .B(_01435_),
    .C(_01436_),
    .X(_01438_));
 sky130_fd_sc_hd__o211a_1 _20261_ (.A1(_01437_),
    .A2(_01438_),
    .B1(_01275_),
    .C1(_01299_),
    .X(_01439_));
 sky130_fd_sc_hd__a211oi_4 _20262_ (.A1(_01275_),
    .A2(_01299_),
    .B1(_01437_),
    .C1(_01438_),
    .Y(_01440_));
 sky130_fd_sc_hd__a21o_1 _20263_ (.A1(_01321_),
    .A2(_01335_),
    .B1(_01334_),
    .X(_01441_));
 sky130_fd_sc_hd__a22o_1 _20264_ (.A1(net236),
    .A2(net95),
    .B1(net91),
    .B2(net241),
    .X(_01442_));
 sky130_fd_sc_hd__nand4_1 _20265_ (.A(net241),
    .B(net236),
    .C(net95),
    .D(net92),
    .Y(_01443_));
 sky130_fd_sc_hd__a22o_1 _20266_ (.A1(net246),
    .A2(net86),
    .B1(_01442_),
    .B2(_01443_),
    .X(_01444_));
 sky130_fd_sc_hd__nand4_1 _20267_ (.A(net245),
    .B(net86),
    .C(_01442_),
    .D(_01443_),
    .Y(_01445_));
 sky130_fd_sc_hd__nand2_1 _20268_ (.A(_01444_),
    .B(_01445_),
    .Y(_01446_));
 sky130_fd_sc_hd__a22o_1 _20269_ (.A1(net105),
    .A2(net227),
    .B1(net222),
    .B2(net110),
    .X(_01447_));
 sky130_fd_sc_hd__and4_1 _20270_ (.A(net110),
    .B(net105),
    .C(net227),
    .D(net222),
    .X(_01448_));
 sky130_fd_sc_hd__inv_2 _20271_ (.A(_01448_),
    .Y(_01449_));
 sky130_fd_sc_hd__a22oi_1 _20272_ (.A1(net231),
    .A2(net101),
    .B1(_01447_),
    .B2(_01449_),
    .Y(_01450_));
 sky130_fd_sc_hd__and4_1 _20273_ (.A(net231),
    .B(net101),
    .C(_01447_),
    .D(_01449_),
    .X(_01451_));
 sky130_fd_sc_hd__or2_1 _20274_ (.A(_01450_),
    .B(_01451_),
    .X(_01452_));
 sky130_fd_sc_hd__or2_1 _20275_ (.A(_01312_),
    .B(_01315_),
    .X(_01453_));
 sky130_fd_sc_hd__nand2b_1 _20276_ (.A_N(_01452_),
    .B(_01453_),
    .Y(_01454_));
 sky130_fd_sc_hd__xor2_1 _20277_ (.A(_01452_),
    .B(_01453_),
    .X(_01455_));
 sky130_fd_sc_hd__or2_1 _20278_ (.A(_01446_),
    .B(_01455_),
    .X(_01456_));
 sky130_fd_sc_hd__nand2_1 _20279_ (.A(_01446_),
    .B(_01455_),
    .Y(_01457_));
 sky130_fd_sc_hd__and2_1 _20280_ (.A(_01456_),
    .B(_01457_),
    .X(_01458_));
 sky130_fd_sc_hd__or2_1 _20281_ (.A(_01325_),
    .B(_01327_),
    .X(_01459_));
 sky130_fd_sc_hd__nand2_1 _20282_ (.A(_01280_),
    .B(_01282_),
    .Y(_01460_));
 sky130_fd_sc_hd__a22o_1 _20283_ (.A1(net121),
    .A2(net213),
    .B1(net210),
    .B2(net126),
    .X(_01461_));
 sky130_fd_sc_hd__inv_2 _20284_ (.A(_01461_),
    .Y(_01462_));
 sky130_fd_sc_hd__and4_1 _20285_ (.A(net126),
    .B(net121),
    .C(net213),
    .D(net210),
    .X(_01463_));
 sky130_fd_sc_hd__o2bb2a_1 _20286_ (.A1_N(\mul1.b[17] ),
    .A2_N(net217),
    .B1(_01462_),
    .B2(_01463_),
    .X(_01464_));
 sky130_fd_sc_hd__and4b_1 _20287_ (.A_N(_01463_),
    .B(net217),
    .C(net113),
    .D(_01461_),
    .X(_01465_));
 sky130_fd_sc_hd__or2_1 _20288_ (.A(_01464_),
    .B(_01465_),
    .X(_01466_));
 sky130_fd_sc_hd__nand2b_1 _20289_ (.A_N(_01466_),
    .B(_01460_),
    .Y(_01467_));
 sky130_fd_sc_hd__xnor2_1 _20290_ (.A(_01460_),
    .B(_01466_),
    .Y(_01468_));
 sky130_fd_sc_hd__nand2_1 _20291_ (.A(_01459_),
    .B(_01468_),
    .Y(_01469_));
 sky130_fd_sc_hd__xnor2_1 _20292_ (.A(_01459_),
    .B(_01468_),
    .Y(_01470_));
 sky130_fd_sc_hd__a21o_1 _20293_ (.A1(_01329_),
    .A2(_01331_),
    .B1(_01470_),
    .X(_01471_));
 sky130_fd_sc_hd__nand3_1 _20294_ (.A(_01329_),
    .B(_01331_),
    .C(_01470_),
    .Y(_01472_));
 sky130_fd_sc_hd__nand3_2 _20295_ (.A(_01458_),
    .B(_01471_),
    .C(_01472_),
    .Y(_01473_));
 sky130_fd_sc_hd__a21o_1 _20296_ (.A1(_01471_),
    .A2(_01472_),
    .B1(_01458_),
    .X(_01474_));
 sky130_fd_sc_hd__o211a_1 _20297_ (.A1(_01294_),
    .A2(_01297_),
    .B1(_01473_),
    .C1(_01474_),
    .X(_01475_));
 sky130_fd_sc_hd__a211oi_1 _20298_ (.A1(_01473_),
    .A2(_01474_),
    .B1(_01294_),
    .C1(_01297_),
    .Y(_01476_));
 sky130_fd_sc_hd__nor2_1 _20299_ (.A(_01475_),
    .B(_01476_),
    .Y(_01477_));
 sky130_fd_sc_hd__and2_1 _20300_ (.A(_01441_),
    .B(_01477_),
    .X(_01478_));
 sky130_fd_sc_hd__xnor2_2 _20301_ (.A(_01441_),
    .B(_01477_),
    .Y(_01479_));
 sky130_fd_sc_hd__nor3_4 _20302_ (.A(_01439_),
    .B(_01440_),
    .C(_01479_),
    .Y(_01480_));
 sky130_fd_sc_hd__o21a_1 _20303_ (.A1(_01439_),
    .A2(_01440_),
    .B1(_01479_),
    .X(_01481_));
 sky130_fd_sc_hd__a211o_2 _20304_ (.A1(_01302_),
    .A2(_01341_),
    .B1(_01480_),
    .C1(_01481_),
    .X(_01482_));
 sky130_fd_sc_hd__o211ai_4 _20305_ (.A1(_01480_),
    .A2(_01481_),
    .B1(_01302_),
    .C1(_01341_),
    .Y(_01483_));
 sky130_fd_sc_hd__o21a_1 _20306_ (.A1(_01364_),
    .A2(_01384_),
    .B1(_01383_),
    .X(_01484_));
 sky130_fd_sc_hd__nand2_1 _20307_ (.A(_01337_),
    .B(_01339_),
    .Y(_01485_));
 sky130_fd_sc_hd__a22o_1 _20308_ (.A1(net261),
    .A2(net72),
    .B1(net69),
    .B2(net265),
    .X(_01486_));
 sky130_fd_sc_hd__and4_1 _20309_ (.A(net261),
    .B(net265),
    .C(net72),
    .D(net69),
    .X(_01487_));
 sky130_fd_sc_hd__inv_2 _20310_ (.A(_01487_),
    .Y(_01488_));
 sky130_fd_sc_hd__a22oi_1 _20311_ (.A1(net269),
    .A2(net66),
    .B1(_01486_),
    .B2(_01488_),
    .Y(_01489_));
 sky130_fd_sc_hd__and4_1 _20312_ (.A(net269),
    .B(net66),
    .C(_01486_),
    .D(_01488_),
    .X(_01490_));
 sky130_fd_sc_hd__or2_1 _20313_ (.A(_01489_),
    .B(_01490_),
    .X(_01491_));
 sky130_fd_sc_hd__or2_1 _20314_ (.A(_01349_),
    .B(_01352_),
    .X(_01492_));
 sky130_fd_sc_hd__and2b_1 _20315_ (.A_N(_01491_),
    .B(_01492_),
    .X(_01493_));
 sky130_fd_sc_hd__xor2_1 _20316_ (.A(_01491_),
    .B(_01492_),
    .X(_01494_));
 sky130_fd_sc_hd__and4b_1 _20317_ (.A_N(net280),
    .B(net63),
    .C(net62),
    .D(net276),
    .X(_01495_));
 sky130_fd_sc_hd__inv_2 _20318_ (.A(_01495_),
    .Y(_01496_));
 sky130_fd_sc_hd__o2bb2a_1 _20319_ (.A1_N(net276),
    .A2_N(net64),
    .B1(net56),
    .B2(net281),
    .X(_01497_));
 sky130_fd_sc_hd__o21a_1 _20320_ (.A1(_01495_),
    .A2(_01497_),
    .B1(_01494_),
    .X(_01498_));
 sky130_fd_sc_hd__nor3_1 _20321_ (.A(_01494_),
    .B(_01495_),
    .C(_01497_),
    .Y(_01499_));
 sky130_fd_sc_hd__nor2_1 _20322_ (.A(_01498_),
    .B(_01499_),
    .Y(_01500_));
 sky130_fd_sc_hd__o31ai_2 _20323_ (.A1(_01356_),
    .A2(_01357_),
    .A3(_01358_),
    .B1(_01355_),
    .Y(_01501_));
 sky130_fd_sc_hd__nand2_1 _20324_ (.A(_01500_),
    .B(_01501_),
    .Y(_01502_));
 sky130_fd_sc_hd__xnor2_1 _20325_ (.A(_01500_),
    .B(_01501_),
    .Y(_01503_));
 sky130_fd_sc_hd__inv_2 _20326_ (.A(_01503_),
    .Y(_01504_));
 sky130_fd_sc_hd__nand2_1 _20327_ (.A(_01357_),
    .B(_01504_),
    .Y(_01505_));
 sky130_fd_sc_hd__xor2_1 _20328_ (.A(_01357_),
    .B(_01503_),
    .X(_01506_));
 sky130_fd_sc_hd__or2_1 _20329_ (.A(_01370_),
    .B(_01372_),
    .X(_01507_));
 sky130_fd_sc_hd__nand2_1 _20330_ (.A(_01307_),
    .B(_01309_),
    .Y(_01508_));
 sky130_fd_sc_hd__a22o_1 _20331_ (.A1(net628),
    .A2(net83),
    .B1(net79),
    .B2(net250),
    .X(_01509_));
 sky130_fd_sc_hd__inv_2 _20332_ (.A(_01509_),
    .Y(_01510_));
 sky130_fd_sc_hd__and4_1 _20333_ (.A(net628),
    .B(net250),
    .C(net83),
    .D(net79),
    .X(_01511_));
 sky130_fd_sc_hd__o2bb2a_1 _20334_ (.A1_N(net255),
    .A2_N(net76),
    .B1(_01510_),
    .B2(_01511_),
    .X(_01512_));
 sky130_fd_sc_hd__and4b_1 _20335_ (.A_N(_01511_),
    .B(net76),
    .C(net255),
    .D(_01509_),
    .X(_01513_));
 sky130_fd_sc_hd__or2_1 _20336_ (.A(_01512_),
    .B(_01513_),
    .X(_01514_));
 sky130_fd_sc_hd__nand2b_1 _20337_ (.A_N(_01514_),
    .B(_01508_),
    .Y(_01515_));
 sky130_fd_sc_hd__xnor2_1 _20338_ (.A(_01508_),
    .B(_01514_),
    .Y(_01516_));
 sky130_fd_sc_hd__nand2_1 _20339_ (.A(_01507_),
    .B(_01516_),
    .Y(_01517_));
 sky130_fd_sc_hd__xnor2_1 _20340_ (.A(_01507_),
    .B(_01516_),
    .Y(_01518_));
 sky130_fd_sc_hd__a21oi_1 _20341_ (.A1(_01318_),
    .A2(_01320_),
    .B1(_01518_),
    .Y(_01519_));
 sky130_fd_sc_hd__a21o_1 _20342_ (.A1(_01318_),
    .A2(_01320_),
    .B1(_01518_),
    .X(_01520_));
 sky130_fd_sc_hd__and3_1 _20343_ (.A(_01318_),
    .B(_01320_),
    .C(_01518_),
    .X(_01521_));
 sky130_fd_sc_hd__a211o_2 _20344_ (.A1(_01374_),
    .A2(_01376_),
    .B1(_01519_),
    .C1(_01521_),
    .X(_01522_));
 sky130_fd_sc_hd__o211ai_2 _20345_ (.A1(_01519_),
    .A2(_01521_),
    .B1(_01374_),
    .C1(_01376_),
    .Y(_01523_));
 sky130_fd_sc_hd__o211a_1 _20346_ (.A1(_01378_),
    .A2(_01380_),
    .B1(_01522_),
    .C1(_01523_),
    .X(_01524_));
 sky130_fd_sc_hd__a211oi_1 _20347_ (.A1(_01522_),
    .A2(_01523_),
    .B1(_01378_),
    .C1(_01380_),
    .Y(_01525_));
 sky130_fd_sc_hd__nor3_1 _20348_ (.A(_01506_),
    .B(_01524_),
    .C(_01525_),
    .Y(_01526_));
 sky130_fd_sc_hd__o21a_1 _20349_ (.A1(_01524_),
    .A2(_01525_),
    .B1(_01506_),
    .X(_01527_));
 sky130_fd_sc_hd__nor2_1 _20350_ (.A(_01526_),
    .B(_01527_),
    .Y(_01528_));
 sky130_fd_sc_hd__nand2_1 _20351_ (.A(_01485_),
    .B(_01528_),
    .Y(_01529_));
 sky130_fd_sc_hd__xnor2_1 _20352_ (.A(_01485_),
    .B(_01528_),
    .Y(_01530_));
 sky130_fd_sc_hd__or2_1 _20353_ (.A(_01484_),
    .B(_01530_),
    .X(_01531_));
 sky130_fd_sc_hd__xnor2_1 _20354_ (.A(_01484_),
    .B(_01530_),
    .Y(_01532_));
 sky130_fd_sc_hd__nand3b_4 _20355_ (.A_N(_01532_),
    .B(_01483_),
    .C(_01482_),
    .Y(_01533_));
 sky130_fd_sc_hd__a21bo_1 _20356_ (.A1(_01482_),
    .A2(_01483_),
    .B1_N(_01532_),
    .X(_01534_));
 sky130_fd_sc_hd__o211ai_4 _20357_ (.A1(_01344_),
    .A2(_01390_),
    .B1(_01533_),
    .C1(_01534_),
    .Y(_01535_));
 sky130_fd_sc_hd__a211o_1 _20358_ (.A1(_01533_),
    .A2(_01534_),
    .B1(_01344_),
    .C1(_01390_),
    .X(_01536_));
 sky130_fd_sc_hd__o211ai_4 _20359_ (.A1(_01386_),
    .A2(_01388_),
    .B1(_01535_),
    .C1(_01536_),
    .Y(_01537_));
 sky130_fd_sc_hd__a211o_1 _20360_ (.A1(_01535_),
    .A2(_01536_),
    .B1(_01386_),
    .C1(_01388_),
    .X(_01538_));
 sky130_fd_sc_hd__o211ai_2 _20361_ (.A1(_01393_),
    .A2(_01396_),
    .B1(_01537_),
    .C1(_01538_),
    .Y(_01539_));
 sky130_fd_sc_hd__a211o_1 _20362_ (.A1(_01537_),
    .A2(_01538_),
    .B1(_01393_),
    .C1(_01396_),
    .X(_01540_));
 sky130_fd_sc_hd__and2_1 _20363_ (.A(_01539_),
    .B(_01540_),
    .X(_01541_));
 sky130_fd_sc_hd__o21ai_1 _20364_ (.A1(_01213_),
    .A2(_01363_),
    .B1(_01362_),
    .Y(_01542_));
 sky130_fd_sc_hd__nand2_1 _20365_ (.A(_01541_),
    .B(_01542_),
    .Y(_01543_));
 sky130_fd_sc_hd__or2_1 _20366_ (.A(_01541_),
    .B(_01542_),
    .X(_01544_));
 sky130_fd_sc_hd__nand2_1 _20367_ (.A(_01543_),
    .B(_01544_),
    .Y(_01545_));
 sky130_fd_sc_hd__o21ba_1 _20368_ (.A1(_01397_),
    .A2(_01398_),
    .B1_N(_01400_),
    .X(_01546_));
 sky130_fd_sc_hd__nor2_1 _20369_ (.A(_01545_),
    .B(_01546_),
    .Y(_01547_));
 sky130_fd_sc_hd__and2_1 _20370_ (.A(_01545_),
    .B(_01546_),
    .X(_01548_));
 sky130_fd_sc_hd__nor2_1 _20371_ (.A(_01547_),
    .B(_01548_),
    .Y(_01549_));
 sky130_fd_sc_hd__or2_1 _20372_ (.A(_01259_),
    .B(_01405_),
    .X(_01550_));
 sky130_fd_sc_hd__o221a_1 _20373_ (.A1(_01257_),
    .A2(_01403_),
    .B1(_01550_),
    .B2(_01260_),
    .C1(_01404_),
    .X(_01551_));
 sky130_fd_sc_hd__o31a_2 _20374_ (.A1(_00972_),
    .A2(_01261_),
    .A3(_01550_),
    .B1(_01551_),
    .X(_01552_));
 sky130_fd_sc_hd__and2b_1 _20375_ (.A_N(_01552_),
    .B(_01549_),
    .X(_01553_));
 sky130_fd_sc_hd__xor2_1 _20376_ (.A(_01549_),
    .B(_01552_),
    .X(_01554_));
 sky130_fd_sc_hd__nor2_1 _20377_ (.A(_03049_),
    .B(_01554_),
    .Y(_01555_));
 sky130_fd_sc_hd__a221o_1 _20378_ (.A1(net741),
    .A2(net7),
    .B1(_06977_),
    .B2(_03052_),
    .C1(_01555_),
    .X(_01556_));
 sky130_fd_sc_hd__mux2_1 _20379_ (.A0(net747),
    .A1(_01556_),
    .S(net4),
    .X(_00322_));
 sky130_fd_sc_hd__nor2_4 _20380_ (.A(_01026_),
    .B(_01414_),
    .Y(_01557_));
 sky130_fd_sc_hd__and2_1 _20381_ (.A(_01027_),
    .B(_01414_),
    .X(_01558_));
 sky130_fd_sc_hd__nor2_2 _20382_ (.A(_01557_),
    .B(_01558_),
    .Y(_01559_));
 sky130_fd_sc_hd__or2_2 _20383_ (.A(_01557_),
    .B(_01558_),
    .X(_01560_));
 sky130_fd_sc_hd__a31o_1 _20384_ (.A1(_01421_),
    .A2(_01422_),
    .A3(_01431_),
    .B1(_01430_),
    .X(_01561_));
 sky130_fd_sc_hd__nor2_2 _20385_ (.A(_01269_),
    .B(_01412_),
    .Y(_01562_));
 sky130_fd_sc_hd__or2_4 _20386_ (.A(_01269_),
    .B(_01412_),
    .X(_01563_));
 sky130_fd_sc_hd__a22o_1 _20387_ (.A1(net132),
    .A2(net201),
    .B1(net198),
    .B2(net137),
    .X(_01564_));
 sky130_fd_sc_hd__nand4_2 _20388_ (.A(net137),
    .B(net132),
    .C(net201),
    .D(net198),
    .Y(_01565_));
 sky130_fd_sc_hd__a22o_1 _20389_ (.A1(net128),
    .A2(net204),
    .B1(_01564_),
    .B2(_01565_),
    .X(_01566_));
 sky130_fd_sc_hd__nand4_2 _20390_ (.A(net128),
    .B(net204),
    .C(_01564_),
    .D(_01565_),
    .Y(_01567_));
 sky130_fd_sc_hd__nand2_1 _20391_ (.A(_01566_),
    .B(_01567_),
    .Y(_01568_));
 sky130_fd_sc_hd__a31o_1 _20392_ (.A1(net142),
    .A2(net197),
    .A3(_01426_),
    .B1(_01425_),
    .X(_01569_));
 sky130_fd_sc_hd__nand2_1 _20393_ (.A(net143),
    .B(net196),
    .Y(_01570_));
 sky130_fd_sc_hd__and3_1 _20394_ (.A(\mul1.b[9] ),
    .B(net148),
    .C(net194),
    .X(_01571_));
 sky130_fd_sc_hd__o21a_1 _20395_ (.A1(net153),
    .A2(net148),
    .B1(net193),
    .X(_01572_));
 sky130_fd_sc_hd__and2b_1 _20396_ (.A_N(_01571_),
    .B(_01572_),
    .X(_01573_));
 sky130_fd_sc_hd__xnor2_1 _20397_ (.A(_01570_),
    .B(_01573_),
    .Y(_01574_));
 sky130_fd_sc_hd__xor2_1 _20398_ (.A(_01569_),
    .B(_01574_),
    .X(_01575_));
 sky130_fd_sc_hd__xnor2_1 _20399_ (.A(_01568_),
    .B(_01575_),
    .Y(_01576_));
 sky130_fd_sc_hd__and2_1 _20400_ (.A(_01563_),
    .B(_01576_),
    .X(_01577_));
 sky130_fd_sc_hd__xnor2_1 _20401_ (.A(_01563_),
    .B(_01576_),
    .Y(_01578_));
 sky130_fd_sc_hd__and2b_1 _20402_ (.A_N(_01578_),
    .B(_01561_),
    .X(_01579_));
 sky130_fd_sc_hd__xor2_1 _20403_ (.A(_01561_),
    .B(_01578_),
    .X(_01580_));
 sky130_fd_sc_hd__xnor2_1 _20404_ (.A(_01559_),
    .B(_01580_),
    .Y(_01581_));
 sky130_fd_sc_hd__a21o_1 _20405_ (.A1(_01410_),
    .A2(_01416_),
    .B1(_01438_),
    .X(_01582_));
 sky130_fd_sc_hd__or2_1 _20406_ (.A(_01581_),
    .B(_01582_),
    .X(_01583_));
 sky130_fd_sc_hd__nand2_2 _20407_ (.A(_01581_),
    .B(_01582_),
    .Y(_01584_));
 sky130_fd_sc_hd__nand2_1 _20408_ (.A(_01583_),
    .B(_01584_),
    .Y(_01585_));
 sky130_fd_sc_hd__a21bo_1 _20409_ (.A1(_01418_),
    .A2(_01433_),
    .B1_N(_01435_),
    .X(_01586_));
 sky130_fd_sc_hd__a22o_1 _20410_ (.A1(net230),
    .A2(net95),
    .B1(net91),
    .B2(net236),
    .X(_01587_));
 sky130_fd_sc_hd__nand4_2 _20411_ (.A(net236),
    .B(net230),
    .C(net95),
    .D(net91),
    .Y(_01588_));
 sky130_fd_sc_hd__a22o_1 _20412_ (.A1(net241),
    .A2(net86),
    .B1(_01587_),
    .B2(_01588_),
    .X(_01589_));
 sky130_fd_sc_hd__nand4_1 _20413_ (.A(net241),
    .B(net86),
    .C(_01587_),
    .D(_01588_),
    .Y(_01590_));
 sky130_fd_sc_hd__nand2_1 _20414_ (.A(_01589_),
    .B(_01590_),
    .Y(_01591_));
 sky130_fd_sc_hd__a22o_1 _20415_ (.A1(net105),
    .A2(net222),
    .B1(net217),
    .B2(net110),
    .X(_01592_));
 sky130_fd_sc_hd__and4_1 _20416_ (.A(net110),
    .B(net105),
    .C(net222),
    .D(net217),
    .X(_01593_));
 sky130_fd_sc_hd__inv_2 _20417_ (.A(_01593_),
    .Y(_01594_));
 sky130_fd_sc_hd__a22oi_1 _20418_ (.A1(\mul1.b[20] ),
    .A2(net227),
    .B1(_01592_),
    .B2(_01594_),
    .Y(_01595_));
 sky130_fd_sc_hd__and4_1 _20419_ (.A(net101),
    .B(net226),
    .C(_01592_),
    .D(_01594_),
    .X(_01596_));
 sky130_fd_sc_hd__or2_1 _20420_ (.A(_01595_),
    .B(_01596_),
    .X(_01597_));
 sky130_fd_sc_hd__or2_1 _20421_ (.A(_01448_),
    .B(_01451_),
    .X(_01598_));
 sky130_fd_sc_hd__nand2b_1 _20422_ (.A_N(_01597_),
    .B(_01598_),
    .Y(_01599_));
 sky130_fd_sc_hd__xor2_1 _20423_ (.A(_01597_),
    .B(_01598_),
    .X(_01600_));
 sky130_fd_sc_hd__or2_1 _20424_ (.A(_01591_),
    .B(_01600_),
    .X(_01601_));
 sky130_fd_sc_hd__nand2_1 _20425_ (.A(_01591_),
    .B(_01600_),
    .Y(_01602_));
 sky130_fd_sc_hd__and2_1 _20426_ (.A(_01601_),
    .B(_01602_),
    .X(_01603_));
 sky130_fd_sc_hd__or2_1 _20427_ (.A(_01463_),
    .B(_01465_),
    .X(_01604_));
 sky130_fd_sc_hd__nand2_1 _20428_ (.A(_01420_),
    .B(_01422_),
    .Y(_01605_));
 sky130_fd_sc_hd__a22o_1 _20429_ (.A1(net118),
    .A2(net210),
    .B1(net207),
    .B2(net123),
    .X(_01606_));
 sky130_fd_sc_hd__inv_2 _20430_ (.A(_01606_),
    .Y(_01607_));
 sky130_fd_sc_hd__and4_1 _20431_ (.A(net123),
    .B(net118),
    .C(net210),
    .D(net207),
    .X(_01608_));
 sky130_fd_sc_hd__o2bb2a_1 _20432_ (.A1_N(net113),
    .A2_N(net213),
    .B1(_01607_),
    .B2(_01608_),
    .X(_01609_));
 sky130_fd_sc_hd__and4b_1 _20433_ (.A_N(_01608_),
    .B(net214),
    .C(net113),
    .D(_01606_),
    .X(_01610_));
 sky130_fd_sc_hd__or2_1 _20434_ (.A(_01609_),
    .B(_01610_),
    .X(_01611_));
 sky130_fd_sc_hd__nand2b_1 _20435_ (.A_N(_01611_),
    .B(_01605_),
    .Y(_01612_));
 sky130_fd_sc_hd__xnor2_1 _20436_ (.A(_01605_),
    .B(_01611_),
    .Y(_01613_));
 sky130_fd_sc_hd__nand2_1 _20437_ (.A(_01604_),
    .B(_01613_),
    .Y(_01614_));
 sky130_fd_sc_hd__xnor2_1 _20438_ (.A(_01604_),
    .B(_01613_),
    .Y(_01615_));
 sky130_fd_sc_hd__a21o_1 _20439_ (.A1(_01467_),
    .A2(_01469_),
    .B1(_01615_),
    .X(_01616_));
 sky130_fd_sc_hd__nand3_1 _20440_ (.A(_01467_),
    .B(_01469_),
    .C(_01615_),
    .Y(_01617_));
 sky130_fd_sc_hd__and3_1 _20441_ (.A(_01603_),
    .B(_01616_),
    .C(_01617_),
    .X(_01618_));
 sky130_fd_sc_hd__inv_2 _20442_ (.A(_01618_),
    .Y(_01619_));
 sky130_fd_sc_hd__a21oi_1 _20443_ (.A1(_01616_),
    .A2(_01617_),
    .B1(_01603_),
    .Y(_01620_));
 sky130_fd_sc_hd__nor2_1 _20444_ (.A(_01618_),
    .B(_01620_),
    .Y(_01621_));
 sky130_fd_sc_hd__nand2_2 _20445_ (.A(_01586_),
    .B(_01621_),
    .Y(_01622_));
 sky130_fd_sc_hd__xnor2_1 _20446_ (.A(_01586_),
    .B(_01621_),
    .Y(_01623_));
 sky130_fd_sc_hd__a21oi_2 _20447_ (.A1(_01471_),
    .A2(_01473_),
    .B1(_01623_),
    .Y(_01624_));
 sky130_fd_sc_hd__inv_2 _20448_ (.A(_01624_),
    .Y(_01625_));
 sky130_fd_sc_hd__and3_1 _20449_ (.A(_01471_),
    .B(_01473_),
    .C(_01623_),
    .X(_01626_));
 sky130_fd_sc_hd__or3_4 _20450_ (.A(_01585_),
    .B(_01624_),
    .C(_01626_),
    .X(_01627_));
 sky130_fd_sc_hd__o21ai_2 _20451_ (.A1(_01624_),
    .A2(_01626_),
    .B1(_01585_),
    .Y(_01628_));
 sky130_fd_sc_hd__o211a_2 _20452_ (.A1(_01440_),
    .A2(_01480_),
    .B1(_01627_),
    .C1(_01628_),
    .X(_01629_));
 sky130_fd_sc_hd__a211oi_4 _20453_ (.A1(_01627_),
    .A2(_01628_),
    .B1(_01440_),
    .C1(_01480_),
    .Y(_01630_));
 sky130_fd_sc_hd__a22o_1 _20454_ (.A1(net255),
    .A2(net72),
    .B1(net69),
    .B2(net261),
    .X(_01631_));
 sky130_fd_sc_hd__and4_1 _20455_ (.A(net255),
    .B(net261),
    .C(net72),
    .D(net69),
    .X(_01632_));
 sky130_fd_sc_hd__inv_2 _20456_ (.A(_01632_),
    .Y(_01633_));
 sky130_fd_sc_hd__a22oi_1 _20457_ (.A1(net265),
    .A2(net66),
    .B1(_01631_),
    .B2(_01633_),
    .Y(_01634_));
 sky130_fd_sc_hd__and4_1 _20458_ (.A(net265),
    .B(net66),
    .C(_01631_),
    .D(_01633_),
    .X(_01635_));
 sky130_fd_sc_hd__or2_2 _20459_ (.A(_01634_),
    .B(_01635_),
    .X(_01636_));
 sky130_fd_sc_hd__nor2_2 _20460_ (.A(_01487_),
    .B(_01490_),
    .Y(_01637_));
 sky130_fd_sc_hd__xnor2_2 _20461_ (.A(_01636_),
    .B(_01637_),
    .Y(_01638_));
 sky130_fd_sc_hd__and4b_2 _20462_ (.A_N(net277),
    .B(net63),
    .C(net62),
    .D(net269),
    .X(_01639_));
 sky130_fd_sc_hd__o2bb2a_1 _20463_ (.A1_N(net269),
    .A2_N(net63),
    .B1(net56),
    .B2(net277),
    .X(_01640_));
 sky130_fd_sc_hd__nor2_1 _20464_ (.A(_01639_),
    .B(_01640_),
    .Y(_01641_));
 sky130_fd_sc_hd__xnor2_1 _20465_ (.A(_01638_),
    .B(_01641_),
    .Y(_01642_));
 sky130_fd_sc_hd__nor3_1 _20466_ (.A(_01493_),
    .B(_01499_),
    .C(_01642_),
    .Y(_01643_));
 sky130_fd_sc_hd__o21a_1 _20467_ (.A1(_01493_),
    .A2(_01499_),
    .B1(_01642_),
    .X(_01644_));
 sky130_fd_sc_hd__or2_1 _20468_ (.A(_01643_),
    .B(_01644_),
    .X(_01645_));
 sky130_fd_sc_hd__nor2_1 _20469_ (.A(_01496_),
    .B(_01645_),
    .Y(_01646_));
 sky130_fd_sc_hd__and2_1 _20470_ (.A(_01496_),
    .B(_01645_),
    .X(_01647_));
 sky130_fd_sc_hd__or2_1 _20471_ (.A(_01646_),
    .B(_01647_),
    .X(_01648_));
 sky130_fd_sc_hd__or2_1 _20472_ (.A(_01511_),
    .B(_01513_),
    .X(_01649_));
 sky130_fd_sc_hd__nand2_1 _20473_ (.A(_01443_),
    .B(_01445_),
    .Y(_01650_));
 sky130_fd_sc_hd__a22o_1 _20474_ (.A1(net245),
    .A2(net83),
    .B1(net79),
    .B2(net628),
    .X(_01651_));
 sky130_fd_sc_hd__inv_2 _20475_ (.A(_01651_),
    .Y(_01652_));
 sky130_fd_sc_hd__and4_1 _20476_ (.A(net246),
    .B(net628),
    .C(net83),
    .D(net79),
    .X(_01653_));
 sky130_fd_sc_hd__o2bb2a_1 _20477_ (.A1_N(net251),
    .A2_N(net77),
    .B1(_01652_),
    .B2(_01653_),
    .X(_01654_));
 sky130_fd_sc_hd__and4b_1 _20478_ (.A_N(_01653_),
    .B(net76),
    .C(net251),
    .D(_01651_),
    .X(_01655_));
 sky130_fd_sc_hd__or2_1 _20479_ (.A(_01654_),
    .B(_01655_),
    .X(_01656_));
 sky130_fd_sc_hd__nand2b_1 _20480_ (.A_N(_01656_),
    .B(_01650_),
    .Y(_01657_));
 sky130_fd_sc_hd__xnor2_1 _20481_ (.A(_01650_),
    .B(_01656_),
    .Y(_01658_));
 sky130_fd_sc_hd__nand2_1 _20482_ (.A(_01649_),
    .B(_01658_),
    .Y(_01659_));
 sky130_fd_sc_hd__or2_1 _20483_ (.A(_01649_),
    .B(_01658_),
    .X(_01660_));
 sky130_fd_sc_hd__nand2_1 _20484_ (.A(_01659_),
    .B(_01660_),
    .Y(_01661_));
 sky130_fd_sc_hd__a21oi_4 _20485_ (.A1(_01454_),
    .A2(_01456_),
    .B1(_01661_),
    .Y(_01662_));
 sky130_fd_sc_hd__and3_1 _20486_ (.A(_01454_),
    .B(_01456_),
    .C(_01661_),
    .X(_01663_));
 sky130_fd_sc_hd__a211oi_4 _20487_ (.A1(_01515_),
    .A2(_01517_),
    .B1(_01662_),
    .C1(_01663_),
    .Y(_01664_));
 sky130_fd_sc_hd__o211a_1 _20488_ (.A1(_01662_),
    .A2(_01663_),
    .B1(_01515_),
    .C1(_01517_),
    .X(_01665_));
 sky130_fd_sc_hd__a211oi_4 _20489_ (.A1(_01520_),
    .A2(_01522_),
    .B1(_01664_),
    .C1(_01665_),
    .Y(_01666_));
 sky130_fd_sc_hd__o211a_1 _20490_ (.A1(_01664_),
    .A2(_01665_),
    .B1(_01520_),
    .C1(_01522_),
    .X(_01667_));
 sky130_fd_sc_hd__or3_2 _20491_ (.A(_01648_),
    .B(_01666_),
    .C(_01667_),
    .X(_01668_));
 sky130_fd_sc_hd__inv_2 _20492_ (.A(_01668_),
    .Y(_01669_));
 sky130_fd_sc_hd__o21ai_1 _20493_ (.A1(_01666_),
    .A2(_01667_),
    .B1(_01648_),
    .Y(_01670_));
 sky130_fd_sc_hd__o211a_1 _20494_ (.A1(_01475_),
    .A2(_01478_),
    .B1(_01668_),
    .C1(_01670_),
    .X(_01671_));
 sky130_fd_sc_hd__a211oi_1 _20495_ (.A1(_01668_),
    .A2(_01670_),
    .B1(_01475_),
    .C1(_01478_),
    .Y(_01672_));
 sky130_fd_sc_hd__nor2_1 _20496_ (.A(_01671_),
    .B(_01672_),
    .Y(_01673_));
 sky130_fd_sc_hd__o21a_2 _20497_ (.A1(_01524_),
    .A2(_01526_),
    .B1(_01673_),
    .X(_01674_));
 sky130_fd_sc_hd__nor3_2 _20498_ (.A(_01524_),
    .B(_01526_),
    .C(_01673_),
    .Y(_01675_));
 sky130_fd_sc_hd__nor4_4 _20499_ (.A(_01629_),
    .B(_01630_),
    .C(_01674_),
    .D(_01675_),
    .Y(_01676_));
 sky130_fd_sc_hd__o22a_1 _20500_ (.A1(_01629_),
    .A2(_01630_),
    .B1(_01674_),
    .B2(_01675_),
    .X(_01677_));
 sky130_fd_sc_hd__a211oi_4 _20501_ (.A1(_01482_),
    .A2(_01533_),
    .B1(_01676_),
    .C1(_01677_),
    .Y(_01678_));
 sky130_fd_sc_hd__o211a_1 _20502_ (.A1(_01676_),
    .A2(_01677_),
    .B1(_01482_),
    .C1(_01533_),
    .X(_01679_));
 sky130_fd_sc_hd__a211oi_4 _20503_ (.A1(_01529_),
    .A2(_01531_),
    .B1(_01678_),
    .C1(_01679_),
    .Y(_01680_));
 sky130_fd_sc_hd__o211a_1 _20504_ (.A1(_01678_),
    .A2(_01679_),
    .B1(_01529_),
    .C1(_01531_),
    .X(_01681_));
 sky130_fd_sc_hd__a211oi_2 _20505_ (.A1(_01535_),
    .A2(_01537_),
    .B1(_01680_),
    .C1(_01681_),
    .Y(_01682_));
 sky130_fd_sc_hd__o211a_1 _20506_ (.A1(_01680_),
    .A2(_01681_),
    .B1(_01535_),
    .C1(_01537_),
    .X(_01683_));
 sky130_fd_sc_hd__a211oi_2 _20507_ (.A1(_01502_),
    .A2(_01505_),
    .B1(_01682_),
    .C1(_01683_),
    .Y(_01684_));
 sky130_fd_sc_hd__o211a_1 _20508_ (.A1(_01682_),
    .A2(_01683_),
    .B1(_01502_),
    .C1(_01505_),
    .X(_01685_));
 sky130_fd_sc_hd__a211oi_1 _20509_ (.A1(_01539_),
    .A2(_01543_),
    .B1(_01684_),
    .C1(_01685_),
    .Y(_01686_));
 sky130_fd_sc_hd__o211ai_1 _20510_ (.A1(_01684_),
    .A2(_01685_),
    .B1(_01539_),
    .C1(_01543_),
    .Y(_01687_));
 sky130_fd_sc_hd__and2b_2 _20511_ (.A_N(_01686_),
    .B(_01687_),
    .X(_01688_));
 sky130_fd_sc_hd__inv_2 _20512_ (.A(_01688_),
    .Y(_01689_));
 sky130_fd_sc_hd__nor2_1 _20513_ (.A(_01547_),
    .B(_01553_),
    .Y(_01690_));
 sky130_fd_sc_hd__xnor2_2 _20514_ (.A(_01688_),
    .B(_01690_),
    .Y(_01691_));
 sky130_fd_sc_hd__a22o_1 _20515_ (.A1(net831),
    .A2(net7),
    .B1(_07105_),
    .B2(_03052_),
    .X(_01692_));
 sky130_fd_sc_hd__a21o_1 _20516_ (.A1(net10),
    .A2(_01691_),
    .B1(_01692_),
    .X(_01693_));
 sky130_fd_sc_hd__mux2_1 _20517_ (.A0(net919),
    .A1(_01693_),
    .S(net1),
    .X(_00323_));
 sky130_fd_sc_hd__a32o_1 _20518_ (.A1(_01566_),
    .A2(_01567_),
    .A3(_01575_),
    .B1(_01574_),
    .B2(_01569_),
    .X(_01694_));
 sky130_fd_sc_hd__a22o_1 _20519_ (.A1(net132),
    .A2(net198),
    .B1(net196),
    .B2(net137),
    .X(_01695_));
 sky130_fd_sc_hd__and4_1 _20520_ (.A(net137),
    .B(net132),
    .C(net198),
    .D(net196),
    .X(_01696_));
 sky130_fd_sc_hd__inv_2 _20521_ (.A(_01696_),
    .Y(_01697_));
 sky130_fd_sc_hd__a22oi_1 _20522_ (.A1(net128),
    .A2(net201),
    .B1(_01695_),
    .B2(_01697_),
    .Y(_01698_));
 sky130_fd_sc_hd__and4_1 _20523_ (.A(net128),
    .B(net201),
    .C(_01695_),
    .D(_01697_),
    .X(_01699_));
 sky130_fd_sc_hd__or2_1 _20524_ (.A(_01698_),
    .B(_01699_),
    .X(_01700_));
 sky130_fd_sc_hd__a21oi_1 _20525_ (.A1(net142),
    .A2(net194),
    .B1(_01572_),
    .Y(_01701_));
 sky130_fd_sc_hd__a21o_1 _20526_ (.A1(_01570_),
    .A2(_01572_),
    .B1(_01571_),
    .X(_01702_));
 sky130_fd_sc_hd__a21oi_1 _20527_ (.A1(net142),
    .A2(_01702_),
    .B1(_01701_),
    .Y(_01703_));
 sky130_fd_sc_hd__or3b_1 _20528_ (.A(_01698_),
    .B(_01699_),
    .C_N(_01703_),
    .X(_01704_));
 sky130_fd_sc_hd__xnor2_1 _20529_ (.A(_01700_),
    .B(_01703_),
    .Y(_01705_));
 sky130_fd_sc_hd__nand2_1 _20530_ (.A(_01563_),
    .B(_01705_),
    .Y(_01706_));
 sky130_fd_sc_hd__xnor2_1 _20531_ (.A(_01562_),
    .B(_01705_),
    .Y(_01707_));
 sky130_fd_sc_hd__nand2_1 _20532_ (.A(_01694_),
    .B(_01707_),
    .Y(_01708_));
 sky130_fd_sc_hd__xnor2_1 _20533_ (.A(_01694_),
    .B(_01707_),
    .Y(_01709_));
 sky130_fd_sc_hd__and2_1 _20534_ (.A(_01560_),
    .B(_01709_),
    .X(_01710_));
 sky130_fd_sc_hd__nor2_1 _20535_ (.A(_01560_),
    .B(_01709_),
    .Y(_01711_));
 sky130_fd_sc_hd__nor2_1 _20536_ (.A(_01710_),
    .B(_01711_),
    .Y(_01712_));
 sky130_fd_sc_hd__o21bai_1 _20537_ (.A1(_01560_),
    .A2(_01580_),
    .B1_N(_01557_),
    .Y(_01713_));
 sky130_fd_sc_hd__nor2_1 _20538_ (.A(_01712_),
    .B(_01713_),
    .Y(_01714_));
 sky130_fd_sc_hd__and2_1 _20539_ (.A(_01712_),
    .B(_01713_),
    .X(_01715_));
 sky130_fd_sc_hd__or2_1 _20540_ (.A(_01714_),
    .B(_01715_),
    .X(_01716_));
 sky130_fd_sc_hd__a22o_1 _20541_ (.A1(net226),
    .A2(net97),
    .B1(net91),
    .B2(net230),
    .X(_01717_));
 sky130_fd_sc_hd__nand4_1 _20542_ (.A(net230),
    .B(net226),
    .C(net97),
    .D(net91),
    .Y(_01718_));
 sky130_fd_sc_hd__a22o_1 _20543_ (.A1(net237),
    .A2(net86),
    .B1(_01717_),
    .B2(_01718_),
    .X(_01719_));
 sky130_fd_sc_hd__nand4_1 _20544_ (.A(net236),
    .B(net86),
    .C(_01717_),
    .D(_01718_),
    .Y(_01720_));
 sky130_fd_sc_hd__nand2_1 _20545_ (.A(_01719_),
    .B(_01720_),
    .Y(_01721_));
 sky130_fd_sc_hd__a22o_1 _20546_ (.A1(net102),
    .A2(net217),
    .B1(net213),
    .B2(net107),
    .X(_01722_));
 sky130_fd_sc_hd__and4_1 _20547_ (.A(net107),
    .B(net102),
    .C(net217),
    .D(net213),
    .X(_01723_));
 sky130_fd_sc_hd__inv_2 _20548_ (.A(_01723_),
    .Y(_01724_));
 sky130_fd_sc_hd__a22oi_1 _20549_ (.A1(net98),
    .A2(net222),
    .B1(_01722_),
    .B2(_01724_),
    .Y(_01725_));
 sky130_fd_sc_hd__and4_1 _20550_ (.A(net98),
    .B(net222),
    .C(_01722_),
    .D(_01724_),
    .X(_01726_));
 sky130_fd_sc_hd__or2_1 _20551_ (.A(_01725_),
    .B(_01726_),
    .X(_01727_));
 sky130_fd_sc_hd__or2_1 _20552_ (.A(_01593_),
    .B(_01596_),
    .X(_01728_));
 sky130_fd_sc_hd__nand2b_1 _20553_ (.A_N(_01727_),
    .B(_01728_),
    .Y(_01729_));
 sky130_fd_sc_hd__xor2_1 _20554_ (.A(_01727_),
    .B(_01728_),
    .X(_01730_));
 sky130_fd_sc_hd__or2_1 _20555_ (.A(_01721_),
    .B(_01730_),
    .X(_01731_));
 sky130_fd_sc_hd__nand2_1 _20556_ (.A(_01721_),
    .B(_01730_),
    .Y(_01732_));
 sky130_fd_sc_hd__and2_1 _20557_ (.A(_01731_),
    .B(_01732_),
    .X(_01733_));
 sky130_fd_sc_hd__or2_1 _20558_ (.A(_01608_),
    .B(_01610_),
    .X(_01734_));
 sky130_fd_sc_hd__nand2_1 _20559_ (.A(_01565_),
    .B(_01567_),
    .Y(_01735_));
 sky130_fd_sc_hd__a22o_1 _20560_ (.A1(net118),
    .A2(net207),
    .B1(net204),
    .B2(net123),
    .X(_01736_));
 sky130_fd_sc_hd__inv_2 _20561_ (.A(_01736_),
    .Y(_01737_));
 sky130_fd_sc_hd__and4_1 _20562_ (.A(net123),
    .B(net121),
    .C(net207),
    .D(net204),
    .X(_01738_));
 sky130_fd_sc_hd__o2bb2a_1 _20563_ (.A1_N(net113),
    .A2_N(net210),
    .B1(_01737_),
    .B2(_01738_),
    .X(_01739_));
 sky130_fd_sc_hd__and4b_1 _20564_ (.A_N(_01738_),
    .B(net210),
    .C(net113),
    .D(_01736_),
    .X(_01740_));
 sky130_fd_sc_hd__or2_1 _20565_ (.A(_01739_),
    .B(_01740_),
    .X(_01741_));
 sky130_fd_sc_hd__nand2b_1 _20566_ (.A_N(_01741_),
    .B(_01735_),
    .Y(_01742_));
 sky130_fd_sc_hd__xnor2_1 _20567_ (.A(_01735_),
    .B(_01741_),
    .Y(_01743_));
 sky130_fd_sc_hd__nand2_1 _20568_ (.A(_01734_),
    .B(_01743_),
    .Y(_01744_));
 sky130_fd_sc_hd__xnor2_1 _20569_ (.A(_01734_),
    .B(_01743_),
    .Y(_01745_));
 sky130_fd_sc_hd__a21o_1 _20570_ (.A1(_01612_),
    .A2(_01614_),
    .B1(_01745_),
    .X(_01746_));
 sky130_fd_sc_hd__nand3_1 _20571_ (.A(_01612_),
    .B(_01614_),
    .C(_01745_),
    .Y(_01747_));
 sky130_fd_sc_hd__nand3_2 _20572_ (.A(_01733_),
    .B(_01746_),
    .C(_01747_),
    .Y(_01748_));
 sky130_fd_sc_hd__a21o_1 _20573_ (.A1(_01746_),
    .A2(_01747_),
    .B1(_01733_),
    .X(_01749_));
 sky130_fd_sc_hd__o211a_2 _20574_ (.A1(_01577_),
    .A2(_01579_),
    .B1(_01748_),
    .C1(_01749_),
    .X(_01750_));
 sky130_fd_sc_hd__a211oi_2 _20575_ (.A1(_01748_),
    .A2(_01749_),
    .B1(_01577_),
    .C1(_01579_),
    .Y(_01751_));
 sky130_fd_sc_hd__a211oi_4 _20576_ (.A1(_01616_),
    .A2(_01619_),
    .B1(_01750_),
    .C1(_01751_),
    .Y(_01752_));
 sky130_fd_sc_hd__o211a_1 _20577_ (.A1(_01750_),
    .A2(_01751_),
    .B1(_01616_),
    .C1(_01619_),
    .X(_01753_));
 sky130_fd_sc_hd__nor3_4 _20578_ (.A(_01716_),
    .B(_01752_),
    .C(_01753_),
    .Y(_01754_));
 sky130_fd_sc_hd__o21a_1 _20579_ (.A1(_01752_),
    .A2(_01753_),
    .B1(_01716_),
    .X(_01755_));
 sky130_fd_sc_hd__a211oi_4 _20580_ (.A1(_01584_),
    .A2(_01627_),
    .B1(_01754_),
    .C1(_01755_),
    .Y(_01756_));
 sky130_fd_sc_hd__o211a_1 _20581_ (.A1(_01754_),
    .A2(_01755_),
    .B1(_01584_),
    .C1(_01627_),
    .X(_01757_));
 sky130_fd_sc_hd__a22o_1 _20582_ (.A1(net250),
    .A2(net72),
    .B1(net69),
    .B2(net255),
    .X(_01758_));
 sky130_fd_sc_hd__and4_1 _20583_ (.A(net251),
    .B(net255),
    .C(net72),
    .D(net69),
    .X(_01759_));
 sky130_fd_sc_hd__inv_2 _20584_ (.A(_01759_),
    .Y(_01760_));
 sky130_fd_sc_hd__a22oi_1 _20585_ (.A1(net261),
    .A2(net66),
    .B1(_01758_),
    .B2(_01760_),
    .Y(_01761_));
 sky130_fd_sc_hd__and4_1 _20586_ (.A(net261),
    .B(net66),
    .C(_01758_),
    .D(_01760_),
    .X(_01762_));
 sky130_fd_sc_hd__or2_2 _20587_ (.A(_01761_),
    .B(_01762_),
    .X(_01763_));
 sky130_fd_sc_hd__nor2_2 _20588_ (.A(_01632_),
    .B(_01635_),
    .Y(_01764_));
 sky130_fd_sc_hd__xnor2_2 _20589_ (.A(_01763_),
    .B(_01764_),
    .Y(_01765_));
 sky130_fd_sc_hd__and4b_2 _20590_ (.A_N(net269),
    .B(net63),
    .C(net62),
    .D(net265),
    .X(_01766_));
 sky130_fd_sc_hd__inv_2 _20591_ (.A(_01766_),
    .Y(_01767_));
 sky130_fd_sc_hd__o2bb2a_1 _20592_ (.A1_N(net265),
    .A2_N(net63),
    .B1(net56),
    .B2(net269),
    .X(_01768_));
 sky130_fd_sc_hd__nor2_1 _20593_ (.A(_01766_),
    .B(_01768_),
    .Y(_01769_));
 sky130_fd_sc_hd__xnor2_1 _20594_ (.A(_01765_),
    .B(_01769_),
    .Y(_01770_));
 sky130_fd_sc_hd__o32ai_4 _20595_ (.A1(_01638_),
    .A2(_01639_),
    .A3(_01640_),
    .B1(_01637_),
    .B2(_01636_),
    .Y(_01771_));
 sky130_fd_sc_hd__nand2_1 _20596_ (.A(_01770_),
    .B(_01771_),
    .Y(_01772_));
 sky130_fd_sc_hd__xnor2_1 _20597_ (.A(_01770_),
    .B(_01771_),
    .Y(_01773_));
 sky130_fd_sc_hd__inv_2 _20598_ (.A(_01773_),
    .Y(_01774_));
 sky130_fd_sc_hd__nand2_1 _20599_ (.A(_01639_),
    .B(_01774_),
    .Y(_01775_));
 sky130_fd_sc_hd__or2_1 _20600_ (.A(_01639_),
    .B(_01774_),
    .X(_01776_));
 sky130_fd_sc_hd__nand2_1 _20601_ (.A(_01775_),
    .B(_01776_),
    .Y(_01777_));
 sky130_fd_sc_hd__or2_1 _20602_ (.A(_01653_),
    .B(_01655_),
    .X(_01778_));
 sky130_fd_sc_hd__nand2_1 _20603_ (.A(_01588_),
    .B(_01590_),
    .Y(_01779_));
 sky130_fd_sc_hd__a22o_1 _20604_ (.A1(net241),
    .A2(net83),
    .B1(net79),
    .B2(net246),
    .X(_01780_));
 sky130_fd_sc_hd__inv_2 _20605_ (.A(_01780_),
    .Y(_01781_));
 sky130_fd_sc_hd__and4_1 _20606_ (.A(net246),
    .B(net241),
    .C(net83),
    .D(net80),
    .X(_01782_));
 sky130_fd_sc_hd__o2bb2a_1 _20607_ (.A1_N(net629),
    .A2_N(net76),
    .B1(_01781_),
    .B2(_01782_),
    .X(_01783_));
 sky130_fd_sc_hd__and4b_1 _20608_ (.A_N(_01782_),
    .B(net76),
    .C(net629),
    .D(_01780_),
    .X(_01784_));
 sky130_fd_sc_hd__or2_1 _20609_ (.A(_01783_),
    .B(_01784_),
    .X(_01785_));
 sky130_fd_sc_hd__nand2b_1 _20610_ (.A_N(_01785_),
    .B(_01779_),
    .Y(_01786_));
 sky130_fd_sc_hd__xnor2_1 _20611_ (.A(_01779_),
    .B(_01785_),
    .Y(_01787_));
 sky130_fd_sc_hd__nand2_1 _20612_ (.A(_01778_),
    .B(_01787_),
    .Y(_01788_));
 sky130_fd_sc_hd__xnor2_1 _20613_ (.A(_01778_),
    .B(_01787_),
    .Y(_01789_));
 sky130_fd_sc_hd__a21oi_1 _20614_ (.A1(_01599_),
    .A2(_01601_),
    .B1(_01789_),
    .Y(_01790_));
 sky130_fd_sc_hd__a21o_1 _20615_ (.A1(_01599_),
    .A2(_01601_),
    .B1(_01789_),
    .X(_01791_));
 sky130_fd_sc_hd__and3_1 _20616_ (.A(_01599_),
    .B(_01601_),
    .C(_01789_),
    .X(_01792_));
 sky130_fd_sc_hd__a211o_1 _20617_ (.A1(_01657_),
    .A2(_01659_),
    .B1(_01790_),
    .C1(_01792_),
    .X(_01793_));
 sky130_fd_sc_hd__o211ai_2 _20618_ (.A1(_01790_),
    .A2(_01792_),
    .B1(_01657_),
    .C1(_01659_),
    .Y(_01794_));
 sky130_fd_sc_hd__o211a_1 _20619_ (.A1(_01662_),
    .A2(_01664_),
    .B1(_01793_),
    .C1(_01794_),
    .X(_01795_));
 sky130_fd_sc_hd__a211oi_2 _20620_ (.A1(_01793_),
    .A2(_01794_),
    .B1(_01662_),
    .C1(_01664_),
    .Y(_01796_));
 sky130_fd_sc_hd__nor3_2 _20621_ (.A(_01777_),
    .B(_01795_),
    .C(_01796_),
    .Y(_01797_));
 sky130_fd_sc_hd__o21a_1 _20622_ (.A1(_01795_),
    .A2(_01796_),
    .B1(_01777_),
    .X(_01798_));
 sky130_fd_sc_hd__a211o_2 _20623_ (.A1(_01622_),
    .A2(_01625_),
    .B1(_01797_),
    .C1(_01798_),
    .X(_01799_));
 sky130_fd_sc_hd__o211ai_4 _20624_ (.A1(_01797_),
    .A2(_01798_),
    .B1(_01622_),
    .C1(_01625_),
    .Y(_01800_));
 sky130_fd_sc_hd__o211ai_4 _20625_ (.A1(_01666_),
    .A2(_01669_),
    .B1(_01799_),
    .C1(_01800_),
    .Y(_01801_));
 sky130_fd_sc_hd__a211o_1 _20626_ (.A1(_01799_),
    .A2(_01800_),
    .B1(_01666_),
    .C1(_01669_),
    .X(_01802_));
 sky130_fd_sc_hd__and4bb_1 _20627_ (.A_N(_01756_),
    .B_N(_01757_),
    .C(_01801_),
    .D(_01802_),
    .X(_01803_));
 sky130_fd_sc_hd__or4bb_2 _20628_ (.A(_01756_),
    .B(_01757_),
    .C_N(_01801_),
    .D_N(_01802_),
    .X(_01804_));
 sky130_fd_sc_hd__a2bb2o_1 _20629_ (.A1_N(_01756_),
    .A2_N(_01757_),
    .B1(_01801_),
    .B2(_01802_),
    .X(_01805_));
 sky130_fd_sc_hd__o211ai_4 _20630_ (.A1(_01629_),
    .A2(_01676_),
    .B1(_01804_),
    .C1(_01805_),
    .Y(_01806_));
 sky130_fd_sc_hd__a211o_1 _20631_ (.A1(_01804_),
    .A2(_01805_),
    .B1(_01629_),
    .C1(_01676_),
    .X(_01807_));
 sky130_fd_sc_hd__o211ai_4 _20632_ (.A1(_01671_),
    .A2(_01674_),
    .B1(_01806_),
    .C1(_01807_),
    .Y(_01808_));
 sky130_fd_sc_hd__a211o_1 _20633_ (.A1(_01806_),
    .A2(_01807_),
    .B1(_01671_),
    .C1(_01674_),
    .X(_01809_));
 sky130_fd_sc_hd__o211ai_4 _20634_ (.A1(_01678_),
    .A2(_01680_),
    .B1(_01808_),
    .C1(_01809_),
    .Y(_01810_));
 sky130_fd_sc_hd__a211o_1 _20635_ (.A1(_01808_),
    .A2(_01809_),
    .B1(_01678_),
    .C1(_01680_),
    .X(_01811_));
 sky130_fd_sc_hd__o211ai_2 _20636_ (.A1(_01644_),
    .A2(_01646_),
    .B1(_01810_),
    .C1(_01811_),
    .Y(_01812_));
 sky130_fd_sc_hd__a211o_1 _20637_ (.A1(_01810_),
    .A2(_01811_),
    .B1(_01644_),
    .C1(_01646_),
    .X(_01813_));
 sky130_fd_sc_hd__nand2_1 _20638_ (.A(_01812_),
    .B(_01813_),
    .Y(_01814_));
 sky130_fd_sc_hd__or2_2 _20639_ (.A(_01682_),
    .B(_01684_),
    .X(_01815_));
 sky130_fd_sc_hd__and2b_1 _20640_ (.A_N(_01814_),
    .B(_01815_),
    .X(_01816_));
 sky130_fd_sc_hd__xnor2_2 _20641_ (.A(_01814_),
    .B(_01815_),
    .Y(_01817_));
 sky130_fd_sc_hd__o21ai_1 _20642_ (.A1(_01547_),
    .A2(_01686_),
    .B1(_01687_),
    .Y(_01818_));
 sky130_fd_sc_hd__nand2_1 _20643_ (.A(_01549_),
    .B(_01688_),
    .Y(_01819_));
 sky130_fd_sc_hd__o21ai_2 _20644_ (.A1(_01552_),
    .A2(_01819_),
    .B1(_01818_),
    .Y(_01820_));
 sky130_fd_sc_hd__xor2_2 _20645_ (.A(_01817_),
    .B(_01820_),
    .X(_01821_));
 sky130_fd_sc_hd__nor2_1 _20646_ (.A(net43),
    .B(_07236_),
    .Y(_01822_));
 sky130_fd_sc_hd__a221o_1 _20647_ (.A1(net758),
    .A2(net8),
    .B1(_01821_),
    .B2(_03050_),
    .C1(_01822_),
    .X(_01823_));
 sky130_fd_sc_hd__mux2_1 _20648_ (.A0(net922),
    .A1(_01823_),
    .S(net2),
    .X(_00324_));
 sky130_fd_sc_hd__and2_1 _20649_ (.A(net143),
    .B(_01571_),
    .X(_01824_));
 sky130_fd_sc_hd__nand2_2 _20650_ (.A(net143),
    .B(_01571_),
    .Y(_01825_));
 sky130_fd_sc_hd__nand2_1 _20651_ (.A(_01704_),
    .B(_01825_),
    .Y(_01826_));
 sky130_fd_sc_hd__a22oi_1 _20652_ (.A1(net132),
    .A2(\mul1.a[30] ),
    .B1(net194),
    .B2(net137),
    .Y(_01827_));
 sky130_fd_sc_hd__and4_1 _20653_ (.A(net137),
    .B(net132),
    .C(\mul1.a[30] ),
    .D(net194),
    .X(_01828_));
 sky130_fd_sc_hd__nor2_1 _20654_ (.A(_01827_),
    .B(_01828_),
    .Y(_01829_));
 sky130_fd_sc_hd__nand2_1 _20655_ (.A(net128),
    .B(net198),
    .Y(_01830_));
 sky130_fd_sc_hd__xor2_1 _20656_ (.A(_01829_),
    .B(_01830_),
    .X(_01831_));
 sky130_fd_sc_hd__or2_4 _20657_ (.A(_01701_),
    .B(_01824_),
    .X(_01832_));
 sky130_fd_sc_hd__xor2_1 _20658_ (.A(_01831_),
    .B(_01832_),
    .X(_01833_));
 sky130_fd_sc_hd__nand2_1 _20659_ (.A(_01563_),
    .B(_01833_),
    .Y(_01834_));
 sky130_fd_sc_hd__xnor2_1 _20660_ (.A(_01563_),
    .B(_01833_),
    .Y(_01835_));
 sky130_fd_sc_hd__nand2b_1 _20661_ (.A_N(_01835_),
    .B(_01826_),
    .Y(_01836_));
 sky130_fd_sc_hd__xor2_1 _20662_ (.A(_01826_),
    .B(_01835_),
    .X(_01837_));
 sky130_fd_sc_hd__nor2_1 _20663_ (.A(_01560_),
    .B(_01837_),
    .Y(_01838_));
 sky130_fd_sc_hd__xnor2_1 _20664_ (.A(_01559_),
    .B(_01837_),
    .Y(_01839_));
 sky130_fd_sc_hd__or3_1 _20665_ (.A(_01557_),
    .B(_01711_),
    .C(_01839_),
    .X(_01840_));
 sky130_fd_sc_hd__o21ai_2 _20666_ (.A1(_01557_),
    .A2(_01711_),
    .B1(_01839_),
    .Y(_01841_));
 sky130_fd_sc_hd__nand2_1 _20667_ (.A(_01840_),
    .B(_01841_),
    .Y(_01842_));
 sky130_fd_sc_hd__a22o_1 _20668_ (.A1(net97),
    .A2(net222),
    .B1(net91),
    .B2(net226),
    .X(_01843_));
 sky130_fd_sc_hd__nand4_2 _20669_ (.A(net226),
    .B(net97),
    .C(net222),
    .D(net91),
    .Y(_01844_));
 sky130_fd_sc_hd__a22o_1 _20670_ (.A1(net230),
    .A2(net86),
    .B1(_01843_),
    .B2(_01844_),
    .X(_01845_));
 sky130_fd_sc_hd__nand4_1 _20671_ (.A(net230),
    .B(net87),
    .C(_01843_),
    .D(_01844_),
    .Y(_01846_));
 sky130_fd_sc_hd__nand2_1 _20672_ (.A(_01845_),
    .B(_01846_),
    .Y(_01847_));
 sky130_fd_sc_hd__a22o_1 _20673_ (.A1(net102),
    .A2(net213),
    .B1(net210),
    .B2(net107),
    .X(_01848_));
 sky130_fd_sc_hd__and4_1 _20674_ (.A(net107),
    .B(net102),
    .C(net213),
    .D(net210),
    .X(_01849_));
 sky130_fd_sc_hd__inv_2 _20675_ (.A(_01849_),
    .Y(_01850_));
 sky130_fd_sc_hd__a22oi_1 _20676_ (.A1(net98),
    .A2(net218),
    .B1(_01848_),
    .B2(_01850_),
    .Y(_01851_));
 sky130_fd_sc_hd__and4_1 _20677_ (.A(net98),
    .B(net218),
    .C(_01848_),
    .D(_01850_),
    .X(_01852_));
 sky130_fd_sc_hd__or2_1 _20678_ (.A(_01851_),
    .B(_01852_),
    .X(_01853_));
 sky130_fd_sc_hd__or2_1 _20679_ (.A(_01723_),
    .B(_01726_),
    .X(_01854_));
 sky130_fd_sc_hd__nand2b_1 _20680_ (.A_N(_01853_),
    .B(_01854_),
    .Y(_01855_));
 sky130_fd_sc_hd__xor2_1 _20681_ (.A(_01853_),
    .B(_01854_),
    .X(_01856_));
 sky130_fd_sc_hd__or2_1 _20682_ (.A(_01847_),
    .B(_01856_),
    .X(_01857_));
 sky130_fd_sc_hd__nand2_1 _20683_ (.A(_01847_),
    .B(_01856_),
    .Y(_01858_));
 sky130_fd_sc_hd__and2_1 _20684_ (.A(_01857_),
    .B(_01858_),
    .X(_01859_));
 sky130_fd_sc_hd__or2_1 _20685_ (.A(_01738_),
    .B(_01740_),
    .X(_01860_));
 sky130_fd_sc_hd__nor2_1 _20686_ (.A(_01696_),
    .B(_01699_),
    .Y(_01861_));
 sky130_fd_sc_hd__a22o_1 _20687_ (.A1(net118),
    .A2(net204),
    .B1(net201),
    .B2(net123),
    .X(_01862_));
 sky130_fd_sc_hd__inv_2 _20688_ (.A(_01862_),
    .Y(_01863_));
 sky130_fd_sc_hd__and4_1 _20689_ (.A(net126),
    .B(net118),
    .C(net204),
    .D(net201),
    .X(_01864_));
 sky130_fd_sc_hd__o2bb2a_1 _20690_ (.A1_N(net113),
    .A2_N(net207),
    .B1(_01863_),
    .B2(_01864_),
    .X(_01865_));
 sky130_fd_sc_hd__and4b_1 _20691_ (.A_N(_01864_),
    .B(net207),
    .C(net113),
    .D(_01862_),
    .X(_01866_));
 sky130_fd_sc_hd__or2_1 _20692_ (.A(_01865_),
    .B(_01866_),
    .X(_01867_));
 sky130_fd_sc_hd__or2_1 _20693_ (.A(_01861_),
    .B(_01867_),
    .X(_01868_));
 sky130_fd_sc_hd__xor2_1 _20694_ (.A(_01861_),
    .B(_01867_),
    .X(_01869_));
 sky130_fd_sc_hd__nand2_1 _20695_ (.A(_01860_),
    .B(_01869_),
    .Y(_01870_));
 sky130_fd_sc_hd__xnor2_1 _20696_ (.A(_01860_),
    .B(_01869_),
    .Y(_01871_));
 sky130_fd_sc_hd__a21o_1 _20697_ (.A1(_01742_),
    .A2(_01744_),
    .B1(_01871_),
    .X(_01872_));
 sky130_fd_sc_hd__nand3_1 _20698_ (.A(_01742_),
    .B(_01744_),
    .C(_01871_),
    .Y(_01873_));
 sky130_fd_sc_hd__and3_1 _20699_ (.A(_01859_),
    .B(_01872_),
    .C(_01873_),
    .X(_01874_));
 sky130_fd_sc_hd__inv_2 _20700_ (.A(_01874_),
    .Y(_01875_));
 sky130_fd_sc_hd__a21oi_1 _20701_ (.A1(_01872_),
    .A2(_01873_),
    .B1(_01859_),
    .Y(_01876_));
 sky130_fd_sc_hd__a211o_1 _20702_ (.A1(_01706_),
    .A2(_01708_),
    .B1(_01874_),
    .C1(_01876_),
    .X(_01877_));
 sky130_fd_sc_hd__inv_2 _20703_ (.A(_01877_),
    .Y(_01878_));
 sky130_fd_sc_hd__o211ai_1 _20704_ (.A1(_01874_),
    .A2(_01876_),
    .B1(_01706_),
    .C1(_01708_),
    .Y(_01879_));
 sky130_fd_sc_hd__nand2_1 _20705_ (.A(_01877_),
    .B(_01879_),
    .Y(_01880_));
 sky130_fd_sc_hd__a21oi_1 _20706_ (.A1(_01746_),
    .A2(_01748_),
    .B1(_01880_),
    .Y(_01881_));
 sky130_fd_sc_hd__and3_1 _20707_ (.A(_01746_),
    .B(_01748_),
    .C(_01880_),
    .X(_01882_));
 sky130_fd_sc_hd__or3_1 _20708_ (.A(_01842_),
    .B(_01881_),
    .C(_01882_),
    .X(_01883_));
 sky130_fd_sc_hd__o21ai_1 _20709_ (.A1(_01881_),
    .A2(_01882_),
    .B1(_01842_),
    .Y(_01884_));
 sky130_fd_sc_hd__and2_1 _20710_ (.A(_01883_),
    .B(_01884_),
    .X(_01885_));
 sky130_fd_sc_hd__o21ai_4 _20711_ (.A1(_01715_),
    .A2(_01754_),
    .B1(_01885_),
    .Y(_01886_));
 sky130_fd_sc_hd__or3_2 _20712_ (.A(_01715_),
    .B(_01754_),
    .C(_01885_),
    .X(_01887_));
 sky130_fd_sc_hd__a22o_1 _20713_ (.A1(net628),
    .A2(net72),
    .B1(net69),
    .B2(net250),
    .X(_01888_));
 sky130_fd_sc_hd__and4_1 _20714_ (.A(net628),
    .B(net250),
    .C(net72),
    .D(net69),
    .X(_01889_));
 sky130_fd_sc_hd__inv_2 _20715_ (.A(_01889_),
    .Y(_01890_));
 sky130_fd_sc_hd__a22oi_1 _20716_ (.A1(net255),
    .A2(net66),
    .B1(_01888_),
    .B2(_01890_),
    .Y(_01891_));
 sky130_fd_sc_hd__and4_1 _20717_ (.A(net255),
    .B(net66),
    .C(_01888_),
    .D(_01890_),
    .X(_01892_));
 sky130_fd_sc_hd__or2_2 _20718_ (.A(_01891_),
    .B(_01892_),
    .X(_01893_));
 sky130_fd_sc_hd__nor2_2 _20719_ (.A(_01759_),
    .B(_01762_),
    .Y(_01894_));
 sky130_fd_sc_hd__xnor2_2 _20720_ (.A(_01893_),
    .B(_01894_),
    .Y(_01895_));
 sky130_fd_sc_hd__and4b_2 _20721_ (.A_N(net265),
    .B(net63),
    .C(net62),
    .D(net261),
    .X(_01896_));
 sky130_fd_sc_hd__o2bb2a_1 _20722_ (.A1_N(net261),
    .A2_N(net63),
    .B1(net56),
    .B2(net265),
    .X(_01897_));
 sky130_fd_sc_hd__nor2_1 _20723_ (.A(_01896_),
    .B(_01897_),
    .Y(_01898_));
 sky130_fd_sc_hd__xnor2_2 _20724_ (.A(_01895_),
    .B(_01898_),
    .Y(_01899_));
 sky130_fd_sc_hd__o32ai_4 _20725_ (.A1(_01765_),
    .A2(_01766_),
    .A3(_01768_),
    .B1(_01764_),
    .B2(_01763_),
    .Y(_01900_));
 sky130_fd_sc_hd__xnor2_1 _20726_ (.A(_01899_),
    .B(_01900_),
    .Y(_01901_));
 sky130_fd_sc_hd__nor2_1 _20727_ (.A(_01767_),
    .B(_01901_),
    .Y(_01902_));
 sky130_fd_sc_hd__xnor2_1 _20728_ (.A(_01767_),
    .B(_01901_),
    .Y(_01903_));
 sky130_fd_sc_hd__or2_1 _20729_ (.A(_01782_),
    .B(_01784_),
    .X(_01904_));
 sky130_fd_sc_hd__nand2_1 _20730_ (.A(_01718_),
    .B(_01720_),
    .Y(_01905_));
 sky130_fd_sc_hd__a22o_1 _20731_ (.A1(net237),
    .A2(net83),
    .B1(net79),
    .B2(net241),
    .X(_01906_));
 sky130_fd_sc_hd__inv_2 _20732_ (.A(_01906_),
    .Y(_01907_));
 sky130_fd_sc_hd__and4_1 _20733_ (.A(net241),
    .B(net237),
    .C(net84),
    .D(net79),
    .X(_01908_));
 sky130_fd_sc_hd__o2bb2a_1 _20734_ (.A1_N(net246),
    .A2_N(net76),
    .B1(_01907_),
    .B2(_01908_),
    .X(_01909_));
 sky130_fd_sc_hd__and4b_1 _20735_ (.A_N(_01908_),
    .B(net76),
    .C(net246),
    .D(_01906_),
    .X(_01910_));
 sky130_fd_sc_hd__or2_1 _20736_ (.A(_01909_),
    .B(_01910_),
    .X(_01911_));
 sky130_fd_sc_hd__nand2b_1 _20737_ (.A_N(_01911_),
    .B(_01905_),
    .Y(_01912_));
 sky130_fd_sc_hd__xnor2_1 _20738_ (.A(_01905_),
    .B(_01911_),
    .Y(_01913_));
 sky130_fd_sc_hd__nand2_1 _20739_ (.A(_01904_),
    .B(_01913_),
    .Y(_01914_));
 sky130_fd_sc_hd__xnor2_1 _20740_ (.A(_01904_),
    .B(_01913_),
    .Y(_01915_));
 sky130_fd_sc_hd__a21oi_2 _20741_ (.A1(_01729_),
    .A2(_01731_),
    .B1(_01915_),
    .Y(_01916_));
 sky130_fd_sc_hd__and3_1 _20742_ (.A(_01729_),
    .B(_01731_),
    .C(_01915_),
    .X(_01917_));
 sky130_fd_sc_hd__a211oi_2 _20743_ (.A1(_01786_),
    .A2(_01788_),
    .B1(_01916_),
    .C1(_01917_),
    .Y(_01918_));
 sky130_fd_sc_hd__o211a_1 _20744_ (.A1(_01916_),
    .A2(_01917_),
    .B1(_01786_),
    .C1(_01788_),
    .X(_01919_));
 sky130_fd_sc_hd__a211oi_1 _20745_ (.A1(_01791_),
    .A2(_01793_),
    .B1(_01918_),
    .C1(_01919_),
    .Y(_01920_));
 sky130_fd_sc_hd__o211a_1 _20746_ (.A1(_01918_),
    .A2(_01919_),
    .B1(_01791_),
    .C1(_01793_),
    .X(_01921_));
 sky130_fd_sc_hd__or3_1 _20747_ (.A(_01903_),
    .B(_01920_),
    .C(_01921_),
    .X(_01922_));
 sky130_fd_sc_hd__o21ai_1 _20748_ (.A1(_01920_),
    .A2(_01921_),
    .B1(_01903_),
    .Y(_01923_));
 sky130_fd_sc_hd__o211a_2 _20749_ (.A1(_01750_),
    .A2(_01752_),
    .B1(_01922_),
    .C1(_01923_),
    .X(_01924_));
 sky130_fd_sc_hd__inv_2 _20750_ (.A(_01924_),
    .Y(_01925_));
 sky130_fd_sc_hd__a211o_1 _20751_ (.A1(_01922_),
    .A2(_01923_),
    .B1(_01750_),
    .C1(_01752_),
    .X(_01926_));
 sky130_fd_sc_hd__o211a_2 _20752_ (.A1(_01795_),
    .A2(_01797_),
    .B1(_01925_),
    .C1(_01926_),
    .X(_01927_));
 sky130_fd_sc_hd__inv_2 _20753_ (.A(_01927_),
    .Y(_01928_));
 sky130_fd_sc_hd__a211o_1 _20754_ (.A1(_01925_),
    .A2(_01926_),
    .B1(_01795_),
    .C1(_01797_),
    .X(_01929_));
 sky130_fd_sc_hd__nand4_4 _20755_ (.A(_01886_),
    .B(_01887_),
    .C(_01928_),
    .D(_01929_),
    .Y(_01930_));
 sky130_fd_sc_hd__a22o_1 _20756_ (.A1(_01886_),
    .A2(_01887_),
    .B1(_01928_),
    .B2(_01929_),
    .X(_01931_));
 sky130_fd_sc_hd__o211a_2 _20757_ (.A1(_01756_),
    .A2(_01803_),
    .B1(_01930_),
    .C1(_01931_),
    .X(_01932_));
 sky130_fd_sc_hd__a211oi_2 _20758_ (.A1(_01930_),
    .A2(_01931_),
    .B1(_01756_),
    .C1(_01803_),
    .Y(_01933_));
 sky130_fd_sc_hd__a211oi_4 _20759_ (.A1(_01799_),
    .A2(_01801_),
    .B1(_01932_),
    .C1(_01933_),
    .Y(_01934_));
 sky130_fd_sc_hd__o211a_1 _20760_ (.A1(_01932_),
    .A2(_01933_),
    .B1(_01799_),
    .C1(_01801_),
    .X(_01935_));
 sky130_fd_sc_hd__a211oi_2 _20761_ (.A1(_01806_),
    .A2(_01808_),
    .B1(_01934_),
    .C1(_01935_),
    .Y(_01936_));
 sky130_fd_sc_hd__o211a_1 _20762_ (.A1(_01934_),
    .A2(_01935_),
    .B1(_01806_),
    .C1(_01808_),
    .X(_01937_));
 sky130_fd_sc_hd__a211oi_2 _20763_ (.A1(_01772_),
    .A2(_01775_),
    .B1(_01936_),
    .C1(_01937_),
    .Y(_01938_));
 sky130_fd_sc_hd__o211a_1 _20764_ (.A1(_01936_),
    .A2(_01937_),
    .B1(_01772_),
    .C1(_01775_),
    .X(_01939_));
 sky130_fd_sc_hd__o211a_1 _20765_ (.A1(_01938_),
    .A2(_01939_),
    .B1(_01810_),
    .C1(_01812_),
    .X(_01940_));
 sky130_fd_sc_hd__a211o_1 _20766_ (.A1(_01810_),
    .A2(_01812_),
    .B1(_01938_),
    .C1(_01939_),
    .X(_01941_));
 sky130_fd_sc_hd__and2b_1 _20767_ (.A_N(_01940_),
    .B(_01941_),
    .X(_01942_));
 sky130_fd_sc_hd__a21oi_1 _20768_ (.A1(_01817_),
    .A2(_01820_),
    .B1(_01816_),
    .Y(_01943_));
 sky130_fd_sc_hd__xnor2_2 _20769_ (.A(_01942_),
    .B(_01943_),
    .Y(_01944_));
 sky130_fd_sc_hd__and3_1 _20770_ (.A(net770),
    .B(_03049_),
    .C(net43),
    .X(_01945_));
 sky130_fd_sc_hd__a221o_1 _20771_ (.A1(_03052_),
    .A2(_07365_),
    .B1(_01944_),
    .B2(net10),
    .C1(_01945_),
    .X(_01946_));
 sky130_fd_sc_hd__mux2_1 _20772_ (.A0(net872),
    .A1(_01946_),
    .S(net2),
    .X(_00325_));
 sky130_fd_sc_hd__o21ai_1 _20773_ (.A1(_01831_),
    .A2(_01832_),
    .B1(_01825_),
    .Y(_01947_));
 sky130_fd_sc_hd__and3_1 _20774_ (.A(net137),
    .B(net132),
    .C(net194),
    .X(_01948_));
 sky130_fd_sc_hd__o21ai_1 _20775_ (.A1(net137),
    .A2(net132),
    .B1(net194),
    .Y(_01949_));
 sky130_fd_sc_hd__nor2_2 _20776_ (.A(_01948_),
    .B(_01949_),
    .Y(_01950_));
 sky130_fd_sc_hd__nand2_1 _20777_ (.A(net128),
    .B(net196),
    .Y(_01951_));
 sky130_fd_sc_hd__xor2_1 _20778_ (.A(_01950_),
    .B(_01951_),
    .X(_01952_));
 sky130_fd_sc_hd__nor2_1 _20779_ (.A(_01832_),
    .B(_01952_),
    .Y(_01953_));
 sky130_fd_sc_hd__and2_1 _20780_ (.A(_01832_),
    .B(_01952_),
    .X(_01954_));
 sky130_fd_sc_hd__nor2_1 _20781_ (.A(_01953_),
    .B(_01954_),
    .Y(_01955_));
 sky130_fd_sc_hd__nand2_1 _20782_ (.A(_01563_),
    .B(_01955_),
    .Y(_01956_));
 sky130_fd_sc_hd__or2_1 _20783_ (.A(_01563_),
    .B(_01955_),
    .X(_01957_));
 sky130_fd_sc_hd__and2_1 _20784_ (.A(_01956_),
    .B(_01957_),
    .X(_01958_));
 sky130_fd_sc_hd__nand2_1 _20785_ (.A(_01947_),
    .B(_01958_),
    .Y(_01959_));
 sky130_fd_sc_hd__xnor2_1 _20786_ (.A(_01947_),
    .B(_01958_),
    .Y(_01960_));
 sky130_fd_sc_hd__xnor2_1 _20787_ (.A(_01559_),
    .B(_01960_),
    .Y(_01961_));
 sky130_fd_sc_hd__nor3_1 _20788_ (.A(_01557_),
    .B(_01838_),
    .C(_01961_),
    .Y(_01962_));
 sky130_fd_sc_hd__o21a_1 _20789_ (.A1(_01557_),
    .A2(_01838_),
    .B1(_01961_),
    .X(_01963_));
 sky130_fd_sc_hd__or2_1 _20790_ (.A(_01962_),
    .B(_01963_),
    .X(_01964_));
 sky130_fd_sc_hd__a22o_1 _20791_ (.A1(net222),
    .A2(net91),
    .B1(net217),
    .B2(net97),
    .X(_01965_));
 sky130_fd_sc_hd__nand4_2 _20792_ (.A(net97),
    .B(net222),
    .C(net91),
    .D(net217),
    .Y(_01966_));
 sky130_fd_sc_hd__a22o_1 _20793_ (.A1(net226),
    .A2(net86),
    .B1(_01965_),
    .B2(_01966_),
    .X(_01967_));
 sky130_fd_sc_hd__nand4_1 _20794_ (.A(net226),
    .B(net86),
    .C(_01965_),
    .D(_01966_),
    .Y(_01968_));
 sky130_fd_sc_hd__nand2_1 _20795_ (.A(_01967_),
    .B(_01968_),
    .Y(_01969_));
 sky130_fd_sc_hd__a22o_1 _20796_ (.A1(net102),
    .A2(net210),
    .B1(net207),
    .B2(net107),
    .X(_01970_));
 sky130_fd_sc_hd__and4_1 _20797_ (.A(net107),
    .B(net102),
    .C(\mul1.a[25] ),
    .D(net207),
    .X(_01971_));
 sky130_fd_sc_hd__inv_2 _20798_ (.A(_01971_),
    .Y(_01972_));
 sky130_fd_sc_hd__a22oi_1 _20799_ (.A1(net98),
    .A2(net213),
    .B1(_01970_),
    .B2(_01972_),
    .Y(_01973_));
 sky130_fd_sc_hd__and4_1 _20800_ (.A(net98),
    .B(net213),
    .C(_01970_),
    .D(_01972_),
    .X(_01974_));
 sky130_fd_sc_hd__or2_1 _20801_ (.A(_01849_),
    .B(_01852_),
    .X(_01975_));
 sky130_fd_sc_hd__or3b_2 _20802_ (.A(_01973_),
    .B(_01974_),
    .C_N(_01975_),
    .X(_01976_));
 sky130_fd_sc_hd__o21bai_1 _20803_ (.A1(_01973_),
    .A2(_01974_),
    .B1_N(_01975_),
    .Y(_01977_));
 sky130_fd_sc_hd__nand2_1 _20804_ (.A(_01976_),
    .B(_01977_),
    .Y(_01978_));
 sky130_fd_sc_hd__or2_1 _20805_ (.A(_01969_),
    .B(_01978_),
    .X(_01979_));
 sky130_fd_sc_hd__nand2_1 _20806_ (.A(_01969_),
    .B(_01978_),
    .Y(_01980_));
 sky130_fd_sc_hd__and2_1 _20807_ (.A(_01979_),
    .B(_01980_),
    .X(_01981_));
 sky130_fd_sc_hd__or2_1 _20808_ (.A(_01864_),
    .B(_01866_),
    .X(_01982_));
 sky130_fd_sc_hd__a31o_1 _20809_ (.A1(net128),
    .A2(\mul1.a[29] ),
    .A3(_01829_),
    .B1(_01828_),
    .X(_01983_));
 sky130_fd_sc_hd__a22o_1 _20810_ (.A1(net121),
    .A2(net201),
    .B1(\mul1.a[29] ),
    .B2(net123),
    .X(_01984_));
 sky130_fd_sc_hd__inv_2 _20811_ (.A(_01984_),
    .Y(_01985_));
 sky130_fd_sc_hd__and4_1 _20812_ (.A(net123),
    .B(net118),
    .C(net201),
    .D(\mul1.a[29] ),
    .X(_01986_));
 sky130_fd_sc_hd__o2bb2a_1 _20813_ (.A1_N(net113),
    .A2_N(net204),
    .B1(_01985_),
    .B2(_01986_),
    .X(_01987_));
 sky130_fd_sc_hd__and4b_1 _20814_ (.A_N(_01986_),
    .B(net204),
    .C(net113),
    .D(_01984_),
    .X(_01988_));
 sky130_fd_sc_hd__or2_1 _20815_ (.A(_01987_),
    .B(_01988_),
    .X(_01989_));
 sky130_fd_sc_hd__nand2b_1 _20816_ (.A_N(_01989_),
    .B(_01983_),
    .Y(_01990_));
 sky130_fd_sc_hd__xnor2_1 _20817_ (.A(_01983_),
    .B(_01989_),
    .Y(_01991_));
 sky130_fd_sc_hd__nand2_1 _20818_ (.A(_01982_),
    .B(_01991_),
    .Y(_01992_));
 sky130_fd_sc_hd__or2_1 _20819_ (.A(_01982_),
    .B(_01991_),
    .X(_01993_));
 sky130_fd_sc_hd__nand2_1 _20820_ (.A(_01992_),
    .B(_01993_),
    .Y(_01994_));
 sky130_fd_sc_hd__a21o_1 _20821_ (.A1(_01868_),
    .A2(_01870_),
    .B1(_01994_),
    .X(_01995_));
 sky130_fd_sc_hd__inv_2 _20822_ (.A(_01995_),
    .Y(_01996_));
 sky130_fd_sc_hd__nand3_1 _20823_ (.A(_01868_),
    .B(_01870_),
    .C(_01994_),
    .Y(_01997_));
 sky130_fd_sc_hd__and3_2 _20824_ (.A(_01981_),
    .B(_01995_),
    .C(_01997_),
    .X(_01998_));
 sky130_fd_sc_hd__a21oi_2 _20825_ (.A1(_01995_),
    .A2(_01997_),
    .B1(_01981_),
    .Y(_01999_));
 sky130_fd_sc_hd__a211oi_4 _20826_ (.A1(_01834_),
    .A2(_01836_),
    .B1(_01998_),
    .C1(_01999_),
    .Y(_02000_));
 sky130_fd_sc_hd__o211a_1 _20827_ (.A1(_01998_),
    .A2(_01999_),
    .B1(_01834_),
    .C1(_01836_),
    .X(_02001_));
 sky130_fd_sc_hd__a211oi_4 _20828_ (.A1(_01872_),
    .A2(_01875_),
    .B1(_02000_),
    .C1(_02001_),
    .Y(_02002_));
 sky130_fd_sc_hd__o211a_1 _20829_ (.A1(_02000_),
    .A2(_02001_),
    .B1(_01872_),
    .C1(_01875_),
    .X(_02003_));
 sky130_fd_sc_hd__nor3_2 _20830_ (.A(_01964_),
    .B(_02002_),
    .C(_02003_),
    .Y(_02004_));
 sky130_fd_sc_hd__o21a_1 _20831_ (.A1(_02002_),
    .A2(_02003_),
    .B1(_01964_),
    .X(_02005_));
 sky130_fd_sc_hd__a211oi_2 _20832_ (.A1(_01841_),
    .A2(_01883_),
    .B1(_02004_),
    .C1(_02005_),
    .Y(_02006_));
 sky130_fd_sc_hd__o211a_1 _20833_ (.A1(_02004_),
    .A2(_02005_),
    .B1(_01841_),
    .C1(_01883_),
    .X(_02007_));
 sky130_fd_sc_hd__nor2_1 _20834_ (.A(_02006_),
    .B(_02007_),
    .Y(_02008_));
 sky130_fd_sc_hd__nand2b_1 _20835_ (.A_N(_01920_),
    .B(_01922_),
    .Y(_02009_));
 sky130_fd_sc_hd__nor2_1 _20836_ (.A(_01878_),
    .B(_01881_),
    .Y(_02010_));
 sky130_fd_sc_hd__a22o_1 _20837_ (.A1(net245),
    .A2(net72),
    .B1(net69),
    .B2(net628),
    .X(_02011_));
 sky130_fd_sc_hd__and4_1 _20838_ (.A(net245),
    .B(net628),
    .C(net73),
    .D(net70),
    .X(_02012_));
 sky130_fd_sc_hd__inv_2 _20839_ (.A(_02012_),
    .Y(_02013_));
 sky130_fd_sc_hd__a22oi_1 _20840_ (.A1(net250),
    .A2(net66),
    .B1(_02011_),
    .B2(_02013_),
    .Y(_02014_));
 sky130_fd_sc_hd__and4_1 _20841_ (.A(net250),
    .B(net67),
    .C(_02011_),
    .D(_02013_),
    .X(_02015_));
 sky130_fd_sc_hd__or2_2 _20842_ (.A(_02014_),
    .B(_02015_),
    .X(_02016_));
 sky130_fd_sc_hd__nor2_2 _20843_ (.A(_01889_),
    .B(_01892_),
    .Y(_02017_));
 sky130_fd_sc_hd__xnor2_2 _20844_ (.A(_02016_),
    .B(_02017_),
    .Y(_02018_));
 sky130_fd_sc_hd__and4b_2 _20845_ (.A_N(net261),
    .B(net63),
    .C(\mul1.b[31] ),
    .D(net255),
    .X(_02019_));
 sky130_fd_sc_hd__inv_2 _20846_ (.A(_02019_),
    .Y(_02020_));
 sky130_fd_sc_hd__o2bb2a_1 _20847_ (.A1_N(net255),
    .A2_N(net63),
    .B1(_02568_),
    .B2(net261),
    .X(_02021_));
 sky130_fd_sc_hd__nor2_1 _20848_ (.A(_02019_),
    .B(_02021_),
    .Y(_02022_));
 sky130_fd_sc_hd__xnor2_1 _20849_ (.A(_02018_),
    .B(_02022_),
    .Y(_02023_));
 sky130_fd_sc_hd__o32ai_4 _20850_ (.A1(_01895_),
    .A2(_01896_),
    .A3(_01897_),
    .B1(_01894_),
    .B2(_01893_),
    .Y(_02024_));
 sky130_fd_sc_hd__nand2_1 _20851_ (.A(_02023_),
    .B(_02024_),
    .Y(_02025_));
 sky130_fd_sc_hd__xnor2_1 _20852_ (.A(_02023_),
    .B(_02024_),
    .Y(_02026_));
 sky130_fd_sc_hd__inv_2 _20853_ (.A(_02026_),
    .Y(_02027_));
 sky130_fd_sc_hd__nand2_1 _20854_ (.A(_01896_),
    .B(_02027_),
    .Y(_02028_));
 sky130_fd_sc_hd__or2_1 _20855_ (.A(_01896_),
    .B(_02027_),
    .X(_02029_));
 sky130_fd_sc_hd__nand2_1 _20856_ (.A(_02028_),
    .B(_02029_),
    .Y(_02030_));
 sky130_fd_sc_hd__or2_1 _20857_ (.A(_01908_),
    .B(_01910_),
    .X(_02031_));
 sky130_fd_sc_hd__nand2_1 _20858_ (.A(_01844_),
    .B(_01846_),
    .Y(_02032_));
 sky130_fd_sc_hd__a22o_1 _20859_ (.A1(net230),
    .A2(net83),
    .B1(net79),
    .B2(net237),
    .X(_02033_));
 sky130_fd_sc_hd__inv_2 _20860_ (.A(_02033_),
    .Y(_02034_));
 sky130_fd_sc_hd__and4_1 _20861_ (.A(net237),
    .B(net230),
    .C(net83),
    .D(net79),
    .X(_02035_));
 sky130_fd_sc_hd__o2bb2a_1 _20862_ (.A1_N(net241),
    .A2_N(net76),
    .B1(_02034_),
    .B2(_02035_),
    .X(_02036_));
 sky130_fd_sc_hd__and4b_1 _20863_ (.A_N(_02035_),
    .B(net76),
    .C(net241),
    .D(_02033_),
    .X(_02037_));
 sky130_fd_sc_hd__or2_1 _20864_ (.A(_02036_),
    .B(_02037_),
    .X(_02038_));
 sky130_fd_sc_hd__nand2b_1 _20865_ (.A_N(_02038_),
    .B(_02032_),
    .Y(_02039_));
 sky130_fd_sc_hd__xnor2_1 _20866_ (.A(_02032_),
    .B(_02038_),
    .Y(_02040_));
 sky130_fd_sc_hd__nand2_1 _20867_ (.A(_02031_),
    .B(_02040_),
    .Y(_02041_));
 sky130_fd_sc_hd__or2_1 _20868_ (.A(_02031_),
    .B(_02040_),
    .X(_02042_));
 sky130_fd_sc_hd__nand2_1 _20869_ (.A(_02041_),
    .B(_02042_),
    .Y(_02043_));
 sky130_fd_sc_hd__a21oi_1 _20870_ (.A1(_01855_),
    .A2(_01857_),
    .B1(_02043_),
    .Y(_02044_));
 sky130_fd_sc_hd__a21o_1 _20871_ (.A1(_01855_),
    .A2(_01857_),
    .B1(_02043_),
    .X(_02045_));
 sky130_fd_sc_hd__and3_1 _20872_ (.A(_01855_),
    .B(_01857_),
    .C(_02043_),
    .X(_02046_));
 sky130_fd_sc_hd__a211o_1 _20873_ (.A1(_01912_),
    .A2(_01914_),
    .B1(_02044_),
    .C1(_02046_),
    .X(_02047_));
 sky130_fd_sc_hd__o211ai_1 _20874_ (.A1(_02044_),
    .A2(_02046_),
    .B1(_01912_),
    .C1(_01914_),
    .Y(_02048_));
 sky130_fd_sc_hd__o211a_1 _20875_ (.A1(_01916_),
    .A2(_01918_),
    .B1(_02047_),
    .C1(_02048_),
    .X(_02049_));
 sky130_fd_sc_hd__a211oi_1 _20876_ (.A1(_02047_),
    .A2(_02048_),
    .B1(_01916_),
    .C1(_01918_),
    .Y(_02050_));
 sky130_fd_sc_hd__nor3_1 _20877_ (.A(_02030_),
    .B(_02049_),
    .C(_02050_),
    .Y(_02051_));
 sky130_fd_sc_hd__o21a_1 _20878_ (.A1(_02049_),
    .A2(_02050_),
    .B1(_02030_),
    .X(_02052_));
 sky130_fd_sc_hd__nor2_1 _20879_ (.A(_02051_),
    .B(_02052_),
    .Y(_02053_));
 sky130_fd_sc_hd__or3_1 _20880_ (.A(_02010_),
    .B(_02051_),
    .C(_02052_),
    .X(_02054_));
 sky130_fd_sc_hd__xnor2_1 _20881_ (.A(_02010_),
    .B(_02053_),
    .Y(_02055_));
 sky130_fd_sc_hd__nand2_1 _20882_ (.A(_02009_),
    .B(_02055_),
    .Y(_02056_));
 sky130_fd_sc_hd__xor2_1 _20883_ (.A(_02009_),
    .B(_02055_),
    .X(_02057_));
 sky130_fd_sc_hd__and2_2 _20884_ (.A(_02008_),
    .B(_02057_),
    .X(_02058_));
 sky130_fd_sc_hd__nor2_1 _20885_ (.A(_02008_),
    .B(_02057_),
    .Y(_02059_));
 sky130_fd_sc_hd__a211o_2 _20886_ (.A1(_01886_),
    .A2(_01930_),
    .B1(_02058_),
    .C1(_02059_),
    .X(_02060_));
 sky130_fd_sc_hd__o211ai_4 _20887_ (.A1(_02058_),
    .A2(_02059_),
    .B1(_01886_),
    .C1(_01930_),
    .Y(_02061_));
 sky130_fd_sc_hd__o211ai_4 _20888_ (.A1(_01924_),
    .A2(_01927_),
    .B1(_02060_),
    .C1(_02061_),
    .Y(_02062_));
 sky130_fd_sc_hd__a211o_1 _20889_ (.A1(_02060_),
    .A2(_02061_),
    .B1(_01924_),
    .C1(_01927_),
    .X(_02063_));
 sky130_fd_sc_hd__o211ai_4 _20890_ (.A1(_01932_),
    .A2(_01934_),
    .B1(_02062_),
    .C1(_02063_),
    .Y(_02064_));
 sky130_fd_sc_hd__a211o_1 _20891_ (.A1(_02062_),
    .A2(_02063_),
    .B1(_01932_),
    .C1(_01934_),
    .X(_02065_));
 sky130_fd_sc_hd__nand2_1 _20892_ (.A(_02064_),
    .B(_02065_),
    .Y(_02066_));
 sky130_fd_sc_hd__a21oi_2 _20893_ (.A1(_01899_),
    .A2(_01900_),
    .B1(_01902_),
    .Y(_02067_));
 sky130_fd_sc_hd__or2_1 _20894_ (.A(_02066_),
    .B(_02067_),
    .X(_02068_));
 sky130_fd_sc_hd__xnor2_2 _20895_ (.A(_02066_),
    .B(_02067_),
    .Y(_02069_));
 sky130_fd_sc_hd__or2_1 _20896_ (.A(_01936_),
    .B(_01938_),
    .X(_02070_));
 sky130_fd_sc_hd__and2b_1 _20897_ (.A_N(_02069_),
    .B(_02070_),
    .X(_02071_));
 sky130_fd_sc_hd__xnor2_2 _20898_ (.A(_02069_),
    .B(_02070_),
    .Y(_02072_));
 sky130_fd_sc_hd__inv_2 _20899_ (.A(_02072_),
    .Y(_02073_));
 sky130_fd_sc_hd__nand2_1 _20900_ (.A(_01817_),
    .B(_01942_),
    .Y(_02074_));
 sky130_fd_sc_hd__or4b_2 _20901_ (.A(_01552_),
    .B(_01689_),
    .C(_02074_),
    .D_N(_01549_),
    .X(_02075_));
 sky130_fd_sc_hd__or2_1 _20902_ (.A(_01818_),
    .B(_02074_),
    .X(_02076_));
 sky130_fd_sc_hd__or3b_2 _20903_ (.A(_01940_),
    .B(_01814_),
    .C_N(_01815_),
    .X(_02077_));
 sky130_fd_sc_hd__and4_1 _20904_ (.A(_01941_),
    .B(_02075_),
    .C(_02076_),
    .D(_02077_),
    .X(_02078_));
 sky130_fd_sc_hd__a41oi_4 _20905_ (.A1(_01941_),
    .A2(_02075_),
    .A3(_02076_),
    .A4(_02077_),
    .B1(_02073_),
    .Y(_02079_));
 sky130_fd_sc_hd__xnor2_1 _20906_ (.A(_02072_),
    .B(_02078_),
    .Y(_02080_));
 sky130_fd_sc_hd__nor2_1 _20907_ (.A(net43),
    .B(_07499_),
    .Y(_02081_));
 sky130_fd_sc_hd__a221o_1 _20908_ (.A1(net763),
    .A2(net8),
    .B1(_02080_),
    .B2(net10),
    .C1(_02081_),
    .X(_02082_));
 sky130_fd_sc_hd__mux2_1 _20909_ (.A0(net791),
    .A1(_02082_),
    .S(net2),
    .X(_00326_));
 sky130_fd_sc_hd__nand2_2 _20910_ (.A(net128),
    .B(net194),
    .Y(_02083_));
 sky130_fd_sc_hd__xor2_4 _20911_ (.A(_01950_),
    .B(_02083_),
    .X(_02084_));
 sky130_fd_sc_hd__xor2_4 _20912_ (.A(_01832_),
    .B(_02084_),
    .X(_02085_));
 sky130_fd_sc_hd__nand2_1 _20913_ (.A(_01563_),
    .B(_02085_),
    .Y(_02086_));
 sky130_fd_sc_hd__xnor2_4 _20914_ (.A(_01562_),
    .B(_02085_),
    .Y(_02087_));
 sky130_fd_sc_hd__o21ai_2 _20915_ (.A1(_01824_),
    .A2(_01953_),
    .B1(_02087_),
    .Y(_02088_));
 sky130_fd_sc_hd__or3_1 _20916_ (.A(_01824_),
    .B(_01953_),
    .C(_02087_),
    .X(_02089_));
 sky130_fd_sc_hd__nand2_1 _20917_ (.A(_02088_),
    .B(_02089_),
    .Y(_02090_));
 sky130_fd_sc_hd__xnor2_1 _20918_ (.A(_01560_),
    .B(_02090_),
    .Y(_02091_));
 sky130_fd_sc_hd__o21ba_1 _20919_ (.A1(_01560_),
    .A2(_01960_),
    .B1_N(_01557_),
    .X(_02092_));
 sky130_fd_sc_hd__xnor2_1 _20920_ (.A(_02091_),
    .B(_02092_),
    .Y(_02093_));
 sky130_fd_sc_hd__a22o_1 _20921_ (.A1(net91),
    .A2(net217),
    .B1(net213),
    .B2(net97),
    .X(_02094_));
 sky130_fd_sc_hd__nand4_1 _20922_ (.A(net97),
    .B(net91),
    .C(net217),
    .D(net213),
    .Y(_02095_));
 sky130_fd_sc_hd__a22o_1 _20923_ (.A1(net222),
    .A2(net86),
    .B1(_02094_),
    .B2(_02095_),
    .X(_02096_));
 sky130_fd_sc_hd__nand4_1 _20924_ (.A(net222),
    .B(net86),
    .C(_02094_),
    .D(_02095_),
    .Y(_02097_));
 sky130_fd_sc_hd__nand2_1 _20925_ (.A(_02096_),
    .B(_02097_),
    .Y(_02098_));
 sky130_fd_sc_hd__a22o_1 _20926_ (.A1(net102),
    .A2(net207),
    .B1(net204),
    .B2(net112),
    .X(_02099_));
 sky130_fd_sc_hd__and4_1 _20927_ (.A(net112),
    .B(\mul1.b[19] ),
    .C(\mul1.a[26] ),
    .D(net204),
    .X(_02100_));
 sky130_fd_sc_hd__inv_2 _20928_ (.A(_02100_),
    .Y(_02101_));
 sky130_fd_sc_hd__a22oi_1 _20929_ (.A1(\mul1.b[20] ),
    .A2(net210),
    .B1(_02099_),
    .B2(_02101_),
    .Y(_02102_));
 sky130_fd_sc_hd__and4_1 _20930_ (.A(\mul1.b[20] ),
    .B(\mul1.a[25] ),
    .C(_02099_),
    .D(_02101_),
    .X(_02103_));
 sky130_fd_sc_hd__or2_1 _20931_ (.A(_01971_),
    .B(_01974_),
    .X(_02104_));
 sky130_fd_sc_hd__or3b_2 _20932_ (.A(_02102_),
    .B(_02103_),
    .C_N(_02104_),
    .X(_02105_));
 sky130_fd_sc_hd__o21bai_1 _20933_ (.A1(_02102_),
    .A2(_02103_),
    .B1_N(_02104_),
    .Y(_02106_));
 sky130_fd_sc_hd__nand2_1 _20934_ (.A(_02105_),
    .B(_02106_),
    .Y(_02107_));
 sky130_fd_sc_hd__or2_1 _20935_ (.A(_02098_),
    .B(_02107_),
    .X(_02108_));
 sky130_fd_sc_hd__nand2_1 _20936_ (.A(_02098_),
    .B(_02107_),
    .Y(_02109_));
 sky130_fd_sc_hd__and2_1 _20937_ (.A(_02108_),
    .B(_02109_),
    .X(_02110_));
 sky130_fd_sc_hd__or2_1 _20938_ (.A(_01986_),
    .B(_01988_),
    .X(_02111_));
 sky130_fd_sc_hd__a31o_1 _20939_ (.A1(net128),
    .A2(net196),
    .A3(_01950_),
    .B1(_01948_),
    .X(_02112_));
 sky130_fd_sc_hd__a22o_1 _20940_ (.A1(net118),
    .A2(\mul1.a[29] ),
    .B1(\mul1.a[30] ),
    .B2(net123),
    .X(_02113_));
 sky130_fd_sc_hd__and4_1 _20941_ (.A(net123),
    .B(net118),
    .C(\mul1.a[29] ),
    .D(\mul1.a[30] ),
    .X(_02114_));
 sky130_fd_sc_hd__inv_2 _20942_ (.A(_02114_),
    .Y(_02115_));
 sky130_fd_sc_hd__a22o_1 _20943_ (.A1(net113),
    .A2(net201),
    .B1(_02113_),
    .B2(_02115_),
    .X(_02116_));
 sky130_fd_sc_hd__and4_1 _20944_ (.A(net113),
    .B(net201),
    .C(_02113_),
    .D(_02115_),
    .X(_02117_));
 sky130_fd_sc_hd__inv_2 _20945_ (.A(_02117_),
    .Y(_02118_));
 sky130_fd_sc_hd__and3_1 _20946_ (.A(_02112_),
    .B(_02116_),
    .C(_02118_),
    .X(_02119_));
 sky130_fd_sc_hd__a21o_1 _20947_ (.A1(_02116_),
    .A2(_02118_),
    .B1(_02112_),
    .X(_02120_));
 sky130_fd_sc_hd__and2b_1 _20948_ (.A_N(_02119_),
    .B(_02120_),
    .X(_02121_));
 sky130_fd_sc_hd__xnor2_1 _20949_ (.A(_02111_),
    .B(_02121_),
    .Y(_02122_));
 sky130_fd_sc_hd__a21o_1 _20950_ (.A1(_01990_),
    .A2(_01992_),
    .B1(_02122_),
    .X(_02123_));
 sky130_fd_sc_hd__nand3_1 _20951_ (.A(_01990_),
    .B(_01992_),
    .C(_02122_),
    .Y(_02124_));
 sky130_fd_sc_hd__and3_1 _20952_ (.A(_02110_),
    .B(_02123_),
    .C(_02124_),
    .X(_02125_));
 sky130_fd_sc_hd__inv_2 _20953_ (.A(_02125_),
    .Y(_02126_));
 sky130_fd_sc_hd__a21oi_1 _20954_ (.A1(_02123_),
    .A2(_02124_),
    .B1(_02110_),
    .Y(_02127_));
 sky130_fd_sc_hd__a211o_2 _20955_ (.A1(_01956_),
    .A2(_01959_),
    .B1(_02125_),
    .C1(_02127_),
    .X(_02128_));
 sky130_fd_sc_hd__o211ai_2 _20956_ (.A1(_02125_),
    .A2(_02127_),
    .B1(_01956_),
    .C1(_01959_),
    .Y(_02129_));
 sky130_fd_sc_hd__o211a_1 _20957_ (.A1(_01996_),
    .A2(_01998_),
    .B1(_02128_),
    .C1(_02129_),
    .X(_02130_));
 sky130_fd_sc_hd__inv_2 _20958_ (.A(_02130_),
    .Y(_02131_));
 sky130_fd_sc_hd__a211oi_2 _20959_ (.A1(_02128_),
    .A2(_02129_),
    .B1(_01996_),
    .C1(_01998_),
    .Y(_02132_));
 sky130_fd_sc_hd__or3_2 _20960_ (.A(_02093_),
    .B(_02130_),
    .C(_02132_),
    .X(_02133_));
 sky130_fd_sc_hd__o21ai_2 _20961_ (.A1(_02130_),
    .A2(_02132_),
    .B1(_02093_),
    .Y(_02134_));
 sky130_fd_sc_hd__o211ai_4 _20962_ (.A1(_01963_),
    .A2(_02004_),
    .B1(_02133_),
    .C1(_02134_),
    .Y(_02135_));
 sky130_fd_sc_hd__a211o_1 _20963_ (.A1(_02133_),
    .A2(_02134_),
    .B1(_01963_),
    .C1(_02004_),
    .X(_02136_));
 sky130_fd_sc_hd__nand2_1 _20964_ (.A(_02135_),
    .B(_02136_),
    .Y(_02137_));
 sky130_fd_sc_hd__a22o_1 _20965_ (.A1(net242),
    .A2(net72),
    .B1(net69),
    .B2(net245),
    .X(_02138_));
 sky130_fd_sc_hd__and4_1 _20966_ (.A(net245),
    .B(net242),
    .C(net72),
    .D(net69),
    .X(_02139_));
 sky130_fd_sc_hd__inv_2 _20967_ (.A(_02139_),
    .Y(_02140_));
 sky130_fd_sc_hd__a22oi_1 _20968_ (.A1(net628),
    .A2(net66),
    .B1(_02138_),
    .B2(_02140_),
    .Y(_02141_));
 sky130_fd_sc_hd__and4_1 _20969_ (.A(net629),
    .B(net66),
    .C(_02138_),
    .D(_02140_),
    .X(_02142_));
 sky130_fd_sc_hd__or2_1 _20970_ (.A(_02141_),
    .B(_02142_),
    .X(_02143_));
 sky130_fd_sc_hd__or2_1 _20971_ (.A(_02012_),
    .B(_02015_),
    .X(_02144_));
 sky130_fd_sc_hd__and2b_1 _20972_ (.A_N(_02144_),
    .B(_02143_),
    .X(_02145_));
 sky130_fd_sc_hd__and2b_1 _20973_ (.A_N(_02143_),
    .B(_02144_),
    .X(_02146_));
 sky130_fd_sc_hd__or2_1 _20974_ (.A(_02145_),
    .B(_02146_),
    .X(_02147_));
 sky130_fd_sc_hd__and4b_2 _20975_ (.A_N(net255),
    .B(net63),
    .C(\mul1.b[31] ),
    .D(net250),
    .X(_02148_));
 sky130_fd_sc_hd__o2bb2a_1 _20976_ (.A1_N(net251),
    .A2_N(net63),
    .B1(net56),
    .B2(net255),
    .X(_02149_));
 sky130_fd_sc_hd__o21a_1 _20977_ (.A1(_02148_),
    .A2(_02149_),
    .B1(_02147_),
    .X(_02150_));
 sky130_fd_sc_hd__nor3_1 _20978_ (.A(_02147_),
    .B(_02148_),
    .C(_02149_),
    .Y(_02151_));
 sky130_fd_sc_hd__nor2_1 _20979_ (.A(_02150_),
    .B(_02151_),
    .Y(_02152_));
 sky130_fd_sc_hd__o32ai_4 _20980_ (.A1(_02018_),
    .A2(_02019_),
    .A3(_02021_),
    .B1(_02017_),
    .B2(_02016_),
    .Y(_02153_));
 sky130_fd_sc_hd__xnor2_1 _20981_ (.A(_02152_),
    .B(_02153_),
    .Y(_02154_));
 sky130_fd_sc_hd__nor2_1 _20982_ (.A(_02020_),
    .B(_02154_),
    .Y(_02155_));
 sky130_fd_sc_hd__and2_1 _20983_ (.A(_02020_),
    .B(_02154_),
    .X(_02156_));
 sky130_fd_sc_hd__or2_1 _20984_ (.A(_02155_),
    .B(_02156_),
    .X(_02157_));
 sky130_fd_sc_hd__or2_1 _20985_ (.A(_02035_),
    .B(_02037_),
    .X(_02158_));
 sky130_fd_sc_hd__nand2_1 _20986_ (.A(_01966_),
    .B(_01968_),
    .Y(_02159_));
 sky130_fd_sc_hd__a22o_1 _20987_ (.A1(net226),
    .A2(net83),
    .B1(net79),
    .B2(net230),
    .X(_02160_));
 sky130_fd_sc_hd__inv_2 _20988_ (.A(_02160_),
    .Y(_02161_));
 sky130_fd_sc_hd__and4_1 _20989_ (.A(net230),
    .B(net226),
    .C(net83),
    .D(net79),
    .X(_02162_));
 sky130_fd_sc_hd__o2bb2a_1 _20990_ (.A1_N(net236),
    .A2_N(net76),
    .B1(_02161_),
    .B2(_02162_),
    .X(_02163_));
 sky130_fd_sc_hd__and4b_1 _20991_ (.A_N(_02162_),
    .B(net76),
    .C(net237),
    .D(_02160_),
    .X(_02164_));
 sky130_fd_sc_hd__or2_1 _20992_ (.A(_02163_),
    .B(_02164_),
    .X(_02165_));
 sky130_fd_sc_hd__nand2b_1 _20993_ (.A_N(_02165_),
    .B(_02159_),
    .Y(_02166_));
 sky130_fd_sc_hd__xnor2_1 _20994_ (.A(_02159_),
    .B(_02165_),
    .Y(_02167_));
 sky130_fd_sc_hd__nand2_1 _20995_ (.A(_02158_),
    .B(_02167_),
    .Y(_02168_));
 sky130_fd_sc_hd__or2_1 _20996_ (.A(_02158_),
    .B(_02167_),
    .X(_02169_));
 sky130_fd_sc_hd__nand2_1 _20997_ (.A(_02168_),
    .B(_02169_),
    .Y(_02170_));
 sky130_fd_sc_hd__a21oi_2 _20998_ (.A1(_01976_),
    .A2(_01979_),
    .B1(_02170_),
    .Y(_02171_));
 sky130_fd_sc_hd__and3_1 _20999_ (.A(_01976_),
    .B(_01979_),
    .C(_02170_),
    .X(_02172_));
 sky130_fd_sc_hd__a211oi_2 _21000_ (.A1(_02039_),
    .A2(_02041_),
    .B1(_02171_),
    .C1(_02172_),
    .Y(_02173_));
 sky130_fd_sc_hd__o211a_1 _21001_ (.A1(_02171_),
    .A2(_02172_),
    .B1(_02039_),
    .C1(_02041_),
    .X(_02174_));
 sky130_fd_sc_hd__a211oi_2 _21002_ (.A1(_02045_),
    .A2(_02047_),
    .B1(_02173_),
    .C1(_02174_),
    .Y(_02175_));
 sky130_fd_sc_hd__inv_2 _21003_ (.A(_02175_),
    .Y(_02176_));
 sky130_fd_sc_hd__o211a_1 _21004_ (.A1(_02173_),
    .A2(_02174_),
    .B1(_02045_),
    .C1(_02047_),
    .X(_02177_));
 sky130_fd_sc_hd__or3_2 _21005_ (.A(_02157_),
    .B(_02175_),
    .C(_02177_),
    .X(_02178_));
 sky130_fd_sc_hd__o21ai_1 _21006_ (.A1(_02175_),
    .A2(_02177_),
    .B1(_02157_),
    .Y(_02179_));
 sky130_fd_sc_hd__o211a_1 _21007_ (.A1(_02000_),
    .A2(_02002_),
    .B1(_02178_),
    .C1(_02179_),
    .X(_02180_));
 sky130_fd_sc_hd__inv_2 _21008_ (.A(_02180_),
    .Y(_02181_));
 sky130_fd_sc_hd__a211o_1 _21009_ (.A1(_02178_),
    .A2(_02179_),
    .B1(_02000_),
    .C1(_02002_),
    .X(_02182_));
 sky130_fd_sc_hd__o211a_1 _21010_ (.A1(_02049_),
    .A2(_02051_),
    .B1(_02181_),
    .C1(_02182_),
    .X(_02183_));
 sky130_fd_sc_hd__a211oi_1 _21011_ (.A1(_02181_),
    .A2(_02182_),
    .B1(_02049_),
    .C1(_02051_),
    .Y(_02184_));
 sky130_fd_sc_hd__or3_1 _21012_ (.A(_02137_),
    .B(_02183_),
    .C(_02184_),
    .X(_02185_));
 sky130_fd_sc_hd__o21ai_1 _21013_ (.A1(_02183_),
    .A2(_02184_),
    .B1(_02137_),
    .Y(_02186_));
 sky130_fd_sc_hd__and2_1 _21014_ (.A(_02185_),
    .B(_02186_),
    .X(_02187_));
 sky130_fd_sc_hd__o21a_1 _21015_ (.A1(_02006_),
    .A2(_02058_),
    .B1(_02187_),
    .X(_02188_));
 sky130_fd_sc_hd__nor3_1 _21016_ (.A(_02006_),
    .B(_02058_),
    .C(_02187_),
    .Y(_02189_));
 sky130_fd_sc_hd__a211oi_2 _21017_ (.A1(_02054_),
    .A2(_02056_),
    .B1(_02188_),
    .C1(_02189_),
    .Y(_02190_));
 sky130_fd_sc_hd__o211a_1 _21018_ (.A1(_02188_),
    .A2(_02189_),
    .B1(_02054_),
    .C1(_02056_),
    .X(_02191_));
 sky130_fd_sc_hd__a211oi_2 _21019_ (.A1(_02060_),
    .A2(_02062_),
    .B1(_02190_),
    .C1(_02191_),
    .Y(_02192_));
 sky130_fd_sc_hd__o211a_1 _21020_ (.A1(_02190_),
    .A2(_02191_),
    .B1(_02060_),
    .C1(_02062_),
    .X(_02193_));
 sky130_fd_sc_hd__a211oi_2 _21021_ (.A1(_02025_),
    .A2(_02028_),
    .B1(_02192_),
    .C1(_02193_),
    .Y(_02194_));
 sky130_fd_sc_hd__o211a_1 _21022_ (.A1(_02192_),
    .A2(_02193_),
    .B1(_02025_),
    .C1(_02028_),
    .X(_02195_));
 sky130_fd_sc_hd__a211oi_2 _21023_ (.A1(_02064_),
    .A2(_02068_),
    .B1(_02194_),
    .C1(_02195_),
    .Y(_02196_));
 sky130_fd_sc_hd__o211ai_2 _21024_ (.A1(_02194_),
    .A2(_02195_),
    .B1(_02064_),
    .C1(_02068_),
    .Y(_02197_));
 sky130_fd_sc_hd__and2b_1 _21025_ (.A_N(_02196_),
    .B(_02197_),
    .X(_02198_));
 sky130_fd_sc_hd__nor2_1 _21026_ (.A(_02071_),
    .B(_02079_),
    .Y(_02199_));
 sky130_fd_sc_hd__xnor2_1 _21027_ (.A(_02198_),
    .B(_02199_),
    .Y(_02200_));
 sky130_fd_sc_hd__nor2_1 _21028_ (.A(net43),
    .B(_07619_),
    .Y(_02201_));
 sky130_fd_sc_hd__a221o_1 _21029_ (.A1(net723),
    .A2(net8),
    .B1(_02200_),
    .B2(net10),
    .C1(_02201_),
    .X(_02202_));
 sky130_fd_sc_hd__mux2_1 _21030_ (.A0(net746),
    .A1(_02202_),
    .S(net1),
    .X(_00327_));
 sky130_fd_sc_hd__o21ba_1 _21031_ (.A1(_01560_),
    .A2(_02090_),
    .B1_N(_01557_),
    .X(_02203_));
 sky130_fd_sc_hd__o21ai_4 _21032_ (.A1(_01832_),
    .A2(_02084_),
    .B1(_01825_),
    .Y(_02204_));
 sky130_fd_sc_hd__xor2_2 _21033_ (.A(_02087_),
    .B(_02204_),
    .X(_02205_));
 sky130_fd_sc_hd__xnor2_1 _21034_ (.A(_01559_),
    .B(_02205_),
    .Y(_02206_));
 sky130_fd_sc_hd__xnor2_1 _21035_ (.A(_02203_),
    .B(_02206_),
    .Y(_02207_));
 sky130_fd_sc_hd__a22o_1 _21036_ (.A1(net91),
    .A2(net214),
    .B1(net210),
    .B2(net97),
    .X(_02208_));
 sky130_fd_sc_hd__and4_1 _21037_ (.A(net97),
    .B(net91),
    .C(net214),
    .D(net210),
    .X(_02209_));
 sky130_fd_sc_hd__inv_2 _21038_ (.A(_02209_),
    .Y(_02210_));
 sky130_fd_sc_hd__a22oi_1 _21039_ (.A1(net218),
    .A2(net86),
    .B1(_02208_),
    .B2(_02210_),
    .Y(_02211_));
 sky130_fd_sc_hd__and4_1 _21040_ (.A(net218),
    .B(net86),
    .C(_02208_),
    .D(_02210_),
    .X(_02212_));
 sky130_fd_sc_hd__or2_1 _21041_ (.A(_02211_),
    .B(_02212_),
    .X(_02213_));
 sky130_fd_sc_hd__a22o_1 _21042_ (.A1(\mul1.b[19] ),
    .A2(net204),
    .B1(\mul1.a[28] ),
    .B2(net112),
    .X(_02214_));
 sky130_fd_sc_hd__and4_1 _21043_ (.A(net112),
    .B(\mul1.b[19] ),
    .C(net204),
    .D(\mul1.a[28] ),
    .X(_02215_));
 sky130_fd_sc_hd__inv_2 _21044_ (.A(_02215_),
    .Y(_02216_));
 sky130_fd_sc_hd__a22oi_1 _21045_ (.A1(net98),
    .A2(\mul1.a[26] ),
    .B1(_02214_),
    .B2(_02216_),
    .Y(_02217_));
 sky130_fd_sc_hd__and4_1 _21046_ (.A(net98),
    .B(net207),
    .C(_02214_),
    .D(_02216_),
    .X(_02218_));
 sky130_fd_sc_hd__or2_1 _21047_ (.A(_02217_),
    .B(_02218_),
    .X(_02219_));
 sky130_fd_sc_hd__or2_1 _21048_ (.A(_02100_),
    .B(_02103_),
    .X(_02220_));
 sky130_fd_sc_hd__nand2b_1 _21049_ (.A_N(_02219_),
    .B(_02220_),
    .Y(_02221_));
 sky130_fd_sc_hd__xor2_1 _21050_ (.A(_02219_),
    .B(_02220_),
    .X(_02222_));
 sky130_fd_sc_hd__or2_1 _21051_ (.A(_02213_),
    .B(_02222_),
    .X(_02223_));
 sky130_fd_sc_hd__nand2_1 _21052_ (.A(_02213_),
    .B(_02222_),
    .Y(_02224_));
 sky130_fd_sc_hd__and2_1 _21053_ (.A(_02223_),
    .B(_02224_),
    .X(_02225_));
 sky130_fd_sc_hd__or2_1 _21054_ (.A(_02114_),
    .B(_02117_),
    .X(_02226_));
 sky130_fd_sc_hd__o21ba_1 _21055_ (.A1(_01949_),
    .A2(_02083_),
    .B1_N(_01948_),
    .X(_02227_));
 sky130_fd_sc_hd__and2_1 _21056_ (.A(net123),
    .B(net194),
    .X(_02228_));
 sky130_fd_sc_hd__a21oi_1 _21057_ (.A1(net118),
    .A2(net196),
    .B1(_02228_),
    .Y(_02229_));
 sky130_fd_sc_hd__and3_1 _21058_ (.A(net118),
    .B(net196),
    .C(_02228_),
    .X(_02230_));
 sky130_fd_sc_hd__or2_1 _21059_ (.A(_02229_),
    .B(_02230_),
    .X(_02231_));
 sky130_fd_sc_hd__nand2_1 _21060_ (.A(net113),
    .B(\mul1.a[29] ),
    .Y(_02232_));
 sky130_fd_sc_hd__xnor2_1 _21061_ (.A(_02231_),
    .B(_02232_),
    .Y(_02233_));
 sky130_fd_sc_hd__xor2_1 _21062_ (.A(_02227_),
    .B(_02233_),
    .X(_02234_));
 sky130_fd_sc_hd__nand2_1 _21063_ (.A(_02226_),
    .B(_02234_),
    .Y(_02235_));
 sky130_fd_sc_hd__or2_1 _21064_ (.A(_02226_),
    .B(_02234_),
    .X(_02236_));
 sky130_fd_sc_hd__nand2_1 _21065_ (.A(_02235_),
    .B(_02236_),
    .Y(_02237_));
 sky130_fd_sc_hd__a21oi_1 _21066_ (.A1(_02111_),
    .A2(_02121_),
    .B1(_02119_),
    .Y(_02238_));
 sky130_fd_sc_hd__xor2_1 _21067_ (.A(_02237_),
    .B(_02238_),
    .X(_02239_));
 sky130_fd_sc_hd__and2_1 _21068_ (.A(_02225_),
    .B(_02239_),
    .X(_02240_));
 sky130_fd_sc_hd__nor2_1 _21069_ (.A(_02225_),
    .B(_02239_),
    .Y(_02241_));
 sky130_fd_sc_hd__a211oi_2 _21070_ (.A1(_02086_),
    .A2(_02088_),
    .B1(_02240_),
    .C1(_02241_),
    .Y(_02242_));
 sky130_fd_sc_hd__o211a_1 _21071_ (.A1(_02240_),
    .A2(_02241_),
    .B1(_02086_),
    .C1(_02088_),
    .X(_02243_));
 sky130_fd_sc_hd__a211oi_2 _21072_ (.A1(_02123_),
    .A2(_02126_),
    .B1(_02242_),
    .C1(_02243_),
    .Y(_02244_));
 sky130_fd_sc_hd__o211a_1 _21073_ (.A1(_02242_),
    .A2(_02243_),
    .B1(_02123_),
    .C1(_02126_),
    .X(_02245_));
 sky130_fd_sc_hd__o21ai_1 _21074_ (.A1(_02244_),
    .A2(_02245_),
    .B1(_02207_),
    .Y(_02246_));
 sky130_fd_sc_hd__or3_1 _21075_ (.A(_02207_),
    .B(_02244_),
    .C(_02245_),
    .X(_02247_));
 sky130_fd_sc_hd__o21ai_1 _21076_ (.A1(_02091_),
    .A2(_02092_),
    .B1(_02133_),
    .Y(_02248_));
 sky130_fd_sc_hd__and3_1 _21077_ (.A(_02246_),
    .B(_02247_),
    .C(_02248_),
    .X(_02249_));
 sky130_fd_sc_hd__a21oi_1 _21078_ (.A1(_02246_),
    .A2(_02247_),
    .B1(_02248_),
    .Y(_02250_));
 sky130_fd_sc_hd__a22o_1 _21079_ (.A1(net236),
    .A2(net72),
    .B1(net69),
    .B2(net242),
    .X(_02251_));
 sky130_fd_sc_hd__and4_1 _21080_ (.A(net242),
    .B(net236),
    .C(net72),
    .D(net69),
    .X(_02252_));
 sky130_fd_sc_hd__inv_2 _21081_ (.A(_02252_),
    .Y(_02253_));
 sky130_fd_sc_hd__a22oi_1 _21082_ (.A1(net245),
    .A2(net66),
    .B1(_02251_),
    .B2(_02253_),
    .Y(_02254_));
 sky130_fd_sc_hd__and4_1 _21083_ (.A(net245),
    .B(net66),
    .C(_02251_),
    .D(_02253_),
    .X(_02255_));
 sky130_fd_sc_hd__or2_2 _21084_ (.A(_02254_),
    .B(_02255_),
    .X(_02256_));
 sky130_fd_sc_hd__nor2_2 _21085_ (.A(_02139_),
    .B(_02142_),
    .Y(_02257_));
 sky130_fd_sc_hd__xnor2_2 _21086_ (.A(_02256_),
    .B(_02257_),
    .Y(_02258_));
 sky130_fd_sc_hd__and4b_2 _21087_ (.A_N(net250),
    .B(net63),
    .C(\mul1.b[31] ),
    .D(net629),
    .X(_02259_));
 sky130_fd_sc_hd__o2bb2a_1 _21088_ (.A1_N(net629),
    .A2_N(net63),
    .B1(net56),
    .B2(net250),
    .X(_02260_));
 sky130_fd_sc_hd__nor2_1 _21089_ (.A(_02259_),
    .B(_02260_),
    .Y(_02261_));
 sky130_fd_sc_hd__xnor2_1 _21090_ (.A(_02258_),
    .B(_02261_),
    .Y(_02262_));
 sky130_fd_sc_hd__nor3_1 _21091_ (.A(_02146_),
    .B(_02151_),
    .C(_02262_),
    .Y(_02263_));
 sky130_fd_sc_hd__o21a_1 _21092_ (.A1(_02146_),
    .A2(_02151_),
    .B1(_02262_),
    .X(_02264_));
 sky130_fd_sc_hd__or2_2 _21093_ (.A(_02263_),
    .B(_02264_),
    .X(_02265_));
 sky130_fd_sc_hd__inv_2 _21094_ (.A(_02265_),
    .Y(_02266_));
 sky130_fd_sc_hd__xor2_2 _21095_ (.A(_02148_),
    .B(_02265_),
    .X(_02267_));
 sky130_fd_sc_hd__or2_1 _21096_ (.A(_02162_),
    .B(_02164_),
    .X(_02268_));
 sky130_fd_sc_hd__nand2_1 _21097_ (.A(_02095_),
    .B(_02097_),
    .Y(_02269_));
 sky130_fd_sc_hd__a22o_1 _21098_ (.A1(net223),
    .A2(net83),
    .B1(net79),
    .B2(net226),
    .X(_02270_));
 sky130_fd_sc_hd__and4_1 _21099_ (.A(net226),
    .B(net223),
    .C(net83),
    .D(net79),
    .X(_02271_));
 sky130_fd_sc_hd__inv_2 _21100_ (.A(_02271_),
    .Y(_02272_));
 sky130_fd_sc_hd__a22oi_1 _21101_ (.A1(net230),
    .A2(net76),
    .B1(_02270_),
    .B2(_02272_),
    .Y(_02273_));
 sky130_fd_sc_hd__and4_1 _21102_ (.A(net230),
    .B(net76),
    .C(_02270_),
    .D(_02272_),
    .X(_02274_));
 sky130_fd_sc_hd__or2_1 _21103_ (.A(_02273_),
    .B(_02274_),
    .X(_02275_));
 sky130_fd_sc_hd__nand2b_1 _21104_ (.A_N(_02275_),
    .B(_02269_),
    .Y(_02276_));
 sky130_fd_sc_hd__xnor2_1 _21105_ (.A(_02269_),
    .B(_02275_),
    .Y(_02277_));
 sky130_fd_sc_hd__nand2_1 _21106_ (.A(_02268_),
    .B(_02277_),
    .Y(_02278_));
 sky130_fd_sc_hd__or2_1 _21107_ (.A(_02268_),
    .B(_02277_),
    .X(_02279_));
 sky130_fd_sc_hd__nand2_1 _21108_ (.A(_02278_),
    .B(_02279_),
    .Y(_02280_));
 sky130_fd_sc_hd__a21oi_2 _21109_ (.A1(_02105_),
    .A2(_02108_),
    .B1(_02280_),
    .Y(_02281_));
 sky130_fd_sc_hd__and3_1 _21110_ (.A(_02105_),
    .B(_02108_),
    .C(_02280_),
    .X(_02282_));
 sky130_fd_sc_hd__a211oi_1 _21111_ (.A1(_02166_),
    .A2(_02168_),
    .B1(_02281_),
    .C1(_02282_),
    .Y(_02283_));
 sky130_fd_sc_hd__a211o_1 _21112_ (.A1(_02166_),
    .A2(_02168_),
    .B1(_02281_),
    .C1(_02282_),
    .X(_02284_));
 sky130_fd_sc_hd__o211ai_1 _21113_ (.A1(_02281_),
    .A2(_02282_),
    .B1(_02166_),
    .C1(_02168_),
    .Y(_02285_));
 sky130_fd_sc_hd__o211a_1 _21114_ (.A1(_02171_),
    .A2(_02173_),
    .B1(_02284_),
    .C1(_02285_),
    .X(_02286_));
 sky130_fd_sc_hd__a211oi_1 _21115_ (.A1(_02284_),
    .A2(_02285_),
    .B1(_02171_),
    .C1(_02173_),
    .Y(_02287_));
 sky130_fd_sc_hd__nor3_1 _21116_ (.A(_02267_),
    .B(_02286_),
    .C(_02287_),
    .Y(_02288_));
 sky130_fd_sc_hd__o21a_1 _21117_ (.A1(_02286_),
    .A2(_02287_),
    .B1(_02267_),
    .X(_02289_));
 sky130_fd_sc_hd__a211oi_2 _21118_ (.A1(_02128_),
    .A2(_02131_),
    .B1(_02288_),
    .C1(_02289_),
    .Y(_02290_));
 sky130_fd_sc_hd__o211a_1 _21119_ (.A1(_02288_),
    .A2(_02289_),
    .B1(_02128_),
    .C1(_02131_),
    .X(_02291_));
 sky130_fd_sc_hd__a211oi_2 _21120_ (.A1(_02176_),
    .A2(_02178_),
    .B1(_02290_),
    .C1(_02291_),
    .Y(_02292_));
 sky130_fd_sc_hd__o211a_1 _21121_ (.A1(_02290_),
    .A2(_02291_),
    .B1(_02176_),
    .C1(_02178_),
    .X(_02293_));
 sky130_fd_sc_hd__nor4_1 _21122_ (.A(_02249_),
    .B(_02250_),
    .C(_02292_),
    .D(_02293_),
    .Y(_02294_));
 sky130_fd_sc_hd__o22a_1 _21123_ (.A1(_02249_),
    .A2(_02250_),
    .B1(_02292_),
    .B2(_02293_),
    .X(_02295_));
 sky130_fd_sc_hd__a211o_1 _21124_ (.A1(_02135_),
    .A2(_02185_),
    .B1(_02294_),
    .C1(_02295_),
    .X(_02296_));
 sky130_fd_sc_hd__o211ai_2 _21125_ (.A1(_02294_),
    .A2(_02295_),
    .B1(_02135_),
    .C1(_02185_),
    .Y(_02297_));
 sky130_fd_sc_hd__o211ai_2 _21126_ (.A1(_02180_),
    .A2(_02183_),
    .B1(_02296_),
    .C1(_02297_),
    .Y(_02298_));
 sky130_fd_sc_hd__a211o_1 _21127_ (.A1(_02296_),
    .A2(_02297_),
    .B1(_02180_),
    .C1(_02183_),
    .X(_02299_));
 sky130_fd_sc_hd__nand2_1 _21128_ (.A(_02298_),
    .B(_02299_),
    .Y(_02300_));
 sky130_fd_sc_hd__or2_1 _21129_ (.A(_02188_),
    .B(_02190_),
    .X(_02301_));
 sky130_fd_sc_hd__and3_1 _21130_ (.A(_02298_),
    .B(_02299_),
    .C(_02301_),
    .X(_02302_));
 sky130_fd_sc_hd__xnor2_1 _21131_ (.A(_02300_),
    .B(_02301_),
    .Y(_02303_));
 sky130_fd_sc_hd__a21oi_1 _21132_ (.A1(_02152_),
    .A2(_02153_),
    .B1(_02155_),
    .Y(_02304_));
 sky130_fd_sc_hd__and2b_1 _21133_ (.A_N(_02304_),
    .B(_02303_),
    .X(_02305_));
 sky130_fd_sc_hd__xor2_1 _21134_ (.A(_02303_),
    .B(_02304_),
    .X(_02306_));
 sky130_fd_sc_hd__or2_1 _21135_ (.A(_02192_),
    .B(_02194_),
    .X(_02307_));
 sky130_fd_sc_hd__and2b_1 _21136_ (.A_N(_02306_),
    .B(_02307_),
    .X(_02308_));
 sky130_fd_sc_hd__xnor2_1 _21137_ (.A(_02306_),
    .B(_02307_),
    .Y(_02309_));
 sky130_fd_sc_hd__or2_1 _21138_ (.A(_02071_),
    .B(_02196_),
    .X(_02310_));
 sky130_fd_sc_hd__a221oi_1 _21139_ (.A1(_02079_),
    .A2(_02198_),
    .B1(_02310_),
    .B2(_02197_),
    .C1(_02309_),
    .Y(_02311_));
 sky130_fd_sc_hd__o311a_1 _21140_ (.A1(_02071_),
    .A2(_02079_),
    .A3(_02196_),
    .B1(_02197_),
    .C1(_02309_),
    .X(_02312_));
 sky130_fd_sc_hd__nor2_1 _21141_ (.A(_02311_),
    .B(_02312_),
    .Y(_02313_));
 sky130_fd_sc_hd__nor2_1 _21142_ (.A(net43),
    .B(_07730_),
    .Y(_02314_));
 sky130_fd_sc_hd__a221o_1 _21143_ (.A1(\temp[29] ),
    .A2(net8),
    .B1(_02313_),
    .B2(net10),
    .C1(_02314_),
    .X(_02315_));
 sky130_fd_sc_hd__mux2_1 _21144_ (.A0(net792),
    .A1(_02315_),
    .S(net1),
    .X(_00328_));
 sky130_fd_sc_hd__o21ai_1 _21145_ (.A1(_02203_),
    .A2(_02206_),
    .B1(_02247_),
    .Y(_02316_));
 sky130_fd_sc_hd__and2b_1 _21146_ (.A_N(_02205_),
    .B(_01558_),
    .X(_02317_));
 sky130_fd_sc_hd__a21o_1 _21147_ (.A1(_01557_),
    .A2(_02205_),
    .B1(_02317_),
    .X(_02318_));
 sky130_fd_sc_hd__o21ba_1 _21148_ (.A1(_02237_),
    .A2(_02238_),
    .B1_N(_02240_),
    .X(_02319_));
 sky130_fd_sc_hd__a21boi_4 _21149_ (.A1(_02087_),
    .A2(_02204_),
    .B1_N(_02086_),
    .Y(_02320_));
 sky130_fd_sc_hd__a22o_1 _21150_ (.A1(net91),
    .A2(net210),
    .B1(net207),
    .B2(net97),
    .X(_02321_));
 sky130_fd_sc_hd__and3_1 _21151_ (.A(net97),
    .B(net91),
    .C(\mul1.a[25] ),
    .X(_02322_));
 sky130_fd_sc_hd__a21bo_1 _21152_ (.A1(net207),
    .A2(_02322_),
    .B1_N(_02321_),
    .X(_02323_));
 sky130_fd_sc_hd__nand2_1 _21153_ (.A(net86),
    .B(net213),
    .Y(_02324_));
 sky130_fd_sc_hd__xnor2_1 _21154_ (.A(_02323_),
    .B(_02324_),
    .Y(_02325_));
 sky130_fd_sc_hd__a22o_1 _21155_ (.A1(\mul1.b[19] ),
    .A2(net201),
    .B1(net198),
    .B2(net112),
    .X(_02326_));
 sky130_fd_sc_hd__and3_1 _21156_ (.A(net112),
    .B(\mul1.b[19] ),
    .C(net201),
    .X(_02327_));
 sky130_fd_sc_hd__a21bo_1 _21157_ (.A1(net198),
    .A2(_02327_),
    .B1_N(_02326_),
    .X(_02328_));
 sky130_fd_sc_hd__nand2_1 _21158_ (.A(net98),
    .B(net204),
    .Y(_02329_));
 sky130_fd_sc_hd__xnor2_1 _21159_ (.A(_02328_),
    .B(_02329_),
    .Y(_02330_));
 sky130_fd_sc_hd__o21bai_1 _21160_ (.A1(_02215_),
    .A2(_02218_),
    .B1_N(_02330_),
    .Y(_02331_));
 sky130_fd_sc_hd__or3b_1 _21161_ (.A(_02215_),
    .B(_02218_),
    .C_N(_02330_),
    .X(_02332_));
 sky130_fd_sc_hd__nand2_1 _21162_ (.A(_02331_),
    .B(_02332_),
    .Y(_02333_));
 sky130_fd_sc_hd__xor2_1 _21163_ (.A(_02325_),
    .B(_02333_),
    .X(_02334_));
 sky130_fd_sc_hd__inv_2 _21164_ (.A(_02334_),
    .Y(_02335_));
 sky130_fd_sc_hd__o21ai_1 _21165_ (.A1(_02227_),
    .A2(_02233_),
    .B1(_02235_),
    .Y(_02336_));
 sky130_fd_sc_hd__o21ba_1 _21166_ (.A1(_02229_),
    .A2(_02232_),
    .B1_N(_02230_),
    .X(_02337_));
 sky130_fd_sc_hd__o21ai_1 _21167_ (.A1(net123),
    .A2(net118),
    .B1(net194),
    .Y(_02338_));
 sky130_fd_sc_hd__inv_2 _21168_ (.A(_02338_),
    .Y(_02339_));
 sky130_fd_sc_hd__nand2_1 _21169_ (.A(net118),
    .B(_02228_),
    .Y(_02340_));
 sky130_fd_sc_hd__a22o_1 _21170_ (.A1(net113),
    .A2(net196),
    .B1(_02339_),
    .B2(_02340_),
    .X(_02341_));
 sky130_fd_sc_hd__nand4_1 _21171_ (.A(net113),
    .B(net196),
    .C(_02339_),
    .D(_02340_),
    .Y(_02342_));
 sky130_fd_sc_hd__and3_1 _21172_ (.A(_02227_),
    .B(_02341_),
    .C(_02342_),
    .X(_02343_));
 sky130_fd_sc_hd__a21oi_1 _21173_ (.A1(_02341_),
    .A2(_02342_),
    .B1(_02227_),
    .Y(_02344_));
 sky130_fd_sc_hd__nor2_1 _21174_ (.A(_02343_),
    .B(_02344_),
    .Y(_02345_));
 sky130_fd_sc_hd__xor2_1 _21175_ (.A(_02337_),
    .B(_02345_),
    .X(_02346_));
 sky130_fd_sc_hd__xnor2_1 _21176_ (.A(_02336_),
    .B(_02346_),
    .Y(_02347_));
 sky130_fd_sc_hd__nor2_1 _21177_ (.A(_02335_),
    .B(_02347_),
    .Y(_02348_));
 sky130_fd_sc_hd__and2_1 _21178_ (.A(_02335_),
    .B(_02347_),
    .X(_02349_));
 sky130_fd_sc_hd__nor2_1 _21179_ (.A(_02348_),
    .B(_02349_),
    .Y(_02350_));
 sky130_fd_sc_hd__xnor2_1 _21180_ (.A(_02320_),
    .B(_02350_),
    .Y(_02351_));
 sky130_fd_sc_hd__nand2b_1 _21181_ (.A_N(_02319_),
    .B(_02351_),
    .Y(_02352_));
 sky130_fd_sc_hd__xnor2_1 _21182_ (.A(_02319_),
    .B(_02351_),
    .Y(_02353_));
 sky130_fd_sc_hd__xnor2_1 _21183_ (.A(_02318_),
    .B(_02353_),
    .Y(_02354_));
 sky130_fd_sc_hd__nand2_1 _21184_ (.A(_02316_),
    .B(_02354_),
    .Y(_02355_));
 sky130_fd_sc_hd__or2_1 _21185_ (.A(_02316_),
    .B(_02354_),
    .X(_02356_));
 sky130_fd_sc_hd__and2_1 _21186_ (.A(_02355_),
    .B(_02356_),
    .X(_02357_));
 sky130_fd_sc_hd__inv_2 _21187_ (.A(_02357_),
    .Y(_02358_));
 sky130_fd_sc_hd__or2_2 _21188_ (.A(_02286_),
    .B(_02288_),
    .X(_02359_));
 sky130_fd_sc_hd__a22oi_1 _21189_ (.A1(net230),
    .A2(net72),
    .B1(net69),
    .B2(net236),
    .Y(_02360_));
 sky130_fd_sc_hd__and4_1 _21190_ (.A(net236),
    .B(net230),
    .C(net72),
    .D(net69),
    .X(_02361_));
 sky130_fd_sc_hd__nor2_1 _21191_ (.A(_02360_),
    .B(_02361_),
    .Y(_02362_));
 sky130_fd_sc_hd__nand2_1 _21192_ (.A(net242),
    .B(net66),
    .Y(_02363_));
 sky130_fd_sc_hd__xor2_1 _21193_ (.A(_02362_),
    .B(_02363_),
    .X(_02364_));
 sky130_fd_sc_hd__or2_1 _21194_ (.A(_02252_),
    .B(_02255_),
    .X(_02365_));
 sky130_fd_sc_hd__and2b_1 _21195_ (.A_N(_02365_),
    .B(_02364_),
    .X(_02366_));
 sky130_fd_sc_hd__and2b_1 _21196_ (.A_N(_02364_),
    .B(_02365_),
    .X(_02367_));
 sky130_fd_sc_hd__nor2_1 _21197_ (.A(_02366_),
    .B(_02367_),
    .Y(_02368_));
 sky130_fd_sc_hd__a22o_1 _21198_ (.A1(net245),
    .A2(net63),
    .B1(\mul1.b[31] ),
    .B2(_02565_),
    .X(_02369_));
 sky130_fd_sc_hd__nand4_2 _21199_ (.A(net245),
    .B(_02565_),
    .C(net63),
    .D(\mul1.b[31] ),
    .Y(_02370_));
 sky130_fd_sc_hd__nand2_1 _21200_ (.A(_02369_),
    .B(_02370_),
    .Y(_02371_));
 sky130_fd_sc_hd__xnor2_2 _21201_ (.A(_02368_),
    .B(_02371_),
    .Y(_02372_));
 sky130_fd_sc_hd__o32ai_4 _21202_ (.A1(_02258_),
    .A2(_02259_),
    .A3(_02260_),
    .B1(_02257_),
    .B2(_02256_),
    .Y(_02373_));
 sky130_fd_sc_hd__and2_1 _21203_ (.A(_02372_),
    .B(_02373_),
    .X(_02374_));
 sky130_fd_sc_hd__xnor2_2 _21204_ (.A(_02372_),
    .B(_02373_),
    .Y(_02375_));
 sky130_fd_sc_hd__inv_2 _21205_ (.A(_02375_),
    .Y(_02376_));
 sky130_fd_sc_hd__xor2_2 _21206_ (.A(_02259_),
    .B(_02375_),
    .X(_02377_));
 sky130_fd_sc_hd__nand2_1 _21207_ (.A(_02221_),
    .B(_02223_),
    .Y(_02378_));
 sky130_fd_sc_hd__or2_1 _21208_ (.A(_02271_),
    .B(_02274_),
    .X(_02379_));
 sky130_fd_sc_hd__nor2_1 _21209_ (.A(_02209_),
    .B(_02212_),
    .Y(_02380_));
 sky130_fd_sc_hd__a22oi_1 _21210_ (.A1(net217),
    .A2(net83),
    .B1(net79),
    .B2(net223),
    .Y(_02381_));
 sky130_fd_sc_hd__and4_1 _21211_ (.A(net223),
    .B(net217),
    .C(net83),
    .D(net79),
    .X(_02382_));
 sky130_fd_sc_hd__nor2_1 _21212_ (.A(_02381_),
    .B(_02382_),
    .Y(_02383_));
 sky130_fd_sc_hd__nand2_1 _21213_ (.A(net226),
    .B(net76),
    .Y(_02384_));
 sky130_fd_sc_hd__xor2_1 _21214_ (.A(_02383_),
    .B(_02384_),
    .X(_02385_));
 sky130_fd_sc_hd__nor2_1 _21215_ (.A(_02380_),
    .B(_02385_),
    .Y(_02386_));
 sky130_fd_sc_hd__nand2_1 _21216_ (.A(_02380_),
    .B(_02385_),
    .Y(_02387_));
 sky130_fd_sc_hd__and2b_1 _21217_ (.A_N(_02386_),
    .B(_02387_),
    .X(_02388_));
 sky130_fd_sc_hd__xnor2_1 _21218_ (.A(_02379_),
    .B(_02388_),
    .Y(_02389_));
 sky130_fd_sc_hd__nand2b_1 _21219_ (.A_N(_02389_),
    .B(_02378_),
    .Y(_02390_));
 sky130_fd_sc_hd__xor2_1 _21220_ (.A(_02378_),
    .B(_02389_),
    .X(_02391_));
 sky130_fd_sc_hd__a21o_1 _21221_ (.A1(_02276_),
    .A2(_02278_),
    .B1(_02391_),
    .X(_02392_));
 sky130_fd_sc_hd__nand3_1 _21222_ (.A(_02276_),
    .B(_02278_),
    .C(_02391_),
    .Y(_02393_));
 sky130_fd_sc_hd__o211a_1 _21223_ (.A1(_02281_),
    .A2(_02283_),
    .B1(_02392_),
    .C1(_02393_),
    .X(_02394_));
 sky130_fd_sc_hd__a211oi_1 _21224_ (.A1(_02392_),
    .A2(_02393_),
    .B1(_02281_),
    .C1(_02283_),
    .Y(_02395_));
 sky130_fd_sc_hd__nor2_1 _21225_ (.A(_02394_),
    .B(_02395_),
    .Y(_02396_));
 sky130_fd_sc_hd__xnor2_2 _21226_ (.A(_02377_),
    .B(_02396_),
    .Y(_02397_));
 sky130_fd_sc_hd__o21a_1 _21227_ (.A1(_02242_),
    .A2(_02244_),
    .B1(_02397_),
    .X(_02398_));
 sky130_fd_sc_hd__nor3_1 _21228_ (.A(_02242_),
    .B(_02244_),
    .C(_02397_),
    .Y(_02399_));
 sky130_fd_sc_hd__nor2_1 _21229_ (.A(_02398_),
    .B(_02399_),
    .Y(_02400_));
 sky130_fd_sc_hd__xnor2_2 _21230_ (.A(_02359_),
    .B(_02400_),
    .Y(_02401_));
 sky130_fd_sc_hd__xor2_2 _21231_ (.A(_02357_),
    .B(_02401_),
    .X(_02402_));
 sky130_fd_sc_hd__or2_1 _21232_ (.A(_02249_),
    .B(_02294_),
    .X(_02403_));
 sky130_fd_sc_hd__nand2b_1 _21233_ (.A_N(_02402_),
    .B(_02403_),
    .Y(_02404_));
 sky130_fd_sc_hd__xnor2_1 _21234_ (.A(_02402_),
    .B(_02403_),
    .Y(_02405_));
 sky130_fd_sc_hd__o21ai_1 _21235_ (.A1(_02290_),
    .A2(_02292_),
    .B1(_02405_),
    .Y(_02406_));
 sky130_fd_sc_hd__or3_1 _21236_ (.A(_02290_),
    .B(_02292_),
    .C(_02405_),
    .X(_02407_));
 sky130_fd_sc_hd__nand2_1 _21237_ (.A(_02406_),
    .B(_02407_),
    .Y(_02408_));
 sky130_fd_sc_hd__and2_1 _21238_ (.A(_02296_),
    .B(_02298_),
    .X(_02409_));
 sky130_fd_sc_hd__nor2_1 _21239_ (.A(_02408_),
    .B(_02409_),
    .Y(_02410_));
 sky130_fd_sc_hd__nand2_1 _21240_ (.A(_02408_),
    .B(_02409_),
    .Y(_02411_));
 sky130_fd_sc_hd__and2b_1 _21241_ (.A_N(_02410_),
    .B(_02411_),
    .X(_02412_));
 sky130_fd_sc_hd__a21o_1 _21242_ (.A1(_02148_),
    .A2(_02266_),
    .B1(_02264_),
    .X(_02413_));
 sky130_fd_sc_hd__xor2_1 _21243_ (.A(_02412_),
    .B(_02413_),
    .X(_02414_));
 sky130_fd_sc_hd__nor3_1 _21244_ (.A(_02302_),
    .B(_02305_),
    .C(_02414_),
    .Y(_02415_));
 sky130_fd_sc_hd__o21a_1 _21245_ (.A1(_02302_),
    .A2(_02305_),
    .B1(_02414_),
    .X(_02416_));
 sky130_fd_sc_hd__nor2_1 _21246_ (.A(_02415_),
    .B(_02416_),
    .Y(_02417_));
 sky130_fd_sc_hd__nor2_1 _21247_ (.A(_02308_),
    .B(_02312_),
    .Y(_02418_));
 sky130_fd_sc_hd__xnor2_1 _21248_ (.A(_02417_),
    .B(_02418_),
    .Y(_02419_));
 sky130_fd_sc_hd__a21o_1 _21249_ (.A1(_03052_),
    .A2(_07835_),
    .B1(net8),
    .X(_02420_));
 sky130_fd_sc_hd__a21o_1 _21250_ (.A1(net10),
    .A2(_02419_),
    .B1(_02420_),
    .X(_02421_));
 sky130_fd_sc_hd__o21a_1 _21251_ (.A1(\temp[30] ),
    .A2(_03054_),
    .B1(net1),
    .X(_02422_));
 sky130_fd_sc_hd__a22o_1 _21252_ (.A1(net817),
    .A2(_03056_),
    .B1(_02421_),
    .B2(_02422_),
    .X(_00329_));
 sky130_fd_sc_hd__and2b_1 _21253_ (.A_N(_02415_),
    .B(_02308_),
    .X(_02423_));
 sky130_fd_sc_hd__a211o_1 _21254_ (.A1(_02312_),
    .A2(_02417_),
    .B1(_02423_),
    .C1(_02416_),
    .X(_02424_));
 sky130_fd_sc_hd__nand2_1 _21255_ (.A(_02404_),
    .B(_02406_),
    .Y(_02425_));
 sky130_fd_sc_hd__nand2_1 _21256_ (.A(net98),
    .B(net201),
    .Y(_02426_));
 sky130_fd_sc_hd__xnor2_1 _21257_ (.A(_02425_),
    .B(_02426_),
    .Y(_02427_));
 sky130_fd_sc_hd__nand2_1 _21258_ (.A(net102),
    .B(net198),
    .Y(_02428_));
 sky130_fd_sc_hd__xnor2_2 _21259_ (.A(_02320_),
    .B(_02428_),
    .Y(_02429_));
 sky130_fd_sc_hd__xnor2_1 _21260_ (.A(_02427_),
    .B(_02429_),
    .Y(_02430_));
 sky130_fd_sc_hd__or2_1 _21261_ (.A(net246),
    .B(net56),
    .X(_02431_));
 sky130_fd_sc_hd__a21oi_1 _21262_ (.A1(_02379_),
    .A2(_02387_),
    .B1(_02386_),
    .Y(_02432_));
 sky130_fd_sc_hd__xnor2_1 _21263_ (.A(_02431_),
    .B(_02432_),
    .Y(_02433_));
 sky130_fd_sc_hd__nand2_1 _21264_ (.A(net86),
    .B(net210),
    .Y(_02434_));
 sky130_fd_sc_hd__xnor2_1 _21265_ (.A(_02433_),
    .B(_02434_),
    .Y(_02435_));
 sky130_fd_sc_hd__xnor2_1 _21266_ (.A(_02430_),
    .B(_02435_),
    .Y(_02436_));
 sky130_fd_sc_hd__nand2_1 _21267_ (.A(net112),
    .B(\mul1.a[30] ),
    .Y(_02437_));
 sky130_fd_sc_hd__o21a_1 _21268_ (.A1(_02358_),
    .A2(_02401_),
    .B1(_02355_),
    .X(_02438_));
 sky130_fd_sc_hd__xnor2_1 _21269_ (.A(_02437_),
    .B(_02438_),
    .Y(_02439_));
 sky130_fd_sc_hd__mux2_1 _21270_ (.A0(_02343_),
    .A1(_02344_),
    .S(_02337_),
    .X(_02440_));
 sky130_fd_sc_hd__xnor2_2 _21271_ (.A(_02439_),
    .B(_02440_),
    .Y(_02441_));
 sky130_fd_sc_hd__a21o_1 _21272_ (.A1(_02411_),
    .A2(_02413_),
    .B1(_02410_),
    .X(_02442_));
 sky130_fd_sc_hd__a32o_1 _21273_ (.A1(net98),
    .A2(net204),
    .A3(_02326_),
    .B1(_02327_),
    .B2(net198),
    .X(_02443_));
 sky130_fd_sc_hd__xnor2_1 _21274_ (.A(_02442_),
    .B(_02443_),
    .Y(_02444_));
 sky130_fd_sc_hd__nand2_1 _21275_ (.A(_02390_),
    .B(_02392_),
    .Y(_02445_));
 sky130_fd_sc_hd__a21oi_1 _21276_ (.A1(_02259_),
    .A2(_02376_),
    .B1(_02374_),
    .Y(_02446_));
 sky130_fd_sc_hd__xnor2_1 _21277_ (.A(_02445_),
    .B(_02446_),
    .Y(_02447_));
 sky130_fd_sc_hd__nand2_1 _21278_ (.A(net95),
    .B(net204),
    .Y(_02448_));
 sky130_fd_sc_hd__xnor2_1 _21279_ (.A(_02447_),
    .B(_02448_),
    .Y(_02449_));
 sky130_fd_sc_hd__xnor2_1 _21280_ (.A(_02444_),
    .B(_02449_),
    .Y(_02450_));
 sky130_fd_sc_hd__xnor2_1 _21281_ (.A(_02441_),
    .B(_02450_),
    .Y(_02451_));
 sky130_fd_sc_hd__a31o_1 _21282_ (.A1(_02368_),
    .A2(_02369_),
    .A3(_02370_),
    .B1(_02367_),
    .X(_02452_));
 sky130_fd_sc_hd__nand2_1 _21283_ (.A(net214),
    .B(net83),
    .Y(_02453_));
 sky130_fd_sc_hd__o21ba_1 _21284_ (.A1(_02377_),
    .A2(_02395_),
    .B1_N(_02394_),
    .X(_02454_));
 sky130_fd_sc_hd__xnor2_1 _21285_ (.A(_02453_),
    .B(_02454_),
    .Y(_02455_));
 sky130_fd_sc_hd__nand2_1 _21286_ (.A(net226),
    .B(net72),
    .Y(_02456_));
 sky130_fd_sc_hd__xor2_1 _21287_ (.A(_02370_),
    .B(_02456_),
    .X(_02457_));
 sky130_fd_sc_hd__a32o_1 _21288_ (.A1(net86),
    .A2(net214),
    .A3(_02321_),
    .B1(_02322_),
    .B2(net207),
    .X(_02458_));
 sky130_fd_sc_hd__a31o_1 _21289_ (.A1(net242),
    .A2(net66),
    .A3(_02362_),
    .B1(_02361_),
    .X(_02459_));
 sky130_fd_sc_hd__xnor2_1 _21290_ (.A(_02458_),
    .B(_02459_),
    .Y(_02460_));
 sky130_fd_sc_hd__nand2_1 _21291_ (.A(net236),
    .B(net66),
    .Y(_02461_));
 sky130_fd_sc_hd__o31a_1 _21292_ (.A1(_02320_),
    .A2(_02348_),
    .A3(_02349_),
    .B1(_02352_),
    .X(_02462_));
 sky130_fd_sc_hd__nand2_1 _21293_ (.A(net242),
    .B(net63),
    .Y(_02463_));
 sky130_fd_sc_hd__xnor2_1 _21294_ (.A(_02462_),
    .B(_02463_),
    .Y(_02464_));
 sky130_fd_sc_hd__xnor2_1 _21295_ (.A(_02461_),
    .B(_02464_),
    .Y(_02465_));
 sky130_fd_sc_hd__nand2_1 _21296_ (.A(net230),
    .B(net69),
    .Y(_02466_));
 sky130_fd_sc_hd__xnor2_1 _21297_ (.A(_02465_),
    .B(_02466_),
    .Y(_02467_));
 sky130_fd_sc_hd__xnor2_1 _21298_ (.A(_02460_),
    .B(_02467_),
    .Y(_02468_));
 sky130_fd_sc_hd__xnor2_1 _21299_ (.A(_02457_),
    .B(_02468_),
    .Y(_02469_));
 sky130_fd_sc_hd__xnor2_1 _21300_ (.A(_02455_),
    .B(_02469_),
    .Y(_02470_));
 sky130_fd_sc_hd__nand2_1 _21301_ (.A(net91),
    .B(\mul1.a[26] ),
    .Y(_02471_));
 sky130_fd_sc_hd__a2bb2o_1 _21302_ (.A1_N(_02317_),
    .A2_N(_02353_),
    .B1(_01557_),
    .B2(_02205_),
    .X(_02472_));
 sky130_fd_sc_hd__xnor2_1 _21303_ (.A(_02471_),
    .B(_02472_),
    .Y(_02473_));
 sky130_fd_sc_hd__a31o_1 _21304_ (.A1(net226),
    .A2(net76),
    .A3(_02383_),
    .B1(_02382_),
    .X(_02474_));
 sky130_fd_sc_hd__nand2_1 _21305_ (.A(net217),
    .B(net79),
    .Y(_02475_));
 sky130_fd_sc_hd__o21a_1 _21306_ (.A1(_02325_),
    .A2(_02333_),
    .B1(_02331_),
    .X(_02476_));
 sky130_fd_sc_hd__xnor2_1 _21307_ (.A(_02475_),
    .B(_02476_),
    .Y(_02477_));
 sky130_fd_sc_hd__xnor2_1 _21308_ (.A(_02474_),
    .B(_02477_),
    .Y(_02478_));
 sky130_fd_sc_hd__xnor2_1 _21309_ (.A(_02473_),
    .B(_02478_),
    .Y(_02479_));
 sky130_fd_sc_hd__xnor2_1 _21310_ (.A(_02470_),
    .B(_02479_),
    .Y(_02480_));
 sky130_fd_sc_hd__nand2_1 _21311_ (.A(net223),
    .B(net76),
    .Y(_02481_));
 sky130_fd_sc_hd__a21o_1 _21312_ (.A1(_02359_),
    .A2(_02400_),
    .B1(_02398_),
    .X(_02482_));
 sky130_fd_sc_hd__a21oi_1 _21313_ (.A1(_02336_),
    .A2(_02346_),
    .B1(_02348_),
    .Y(_02483_));
 sky130_fd_sc_hd__o2111a_1 _21314_ (.A1(\mul1.a[30] ),
    .A2(_02338_),
    .B1(_02340_),
    .C1(net194),
    .D1(net113),
    .X(_02484_));
 sky130_fd_sc_hd__o211a_1 _21315_ (.A1(net123),
    .A2(net118),
    .B1(_02566_),
    .C1(net194),
    .X(_02485_));
 sky130_fd_sc_hd__nor2_1 _21316_ (.A(_02484_),
    .B(_02485_),
    .Y(_02486_));
 sky130_fd_sc_hd__xnor2_2 _21317_ (.A(_02483_),
    .B(_02486_),
    .Y(_02487_));
 sky130_fd_sc_hd__xnor2_2 _21318_ (.A(_02482_),
    .B(_02487_),
    .Y(_02488_));
 sky130_fd_sc_hd__xnor2_1 _21319_ (.A(_02481_),
    .B(_02488_),
    .Y(_02489_));
 sky130_fd_sc_hd__xnor2_1 _21320_ (.A(_02480_),
    .B(_02489_),
    .Y(_02490_));
 sky130_fd_sc_hd__xnor2_1 _21321_ (.A(_02452_),
    .B(_02490_),
    .Y(_02491_));
 sky130_fd_sc_hd__xnor2_1 _21322_ (.A(_02451_),
    .B(_02491_),
    .Y(_02492_));
 sky130_fd_sc_hd__xnor2_1 _21323_ (.A(_02436_),
    .B(_02492_),
    .Y(_02493_));
 sky130_fd_sc_hd__xnor2_1 _21324_ (.A(_02424_),
    .B(_02493_),
    .Y(_02494_));
 sky130_fd_sc_hd__a21o_1 _21325_ (.A1(_03052_),
    .A2(_07909_),
    .B1(net8),
    .X(_02495_));
 sky130_fd_sc_hd__a21o_1 _21326_ (.A1(net10),
    .A2(_02494_),
    .B1(_02495_),
    .X(_02496_));
 sky130_fd_sc_hd__o21a_1 _21327_ (.A1(net833),
    .A2(_03054_),
    .B1(net1),
    .X(_02497_));
 sky130_fd_sc_hd__a22o_1 _21328_ (.A1(net767),
    .A2(_03056_),
    .B1(_02496_),
    .B2(_02497_),
    .X(_00330_));
 sky130_fd_sc_hd__o21a_1 _21329_ (.A1(net595),
    .A2(net592),
    .B1(net645),
    .X(_02498_));
 sky130_fd_sc_hd__o21ai_4 _21330_ (.A1(net597),
    .A2(net592),
    .B1(net638),
    .Y(_02499_));
 sky130_fd_sc_hd__nor2_1 _21331_ (.A(net597),
    .B(_08642_),
    .Y(_02500_));
 sky130_fd_sc_hd__o21ai_1 _21332_ (.A1(net61),
    .A2(_03792_),
    .B1(net41),
    .Y(_02501_));
 sky130_fd_sc_hd__o22a_1 _21333_ (.A1(net802),
    .A2(net41),
    .B1(_02500_),
    .B2(_02501_),
    .X(_00331_));
 sky130_fd_sc_hd__nand2_1 _21334_ (.A(net61),
    .B(_08741_),
    .Y(_02502_));
 sky130_fd_sc_hd__a21oi_1 _21335_ (.A1(net597),
    .A2(_03893_),
    .B1(net39),
    .Y(_02503_));
 sky130_fd_sc_hd__a22o_1 _21336_ (.A1(net778),
    .A2(net39),
    .B1(_02502_),
    .B2(_02503_),
    .X(_00332_));
 sky130_fd_sc_hd__nor2_1 _21337_ (.A(net597),
    .B(_08843_),
    .Y(_02504_));
 sky130_fd_sc_hd__o21ai_1 _21338_ (.A1(net61),
    .A2(_03993_),
    .B1(net41),
    .Y(_02505_));
 sky130_fd_sc_hd__o22a_1 _21339_ (.A1(net839),
    .A2(net41),
    .B1(_02504_),
    .B2(_02505_),
    .X(_00333_));
 sky130_fd_sc_hd__nand2_1 _21340_ (.A(net597),
    .B(_04100_),
    .Y(_02506_));
 sky130_fd_sc_hd__o211a_1 _21341_ (.A1(net597),
    .A2(_08952_),
    .B1(net41),
    .C1(_02506_),
    .X(_02507_));
 sky130_fd_sc_hd__a21o_1 _21342_ (.A1(net771),
    .A2(net39),
    .B1(_02507_),
    .X(_00334_));
 sky130_fd_sc_hd__nand2_1 _21343_ (.A(net597),
    .B(_04209_),
    .Y(_02508_));
 sky130_fd_sc_hd__o211a_1 _21344_ (.A1(net597),
    .A2(_09062_),
    .B1(net41),
    .C1(_02508_),
    .X(_02509_));
 sky130_fd_sc_hd__a21o_1 _21345_ (.A1(net706),
    .A2(net39),
    .B1(_02509_),
    .X(_00335_));
 sky130_fd_sc_hd__or2_1 _21346_ (.A(net597),
    .B(_09176_),
    .X(_02510_));
 sky130_fd_sc_hd__a21oi_1 _21347_ (.A1(net597),
    .A2(_04325_),
    .B1(net39),
    .Y(_02511_));
 sky130_fd_sc_hd__a22o_1 _21348_ (.A1(net809),
    .A2(net39),
    .B1(_02510_),
    .B2(_02511_),
    .X(_00336_));
 sky130_fd_sc_hd__nor2_1 _21349_ (.A(net597),
    .B(_09297_),
    .Y(_02512_));
 sky130_fd_sc_hd__o21ai_1 _21350_ (.A1(net61),
    .A2(_04449_),
    .B1(net42),
    .Y(_02513_));
 sky130_fd_sc_hd__o22a_1 _21351_ (.A1(net742),
    .A2(net42),
    .B1(_02512_),
    .B2(_02513_),
    .X(_00337_));
 sky130_fd_sc_hd__nand2_1 _21352_ (.A(net595),
    .B(_04588_),
    .Y(_02514_));
 sky130_fd_sc_hd__o211a_1 _21353_ (.A1(net595),
    .A2(_09434_),
    .B1(net41),
    .C1(_02514_),
    .X(_02515_));
 sky130_fd_sc_hd__a21o_1 _21354_ (.A1(net801),
    .A2(net40),
    .B1(_02515_),
    .X(_00338_));
 sky130_fd_sc_hd__nand2_1 _21355_ (.A(net596),
    .B(_04719_),
    .Y(_02516_));
 sky130_fd_sc_hd__o211a_1 _21356_ (.A1(net596),
    .A2(_09564_),
    .B1(net42),
    .C1(_02516_),
    .X(_02517_));
 sky130_fd_sc_hd__a21o_1 _21357_ (.A1(net709),
    .A2(net39),
    .B1(_02517_),
    .X(_00339_));
 sky130_fd_sc_hd__nand2_1 _21358_ (.A(net60),
    .B(_09707_),
    .Y(_02518_));
 sky130_fd_sc_hd__a21oi_1 _21359_ (.A1(net595),
    .A2(_04862_),
    .B1(net40),
    .Y(_02519_));
 sky130_fd_sc_hd__a22o_1 _21360_ (.A1(net836),
    .A2(net40),
    .B1(_02518_),
    .B2(_02519_),
    .X(_00340_));
 sky130_fd_sc_hd__nand2_1 _21361_ (.A(net595),
    .B(_05006_),
    .Y(_02520_));
 sky130_fd_sc_hd__o211a_1 _21362_ (.A1(net595),
    .A2(_09851_),
    .B1(net41),
    .C1(_02520_),
    .X(_02521_));
 sky130_fd_sc_hd__a21o_1 _21363_ (.A1(net782),
    .A2(net40),
    .B1(_02521_),
    .X(_00341_));
 sky130_fd_sc_hd__nand2_1 _21364_ (.A(net595),
    .B(_05156_),
    .Y(_02522_));
 sky130_fd_sc_hd__o211a_1 _21365_ (.A1(net595),
    .A2(_09997_),
    .B1(net41),
    .C1(_02522_),
    .X(_02523_));
 sky130_fd_sc_hd__a21o_1 _21366_ (.A1(net740),
    .A2(net40),
    .B1(_02523_),
    .X(_00342_));
 sky130_fd_sc_hd__or2_1 _21367_ (.A(net596),
    .B(_10147_),
    .X(_02524_));
 sky130_fd_sc_hd__a21oi_1 _21368_ (.A1(net595),
    .A2(_05305_),
    .B1(net40),
    .Y(_02525_));
 sky130_fd_sc_hd__a22o_1 _21369_ (.A1(net796),
    .A2(net40),
    .B1(_02524_),
    .B2(_02525_),
    .X(_00343_));
 sky130_fd_sc_hd__o21ai_1 _21370_ (.A1(net60),
    .A2(_05457_),
    .B1(net41),
    .Y(_02526_));
 sky130_fd_sc_hd__a21oi_1 _21371_ (.A1(net60),
    .A2(_10299_),
    .B1(_02526_),
    .Y(_02527_));
 sky130_fd_sc_hd__a21o_1 _21372_ (.A1(net693),
    .A2(net40),
    .B1(_02527_),
    .X(_00344_));
 sky130_fd_sc_hd__nand2_1 _21373_ (.A(net60),
    .B(_10458_),
    .Y(_02528_));
 sky130_fd_sc_hd__o21a_1 _21374_ (.A1(net60),
    .A2(_05615_),
    .B1(net42),
    .X(_02529_));
 sky130_fd_sc_hd__a22o_1 _21375_ (.A1(net837),
    .A2(net39),
    .B1(_02528_),
    .B2(_02529_),
    .X(_00345_));
 sky130_fd_sc_hd__mux2_1 _21376_ (.A0(_05784_),
    .A1(_10625_),
    .S(net60),
    .X(_02530_));
 sky130_fd_sc_hd__mux2_1 _21377_ (.A0(net764),
    .A1(_02530_),
    .S(net42),
    .X(_00346_));
 sky130_fd_sc_hd__nand2_1 _21378_ (.A(net703),
    .B(net39),
    .Y(_02531_));
 sky130_fd_sc_hd__mux2_1 _21379_ (.A0(_05935_),
    .A1(_10777_),
    .S(net60),
    .X(_02532_));
 sky130_fd_sc_hd__o21ai_1 _21380_ (.A1(net39),
    .A2(_02532_),
    .B1(_02531_),
    .Y(_00347_));
 sky130_fd_sc_hd__nand2_1 _21381_ (.A(net757),
    .B(net39),
    .Y(_02533_));
 sky130_fd_sc_hd__mux2_1 _21382_ (.A0(_06090_),
    .A1(_00660_),
    .S(net60),
    .X(_02534_));
 sky130_fd_sc_hd__o21ai_1 _21383_ (.A1(net39),
    .A2(_02534_),
    .B1(_02533_),
    .Y(_00348_));
 sky130_fd_sc_hd__or2_1 _21384_ (.A(net596),
    .B(_00818_),
    .X(_02535_));
 sky130_fd_sc_hd__a21oi_1 _21385_ (.A1(net596),
    .A2(_06244_),
    .B1(net40),
    .Y(_02536_));
 sky130_fd_sc_hd__a22o_1 _21386_ (.A1(net815),
    .A2(net39),
    .B1(_02535_),
    .B2(_02536_),
    .X(_00349_));
 sky130_fd_sc_hd__nand2_1 _21387_ (.A(net60),
    .B(_00974_),
    .Y(_02537_));
 sky130_fd_sc_hd__o21a_1 _21388_ (.A1(net60),
    .A2(_06402_),
    .B1(net42),
    .X(_02538_));
 sky130_fd_sc_hd__a22o_1 _21389_ (.A1(net820),
    .A2(_02499_),
    .B1(_02537_),
    .B2(_02538_),
    .X(_00350_));
 sky130_fd_sc_hd__nand2_1 _21390_ (.A(net733),
    .B(_02499_),
    .Y(_02539_));
 sky130_fd_sc_hd__mux2_1 _21391_ (.A0(_06552_),
    .A1(_01125_),
    .S(net60),
    .X(_02540_));
 sky130_fd_sc_hd__o21ai_1 _21392_ (.A1(_02499_),
    .A2(_02540_),
    .B1(_02539_),
    .Y(_00351_));
 sky130_fd_sc_hd__nand2_1 _21393_ (.A(net60),
    .B(_01263_),
    .Y(_02541_));
 sky130_fd_sc_hd__a21oi_1 _21394_ (.A1(net596),
    .A2(_06691_),
    .B1(net39),
    .Y(_02542_));
 sky130_fd_sc_hd__a22o_1 _21395_ (.A1(net684),
    .A2(net40),
    .B1(_02541_),
    .B2(_02542_),
    .X(_00352_));
 sky130_fd_sc_hd__nor2_1 _21396_ (.A(net596),
    .B(_01407_),
    .Y(_02543_));
 sky130_fd_sc_hd__a21o_1 _21397_ (.A1(net596),
    .A2(_06837_),
    .B1(_02543_),
    .X(_02544_));
 sky130_fd_sc_hd__mux2_1 _21398_ (.A0(net813),
    .A1(_02544_),
    .S(net42),
    .X(_00353_));
 sky130_fd_sc_hd__nor2_1 _21399_ (.A(net60),
    .B(_06977_),
    .Y(_02545_));
 sky130_fd_sc_hd__a211o_1 _21400_ (.A1(net60),
    .A2(_01554_),
    .B1(net39),
    .C1(_02545_),
    .X(_02546_));
 sky130_fd_sc_hd__a21bo_1 _21401_ (.A1(net741),
    .A2(net40),
    .B1_N(_02546_),
    .X(_00354_));
 sky130_fd_sc_hd__mux2_1 _21402_ (.A0(_07105_),
    .A1(_01691_),
    .S(net61),
    .X(_02547_));
 sky130_fd_sc_hd__mux2_1 _21403_ (.A0(net831),
    .A1(_02547_),
    .S(net42),
    .X(_00355_));
 sky130_fd_sc_hd__nand2_1 _21404_ (.A(net595),
    .B(_07236_),
    .Y(_02548_));
 sky130_fd_sc_hd__o211a_1 _21405_ (.A1(net596),
    .A2(_01821_),
    .B1(net41),
    .C1(_02548_),
    .X(_02549_));
 sky130_fd_sc_hd__a21o_1 _21406_ (.A1(net758),
    .A2(net39),
    .B1(_02549_),
    .X(_00356_));
 sky130_fd_sc_hd__mux2_1 _21407_ (.A0(_07365_),
    .A1(_01944_),
    .S(net61),
    .X(_02550_));
 sky130_fd_sc_hd__mux2_1 _21408_ (.A0(net770),
    .A1(_02550_),
    .S(net41),
    .X(_00357_));
 sky130_fd_sc_hd__nand2_1 _21409_ (.A(net595),
    .B(_07499_),
    .Y(_02551_));
 sky130_fd_sc_hd__o211a_1 _21410_ (.A1(net595),
    .A2(_02080_),
    .B1(net41),
    .C1(_02551_),
    .X(_02552_));
 sky130_fd_sc_hd__a21o_1 _21411_ (.A1(net763),
    .A2(net40),
    .B1(_02552_),
    .X(_00358_));
 sky130_fd_sc_hd__nand2_1 _21412_ (.A(net595),
    .B(_07619_),
    .Y(_02553_));
 sky130_fd_sc_hd__o211a_1 _21413_ (.A1(net596),
    .A2(_02200_),
    .B1(net41),
    .C1(_02553_),
    .X(_02554_));
 sky130_fd_sc_hd__a21o_1 _21414_ (.A1(net723),
    .A2(net40),
    .B1(_02554_),
    .X(_00359_));
 sky130_fd_sc_hd__or2_1 _21415_ (.A(net596),
    .B(_02313_),
    .X(_02555_));
 sky130_fd_sc_hd__a21oi_1 _21416_ (.A1(net595),
    .A2(_07730_),
    .B1(net40),
    .Y(_02556_));
 sky130_fd_sc_hd__a22o_1 _21417_ (.A1(net835),
    .A2(net40),
    .B1(_02555_),
    .B2(_02556_),
    .X(_00360_));
 sky130_fd_sc_hd__mux2_1 _21418_ (.A0(_07835_),
    .A1(_02419_),
    .S(net60),
    .X(_02557_));
 sky130_fd_sc_hd__mux2_1 _21419_ (.A0(net841),
    .A1(_02557_),
    .S(net41),
    .X(_00361_));
 sky130_fd_sc_hd__mux2_1 _21420_ (.A0(_07909_),
    .A1(_02494_),
    .S(net60),
    .X(_02558_));
 sky130_fd_sc_hd__mux2_1 _21421_ (.A0(net833),
    .A1(_02558_),
    .S(net41),
    .X(_00362_));
 sky130_fd_sc_hd__and3_1 _21422_ (.A(net646),
    .B(sstream_o),
    .C(sstream_i[114]),
    .X(_02559_));
 sky130_fd_sc_hd__mux2_1 _21423_ (.A0(net871),
    .A1(sstream_i[0]),
    .S(net30),
    .X(_00363_));
 sky130_fd_sc_hd__mux2_1 _21424_ (.A0(net870),
    .A1(sstream_i[1]),
    .S(net30),
    .X(_00364_));
 sky130_fd_sc_hd__mux2_1 _21425_ (.A0(net868),
    .A1(sstream_i[2]),
    .S(net30),
    .X(_00365_));
 sky130_fd_sc_hd__mux2_1 _21426_ (.A0(net876),
    .A1(sstream_i[3]),
    .S(net31),
    .X(_00366_));
 sky130_fd_sc_hd__mux2_1 _21427_ (.A0(net895),
    .A1(sstream_i[4]),
    .S(net30),
    .X(_00367_));
 sky130_fd_sc_hd__mux2_1 _21428_ (.A0(net901),
    .A1(sstream_i[5]),
    .S(net30),
    .X(_00368_));
 sky130_fd_sc_hd__mux2_1 _21429_ (.A0(net877),
    .A1(sstream_i[6]),
    .S(net31),
    .X(_00369_));
 sky130_fd_sc_hd__mux2_1 _21430_ (.A0(net906),
    .A1(sstream_i[7]),
    .S(net31),
    .X(_00370_));
 sky130_fd_sc_hd__mux2_1 _21431_ (.A0(net894),
    .A1(sstream_i[8]),
    .S(net30),
    .X(_00371_));
 sky130_fd_sc_hd__mux2_1 _21432_ (.A0(net888),
    .A1(sstream_i[9]),
    .S(net30),
    .X(_00372_));
 sky130_fd_sc_hd__mux2_1 _21433_ (.A0(net924),
    .A1(sstream_i[10]),
    .S(net30),
    .X(_00373_));
 sky130_fd_sc_hd__mux2_1 _21434_ (.A0(net890),
    .A1(sstream_i[11]),
    .S(net30),
    .X(_00374_));
 sky130_fd_sc_hd__mux2_1 _21435_ (.A0(net896),
    .A1(sstream_i[12]),
    .S(net30),
    .X(_00375_));
 sky130_fd_sc_hd__mux2_1 _21436_ (.A0(net900),
    .A1(sstream_i[13]),
    .S(net30),
    .X(_00376_));
 sky130_fd_sc_hd__mux2_1 _21437_ (.A0(net912),
    .A1(sstream_i[14]),
    .S(net30),
    .X(_00377_));
 sky130_fd_sc_hd__mux2_1 _21438_ (.A0(net911),
    .A1(sstream_i[15]),
    .S(net30),
    .X(_00378_));
 sky130_fd_sc_hd__mux2_1 _21439_ (.A0(net928),
    .A1(sstream_i[16]),
    .S(net30),
    .X(_00379_));
 sky130_fd_sc_hd__mux2_1 _21440_ (.A0(net925),
    .A1(sstream_i[17]),
    .S(net31),
    .X(_00380_));
 sky130_fd_sc_hd__mux2_1 _21441_ (.A0(net941),
    .A1(sstream_i[18]),
    .S(net30),
    .X(_00381_));
 sky130_fd_sc_hd__mux2_1 _21442_ (.A0(net947),
    .A1(sstream_i[19]),
    .S(net30),
    .X(_00382_));
 sky130_fd_sc_hd__mux2_1 _21443_ (.A0(net913),
    .A1(sstream_i[20]),
    .S(net38),
    .X(_00383_));
 sky130_fd_sc_hd__mux2_1 _21444_ (.A0(net948),
    .A1(sstream_i[21]),
    .S(net31),
    .X(_00384_));
 sky130_fd_sc_hd__mux2_1 _21445_ (.A0(net943),
    .A1(sstream_i[22]),
    .S(net31),
    .X(_00385_));
 sky130_fd_sc_hd__mux2_1 _21446_ (.A0(net937),
    .A1(sstream_i[23]),
    .S(net31),
    .X(_00386_));
 sky130_fd_sc_hd__mux2_1 _21447_ (.A0(net942),
    .A1(sstream_i[24]),
    .S(net31),
    .X(_00387_));
 sky130_fd_sc_hd__mux2_1 _21448_ (.A0(net939),
    .A1(sstream_i[25]),
    .S(net31),
    .X(_00388_));
 sky130_fd_sc_hd__mux2_1 _21449_ (.A0(net765),
    .A1(sstream_i[26]),
    .S(net33),
    .X(_00389_));
 sky130_fd_sc_hd__mux2_1 _21450_ (.A0(net866),
    .A1(sstream_i[27]),
    .S(net32),
    .X(_00390_));
 sky130_fd_sc_hd__mux2_1 _21451_ (.A0(net860),
    .A1(sstream_i[28]),
    .S(net33),
    .X(_00391_));
 sky130_fd_sc_hd__mux2_1 _21452_ (.A0(net821),
    .A1(sstream_i[29]),
    .S(net34),
    .X(_00392_));
 sky130_fd_sc_hd__mux2_1 _21453_ (.A0(net766),
    .A1(sstream_i[30]),
    .S(net34),
    .X(_00393_));
 sky130_fd_sc_hd__mux2_1 _21454_ (.A0(net794),
    .A1(sstream_i[31]),
    .S(net34),
    .X(_00394_));
 sky130_fd_sc_hd__mux2_1 _21455_ (.A0(net806),
    .A1(sstream_i[32]),
    .S(net31),
    .X(_00395_));
 sky130_fd_sc_hd__mux2_1 _21456_ (.A0(net859),
    .A1(sstream_i[33]),
    .S(net31),
    .X(_00396_));
 sky130_fd_sc_hd__mux2_1 _21457_ (.A0(net855),
    .A1(sstream_i[34]),
    .S(net31),
    .X(_00397_));
 sky130_fd_sc_hd__mux2_1 _21458_ (.A0(net842),
    .A1(sstream_i[35]),
    .S(net32),
    .X(_00398_));
 sky130_fd_sc_hd__mux2_1 _21459_ (.A0(net823),
    .A1(sstream_i[36]),
    .S(net32),
    .X(_00399_));
 sky130_fd_sc_hd__mux2_1 _21460_ (.A0(net785),
    .A1(sstream_i[37]),
    .S(net32),
    .X(_00400_));
 sky130_fd_sc_hd__mux2_1 _21461_ (.A0(net850),
    .A1(sstream_i[38]),
    .S(net33),
    .X(_00401_));
 sky130_fd_sc_hd__mux2_1 _21462_ (.A0(net828),
    .A1(sstream_i[39]),
    .S(net32),
    .X(_00402_));
 sky130_fd_sc_hd__mux2_1 _21463_ (.A0(net829),
    .A1(sstream_i[40]),
    .S(net32),
    .X(_00403_));
 sky130_fd_sc_hd__mux2_1 _21464_ (.A0(net845),
    .A1(sstream_i[41]),
    .S(net32),
    .X(_00404_));
 sky130_fd_sc_hd__mux2_1 _21465_ (.A0(net856),
    .A1(sstream_i[42]),
    .S(net32),
    .X(_00405_));
 sky130_fd_sc_hd__mux2_1 _21466_ (.A0(net857),
    .A1(sstream_i[43]),
    .S(net32),
    .X(_00406_));
 sky130_fd_sc_hd__mux2_1 _21467_ (.A0(net769),
    .A1(sstream_i[44]),
    .S(net32),
    .X(_00407_));
 sky130_fd_sc_hd__mux2_1 _21468_ (.A0(net816),
    .A1(sstream_i[45]),
    .S(net33),
    .X(_00408_));
 sky130_fd_sc_hd__mux2_1 _21469_ (.A0(net844),
    .A1(sstream_i[46]),
    .S(net33),
    .X(_00409_));
 sky130_fd_sc_hd__mux2_1 _21470_ (.A0(net799),
    .A1(sstream_i[47]),
    .S(net32),
    .X(_00410_));
 sky130_fd_sc_hd__mux2_1 _21471_ (.A0(net800),
    .A1(sstream_i[48]),
    .S(net32),
    .X(_00411_));
 sky130_fd_sc_hd__mux2_1 _21472_ (.A0(net830),
    .A1(sstream_i[49]),
    .S(net33),
    .X(_00412_));
 sky130_fd_sc_hd__mux2_1 _21473_ (.A0(net808),
    .A1(sstream_i[50]),
    .S(net33),
    .X(_00413_));
 sky130_fd_sc_hd__mux2_1 _21474_ (.A0(net788),
    .A1(sstream_i[51]),
    .S(net33),
    .X(_00414_));
 sky130_fd_sc_hd__mux2_1 _21475_ (.A0(net812),
    .A1(sstream_i[52]),
    .S(net33),
    .X(_00415_));
 sky130_fd_sc_hd__mux2_1 _21476_ (.A0(net777),
    .A1(sstream_i[53]),
    .S(net33),
    .X(_00416_));
 sky130_fd_sc_hd__mux2_1 _21477_ (.A0(net762),
    .A1(sstream_i[54]),
    .S(net33),
    .X(_00417_));
 sky130_fd_sc_hd__mux2_1 _21478_ (.A0(net810),
    .A1(sstream_i[55]),
    .S(net33),
    .X(_00418_));
 sky130_fd_sc_hd__mux2_1 _21479_ (.A0(net776),
    .A1(sstream_i[56]),
    .S(net33),
    .X(_00419_));
 sky130_fd_sc_hd__mux2_1 _21480_ (.A0(net853),
    .A1(sstream_i[57]),
    .S(net33),
    .X(_00420_));
 sky130_fd_sc_hd__mux2_1 _21481_ (.A0(net824),
    .A1(sstream_i[58]),
    .S(net33),
    .X(_00421_));
 sky130_fd_sc_hd__mux2_1 _21482_ (.A0(net807),
    .A1(sstream_i[59]),
    .S(net34),
    .X(_00422_));
 sky130_fd_sc_hd__mux2_1 _21483_ (.A0(net827),
    .A1(sstream_i[60]),
    .S(net34),
    .X(_00423_));
 sky130_fd_sc_hd__mux2_1 _21484_ (.A0(net826),
    .A1(sstream_i[61]),
    .S(net34),
    .X(_00424_));
 sky130_fd_sc_hd__mux2_1 _21485_ (.A0(net847),
    .A1(sstream_i[62]),
    .S(net34),
    .X(_00425_));
 sky130_fd_sc_hd__mux2_1 _21486_ (.A0(net848),
    .A1(sstream_i[63]),
    .S(net34),
    .X(_00426_));
 sky130_fd_sc_hd__mux2_1 _21487_ (.A0(net846),
    .A1(sstream_i[64]),
    .S(net31),
    .X(_00427_));
 sky130_fd_sc_hd__mux2_1 _21488_ (.A0(net843),
    .A1(sstream_i[65]),
    .S(net31),
    .X(_00428_));
 sky130_fd_sc_hd__mux2_1 _21489_ (.A0(net822),
    .A1(sstream_i[66]),
    .S(net31),
    .X(_00429_));
 sky130_fd_sc_hd__mux2_1 _21490_ (.A0(net838),
    .A1(sstream_i[67]),
    .S(net38),
    .X(_00430_));
 sky130_fd_sc_hd__mux2_1 _21491_ (.A0(net811),
    .A1(sstream_i[68]),
    .S(net32),
    .X(_00431_));
 sky130_fd_sc_hd__mux2_1 _21492_ (.A0(net832),
    .A1(sstream_i[69]),
    .S(net32),
    .X(_00432_));
 sky130_fd_sc_hd__mux2_1 _21493_ (.A0(net825),
    .A1(sstream_i[70]),
    .S(net32),
    .X(_00433_));
 sky130_fd_sc_hd__mux2_1 _21494_ (.A0(net795),
    .A1(sstream_i[71]),
    .S(net32),
    .X(_00434_));
 sky130_fd_sc_hd__mux2_1 _21495_ (.A0(net944),
    .A1(sstream_i[72]),
    .S(net34),
    .X(_00435_));
 sky130_fd_sc_hd__mux2_1 _21496_ (.A0(net954),
    .A1(sstream_i[73]),
    .S(net35),
    .X(_00436_));
 sky130_fd_sc_hd__mux2_1 _21497_ (.A0(net962),
    .A1(sstream_i[74]),
    .S(net34),
    .X(_00437_));
 sky130_fd_sc_hd__mux2_1 _21498_ (.A0(net907),
    .A1(sstream_i[75]),
    .S(net35),
    .X(_00438_));
 sky130_fd_sc_hd__mux2_1 _21499_ (.A0(net949),
    .A1(sstream_i[76]),
    .S(net35),
    .X(_00439_));
 sky130_fd_sc_hd__mux2_1 _21500_ (.A0(net938),
    .A1(sstream_i[77]),
    .S(net35),
    .X(_00440_));
 sky130_fd_sc_hd__mux2_1 _21501_ (.A0(net950),
    .A1(sstream_i[78]),
    .S(net35),
    .X(_00441_));
 sky130_fd_sc_hd__mux2_1 _21502_ (.A0(net915),
    .A1(sstream_i[79]),
    .S(net34),
    .X(_00442_));
 sky130_fd_sc_hd__mux2_1 _21503_ (.A0(net931),
    .A1(sstream_i[80]),
    .S(net34),
    .X(_00443_));
 sky130_fd_sc_hd__mux2_1 _21504_ (.A0(net957),
    .A1(sstream_i[81]),
    .S(net34),
    .X(_00444_));
 sky130_fd_sc_hd__mux2_1 _21505_ (.A0(net927),
    .A1(sstream_i[82]),
    .S(net34),
    .X(_00445_));
 sky130_fd_sc_hd__mux2_1 _21506_ (.A0(net892),
    .A1(sstream_i[83]),
    .S(net34),
    .X(_00446_));
 sky130_fd_sc_hd__mux2_1 _21507_ (.A0(net881),
    .A1(sstream_i[84]),
    .S(net34),
    .X(_00447_));
 sky130_fd_sc_hd__mux2_1 _21508_ (.A0(net926),
    .A1(sstream_i[85]),
    .S(net35),
    .X(_00448_));
 sky130_fd_sc_hd__mux2_1 _21509_ (.A0(net951),
    .A1(sstream_i[86]),
    .S(net35),
    .X(_00449_));
 sky130_fd_sc_hd__mux2_1 _21510_ (.A0(net879),
    .A1(sstream_i[87]),
    .S(net35),
    .X(_00450_));
 sky130_fd_sc_hd__mux2_1 _21511_ (.A0(net917),
    .A1(sstream_i[88]),
    .S(net36),
    .X(_00451_));
 sky130_fd_sc_hd__mux2_1 _21512_ (.A0(net874),
    .A1(sstream_i[89]),
    .S(net36),
    .X(_00452_));
 sky130_fd_sc_hd__mux2_1 _21513_ (.A0(net918),
    .A1(sstream_i[90]),
    .S(net36),
    .X(_00453_));
 sky130_fd_sc_hd__mux2_1 _21514_ (.A0(net884),
    .A1(sstream_i[91]),
    .S(net36),
    .X(_00454_));
 sky130_fd_sc_hd__mux2_1 _21515_ (.A0(net891),
    .A1(sstream_i[92]),
    .S(net36),
    .X(_00455_));
 sky130_fd_sc_hd__mux2_1 _21516_ (.A0(net882),
    .A1(sstream_i[93]),
    .S(net36),
    .X(_00456_));
 sky130_fd_sc_hd__mux2_1 _21517_ (.A0(net883),
    .A1(sstream_i[94]),
    .S(net36),
    .X(_00457_));
 sky130_fd_sc_hd__mux2_1 _21518_ (.A0(net897),
    .A1(sstream_i[95]),
    .S(net36),
    .X(_00458_));
 sky130_fd_sc_hd__mux2_1 _21519_ (.A0(net880),
    .A1(sstream_i[96]),
    .S(net36),
    .X(_00459_));
 sky130_fd_sc_hd__mux2_1 _21520_ (.A0(net904),
    .A1(sstream_i[97]),
    .S(net36),
    .X(_00460_));
 sky130_fd_sc_hd__mux2_1 _21521_ (.A0(net885),
    .A1(sstream_i[98]),
    .S(net36),
    .X(_00461_));
 sky130_fd_sc_hd__mux2_1 _21522_ (.A0(net902),
    .A1(sstream_i[99]),
    .S(net36),
    .X(_00462_));
 sky130_fd_sc_hd__mux2_1 _21523_ (.A0(net936),
    .A1(sstream_i[100]),
    .S(net37),
    .X(_00463_));
 sky130_fd_sc_hd__mux2_1 _21524_ (.A0(net893),
    .A1(sstream_i[101]),
    .S(net37),
    .X(_00464_));
 sky130_fd_sc_hd__mux2_1 _21525_ (.A0(net921),
    .A1(sstream_i[102]),
    .S(net36),
    .X(_00465_));
 sky130_fd_sc_hd__mux2_1 _21526_ (.A0(net955),
    .A1(sstream_i[103]),
    .S(net36),
    .X(_00466_));
 sky130_fd_sc_hd__mux2_1 _21527_ (.A0(net932),
    .A1(sstream_i[104]),
    .S(net36),
    .X(_00467_));
 sky130_fd_sc_hd__mux2_1 _21528_ (.A0(net916),
    .A1(sstream_i[105]),
    .S(net36),
    .X(_00468_));
 sky130_fd_sc_hd__mux2_1 _21529_ (.A0(net945),
    .A1(sstream_i[106]),
    .S(net37),
    .X(_00469_));
 sky130_fd_sc_hd__mux2_1 _21530_ (.A0(net934),
    .A1(sstream_i[107]),
    .S(net37),
    .X(_00470_));
 sky130_fd_sc_hd__mux2_1 _21531_ (.A0(net920),
    .A1(sstream_i[108]),
    .S(net37),
    .X(_00471_));
 sky130_fd_sc_hd__mux2_1 _21532_ (.A0(net908),
    .A1(sstream_i[109]),
    .S(net37),
    .X(_00472_));
 sky130_fd_sc_hd__mux2_1 _21533_ (.A0(net952),
    .A1(sstream_i[110]),
    .S(net37),
    .X(_00473_));
 sky130_fd_sc_hd__mux2_1 _21534_ (.A0(net914),
    .A1(sstream_i[111]),
    .S(net37),
    .X(_00474_));
 sky130_fd_sc_hd__mux2_1 _21535_ (.A0(net923),
    .A1(sstream_i[112]),
    .S(net37),
    .X(_00475_));
 sky130_fd_sc_hd__mux2_1 _21536_ (.A0(net929),
    .A1(sstream_i[113]),
    .S(net37),
    .X(_00476_));
 sky130_fd_sc_hd__mux2_1 _21537_ (.A0(mstream_o[0]),
    .A1(net659),
    .S(net612),
    .X(_00477_));
 sky130_fd_sc_hd__mux2_1 _21538_ (.A0(mstream_o[1]),
    .A1(net655),
    .S(net612),
    .X(_00478_));
 sky130_fd_sc_hd__mux2_1 _21539_ (.A0(mstream_o[2]),
    .A1(net731),
    .S(net612),
    .X(_00479_));
 sky130_fd_sc_hd__mux2_1 _21540_ (.A0(mstream_o[3]),
    .A1(net667),
    .S(net612),
    .X(_00480_));
 sky130_fd_sc_hd__mux2_1 _21541_ (.A0(mstream_o[4]),
    .A1(net650),
    .S(net612),
    .X(_00481_));
 sky130_fd_sc_hd__mux2_1 _21542_ (.A0(mstream_o[5]),
    .A1(net661),
    .S(net612),
    .X(_00482_));
 sky130_fd_sc_hd__mux2_1 _21543_ (.A0(mstream_o[6]),
    .A1(net662),
    .S(net612),
    .X(_00483_));
 sky130_fd_sc_hd__mux2_1 _21544_ (.A0(mstream_o[7]),
    .A1(net665),
    .S(net612),
    .X(_00484_));
 sky130_fd_sc_hd__mux2_1 _21545_ (.A0(mstream_o[8]),
    .A1(net679),
    .S(net612),
    .X(_00485_));
 sky130_fd_sc_hd__mux2_1 _21546_ (.A0(mstream_o[9]),
    .A1(net819),
    .S(net612),
    .X(_00486_));
 sky130_fd_sc_hd__mux2_1 _21547_ (.A0(mstream_o[10]),
    .A1(net728),
    .S(net612),
    .X(_00487_));
 sky130_fd_sc_hd__mux2_1 _21548_ (.A0(mstream_o[11]),
    .A1(net695),
    .S(net612),
    .X(_00488_));
 sky130_fd_sc_hd__mux2_1 _21549_ (.A0(mstream_o[12]),
    .A1(net798),
    .S(net612),
    .X(_00489_));
 sky130_fd_sc_hd__mux2_1 _21550_ (.A0(mstream_o[13]),
    .A1(net677),
    .S(net613),
    .X(_00490_));
 sky130_fd_sc_hd__mux2_1 _21551_ (.A0(mstream_o[14]),
    .A1(net654),
    .S(net613),
    .X(_00491_));
 sky130_fd_sc_hd__mux2_1 _21552_ (.A0(mstream_o[15]),
    .A1(net752),
    .S(net612),
    .X(_00492_));
 sky130_fd_sc_hd__mux2_1 _21553_ (.A0(mstream_o[16]),
    .A1(net719),
    .S(net612),
    .X(_00493_));
 sky130_fd_sc_hd__mux2_1 _21554_ (.A0(mstream_o[17]),
    .A1(net678),
    .S(net612),
    .X(_00494_));
 sky130_fd_sc_hd__mux2_1 _21555_ (.A0(mstream_o[18]),
    .A1(net663),
    .S(net613),
    .X(_00495_));
 sky130_fd_sc_hd__mux2_1 _21556_ (.A0(mstream_o[19]),
    .A1(net790),
    .S(net613),
    .X(_00496_));
 sky130_fd_sc_hd__mux2_1 _21557_ (.A0(mstream_o[20]),
    .A1(net710),
    .S(net613),
    .X(_00497_));
 sky130_fd_sc_hd__mux2_1 _21558_ (.A0(mstream_o[21]),
    .A1(net672),
    .S(net613),
    .X(_00498_));
 sky130_fd_sc_hd__mux2_1 _21559_ (.A0(mstream_o[22]),
    .A1(net814),
    .S(net613),
    .X(_00499_));
 sky130_fd_sc_hd__mux2_1 _21560_ (.A0(mstream_o[23]),
    .A1(net700),
    .S(net613),
    .X(_00500_));
 sky130_fd_sc_hd__mux2_1 _21561_ (.A0(mstream_o[24]),
    .A1(net689),
    .S(net613),
    .X(_00501_));
 sky130_fd_sc_hd__mux2_1 _21562_ (.A0(mstream_o[25]),
    .A1(net674),
    .S(net613),
    .X(_00502_));
 sky130_fd_sc_hd__mux2_1 _21563_ (.A0(mstream_o[26]),
    .A1(net658),
    .S(net614),
    .X(_00503_));
 sky130_fd_sc_hd__mux2_1 _21564_ (.A0(mstream_o[27]),
    .A1(net691),
    .S(net614),
    .X(_00504_));
 sky130_fd_sc_hd__mux2_1 _21565_ (.A0(mstream_o[28]),
    .A1(net651),
    .S(net614),
    .X(_00505_));
 sky130_fd_sc_hd__mux2_1 _21566_ (.A0(mstream_o[29]),
    .A1(net707),
    .S(net614),
    .X(_00506_));
 sky130_fd_sc_hd__mux2_1 _21567_ (.A0(mstream_o[30]),
    .A1(net699),
    .S(net616),
    .X(_00507_));
 sky130_fd_sc_hd__mux2_1 _21568_ (.A0(mstream_o[31]),
    .A1(net713),
    .S(net616),
    .X(_00508_));
 sky130_fd_sc_hd__mux2_1 _21569_ (.A0(mstream_o[32]),
    .A1(_02738_),
    .S(net614),
    .X(_00509_));
 sky130_fd_sc_hd__mux2_1 _21570_ (.A0(mstream_o[33]),
    .A1(_02739_),
    .S(net614),
    .X(_00510_));
 sky130_fd_sc_hd__mux2_1 _21571_ (.A0(mstream_o[34]),
    .A1(_02741_),
    .S(net614),
    .X(_00511_));
 sky130_fd_sc_hd__mux2_1 _21572_ (.A0(mstream_o[35]),
    .A1(_02743_),
    .S(net614),
    .X(_00512_));
 sky130_fd_sc_hd__mux2_1 _21573_ (.A0(mstream_o[36]),
    .A1(_02744_),
    .S(net614),
    .X(_00513_));
 sky130_fd_sc_hd__mux2_1 _21574_ (.A0(mstream_o[37]),
    .A1(_02745_),
    .S(net614),
    .X(_00514_));
 sky130_fd_sc_hd__mux2_1 _21575_ (.A0(mstream_o[38]),
    .A1(_02746_),
    .S(net614),
    .X(_00515_));
 sky130_fd_sc_hd__mux2_1 _21576_ (.A0(mstream_o[39]),
    .A1(_02747_),
    .S(net614),
    .X(_00516_));
 sky130_fd_sc_hd__mux2_1 _21577_ (.A0(mstream_o[40]),
    .A1(_02748_),
    .S(net614),
    .X(_00517_));
 sky130_fd_sc_hd__mux2_1 _21578_ (.A0(mstream_o[41]),
    .A1(_02749_),
    .S(net614),
    .X(_00518_));
 sky130_fd_sc_hd__mux2_1 _21579_ (.A0(mstream_o[42]),
    .A1(_02751_),
    .S(net614),
    .X(_00519_));
 sky130_fd_sc_hd__dfrtp_4 _21580_ (.CLK(clknet_leaf_31_clk_i),
    .D(_00003_),
    .RESET_B(net637),
    .Q(mstream_o[43]));
 sky130_fd_sc_hd__dfrtp_4 _21581_ (.CLK(clknet_leaf_31_clk_i),
    .D(_00004_),
    .RESET_B(net638),
    .Q(mstream_o[44]));
 sky130_fd_sc_hd__dfrtp_4 _21582_ (.CLK(clknet_leaf_31_clk_i),
    .D(_00005_),
    .RESET_B(net637),
    .Q(mstream_o[45]));
 sky130_fd_sc_hd__dfrtp_4 _21583_ (.CLK(clknet_leaf_31_clk_i),
    .D(_00006_),
    .RESET_B(net637),
    .Q(mstream_o[46]));
 sky130_fd_sc_hd__dfrtp_4 _21584_ (.CLK(clknet_leaf_31_clk_i),
    .D(_00007_),
    .RESET_B(net637),
    .Q(mstream_o[47]));
 sky130_fd_sc_hd__dfrtp_4 _21585_ (.CLK(clknet_leaf_26_clk_i),
    .D(_00008_),
    .RESET_B(net640),
    .Q(mstream_o[48]));
 sky130_fd_sc_hd__dfrtp_4 _21586_ (.CLK(clknet_leaf_26_clk_i),
    .D(_00009_),
    .RESET_B(net640),
    .Q(mstream_o[49]));
 sky130_fd_sc_hd__dfrtp_4 _21587_ (.CLK(clknet_leaf_26_clk_i),
    .D(_00010_),
    .RESET_B(net640),
    .Q(mstream_o[50]));
 sky130_fd_sc_hd__dfrtp_4 _21588_ (.CLK(clknet_leaf_26_clk_i),
    .D(_00011_),
    .RESET_B(net640),
    .Q(mstream_o[51]));
 sky130_fd_sc_hd__dfrtp_4 _21589_ (.CLK(clknet_leaf_26_clk_i),
    .D(_00012_),
    .RESET_B(net640),
    .Q(mstream_o[52]));
 sky130_fd_sc_hd__dfrtp_4 _21590_ (.CLK(clknet_leaf_26_clk_i),
    .D(_00013_),
    .RESET_B(net640),
    .Q(mstream_o[53]));
 sky130_fd_sc_hd__dfrtp_4 _21591_ (.CLK(clknet_leaf_26_clk_i),
    .D(_00014_),
    .RESET_B(net640),
    .Q(mstream_o[54]));
 sky130_fd_sc_hd__dfrtp_4 _21592_ (.CLK(clknet_leaf_26_clk_i),
    .D(_00015_),
    .RESET_B(net640),
    .Q(mstream_o[55]));
 sky130_fd_sc_hd__dfrtp_4 _21593_ (.CLK(clknet_leaf_26_clk_i),
    .D(_00016_),
    .RESET_B(net642),
    .Q(mstream_o[56]));
 sky130_fd_sc_hd__dfrtp_4 _21594_ (.CLK(clknet_leaf_26_clk_i),
    .D(_00017_),
    .RESET_B(net642),
    .Q(mstream_o[57]));
 sky130_fd_sc_hd__dfrtp_4 _21595_ (.CLK(clknet_leaf_25_clk_i),
    .D(_00018_),
    .RESET_B(net640),
    .Q(mstream_o[58]));
 sky130_fd_sc_hd__dfrtp_4 _21596_ (.CLK(clknet_leaf_25_clk_i),
    .D(_00019_),
    .RESET_B(net640),
    .Q(mstream_o[59]));
 sky130_fd_sc_hd__dfrtp_4 _21597_ (.CLK(clknet_leaf_26_clk_i),
    .D(_00020_),
    .RESET_B(net640),
    .Q(mstream_o[60]));
 sky130_fd_sc_hd__dfrtp_4 _21598_ (.CLK(clknet_leaf_26_clk_i),
    .D(_00021_),
    .RESET_B(net640),
    .Q(mstream_o[61]));
 sky130_fd_sc_hd__dfrtp_4 _21599_ (.CLK(clknet_leaf_25_clk_i),
    .D(_00022_),
    .RESET_B(net640),
    .Q(mstream_o[62]));
 sky130_fd_sc_hd__dfrtp_4 _21600_ (.CLK(clknet_leaf_25_clk_i),
    .D(_00023_),
    .RESET_B(net641),
    .Q(mstream_o[63]));
 sky130_fd_sc_hd__dfrtp_4 _21601_ (.CLK(clknet_leaf_26_clk_i),
    .D(_00024_),
    .RESET_B(net640),
    .Q(mstream_o[64]));
 sky130_fd_sc_hd__dfrtp_4 _21602_ (.CLK(clknet_leaf_26_clk_i),
    .D(_00025_),
    .RESET_B(net642),
    .Q(mstream_o[65]));
 sky130_fd_sc_hd__dfrtp_4 _21603_ (.CLK(clknet_leaf_26_clk_i),
    .D(_00026_),
    .RESET_B(net640),
    .Q(mstream_o[66]));
 sky130_fd_sc_hd__dfrtp_4 _21604_ (.CLK(clknet_leaf_25_clk_i),
    .D(_00027_),
    .RESET_B(net640),
    .Q(mstream_o[67]));
 sky130_fd_sc_hd__dfrtp_4 _21605_ (.CLK(clknet_leaf_25_clk_i),
    .D(_00028_),
    .RESET_B(net641),
    .Q(mstream_o[68]));
 sky130_fd_sc_hd__dfrtp_4 _21606_ (.CLK(clknet_leaf_25_clk_i),
    .D(_00029_),
    .RESET_B(net642),
    .Q(mstream_o[69]));
 sky130_fd_sc_hd__dfrtp_4 _21607_ (.CLK(clknet_leaf_24_clk_i),
    .D(_00030_),
    .RESET_B(net641),
    .Q(mstream_o[70]));
 sky130_fd_sc_hd__dfrtp_4 _21608_ (.CLK(clknet_leaf_25_clk_i),
    .D(_00031_),
    .RESET_B(net641),
    .Q(mstream_o[71]));
 sky130_fd_sc_hd__dfrtp_4 _21609_ (.CLK(clknet_leaf_25_clk_i),
    .D(_00032_),
    .RESET_B(net641),
    .Q(mstream_o[72]));
 sky130_fd_sc_hd__dfrtp_4 _21610_ (.CLK(clknet_leaf_24_clk_i),
    .D(_00033_),
    .RESET_B(net641),
    .Q(mstream_o[73]));
 sky130_fd_sc_hd__dfrtp_4 _21611_ (.CLK(clknet_leaf_25_clk_i),
    .D(_00034_),
    .RESET_B(net641),
    .Q(mstream_o[74]));
 sky130_fd_sc_hd__dfrtp_4 _21612_ (.CLK(clknet_leaf_24_clk_i),
    .D(_00035_),
    .RESET_B(net641),
    .Q(mstream_o[75]));
 sky130_fd_sc_hd__dfrtp_4 _21613_ (.CLK(clknet_leaf_24_clk_i),
    .D(_00036_),
    .RESET_B(net641),
    .Q(mstream_o[76]));
 sky130_fd_sc_hd__dfrtp_4 _21614_ (.CLK(clknet_leaf_24_clk_i),
    .D(_00037_),
    .RESET_B(net641),
    .Q(mstream_o[77]));
 sky130_fd_sc_hd__dfrtp_4 _21615_ (.CLK(clknet_leaf_24_clk_i),
    .D(_00038_),
    .RESET_B(net641),
    .Q(mstream_o[78]));
 sky130_fd_sc_hd__dfrtp_4 _21616_ (.CLK(clknet_leaf_24_clk_i),
    .D(_00039_),
    .RESET_B(net641),
    .Q(mstream_o[79]));
 sky130_fd_sc_hd__dfrtp_4 _21617_ (.CLK(clknet_leaf_24_clk_i),
    .D(_00040_),
    .RESET_B(net641),
    .Q(mstream_o[80]));
 sky130_fd_sc_hd__dfrtp_4 _21618_ (.CLK(clknet_leaf_24_clk_i),
    .D(_00041_),
    .RESET_B(net641),
    .Q(mstream_o[81]));
 sky130_fd_sc_hd__dfrtp_4 _21619_ (.CLK(clknet_leaf_20_clk_i),
    .D(_00042_),
    .RESET_B(net644),
    .Q(mstream_o[82]));
 sky130_fd_sc_hd__dfrtp_4 _21620_ (.CLK(clknet_leaf_24_clk_i),
    .D(_00043_),
    .RESET_B(net641),
    .Q(mstream_o[83]));
 sky130_fd_sc_hd__dfrtp_4 _21621_ (.CLK(clknet_leaf_20_clk_i),
    .D(_00044_),
    .RESET_B(net644),
    .Q(mstream_o[84]));
 sky130_fd_sc_hd__dfrtp_4 _21622_ (.CLK(clknet_leaf_20_clk_i),
    .D(_00045_),
    .RESET_B(net644),
    .Q(mstream_o[85]));
 sky130_fd_sc_hd__dfrtp_4 _21623_ (.CLK(clknet_leaf_20_clk_i),
    .D(_00046_),
    .RESET_B(net644),
    .Q(mstream_o[86]));
 sky130_fd_sc_hd__dfrtp_4 _21624_ (.CLK(clknet_leaf_20_clk_i),
    .D(_00047_),
    .RESET_B(net644),
    .Q(mstream_o[87]));
 sky130_fd_sc_hd__dfrtp_4 _21625_ (.CLK(clknet_leaf_19_clk_i),
    .D(_00048_),
    .RESET_B(net644),
    .Q(mstream_o[88]));
 sky130_fd_sc_hd__dfrtp_4 _21626_ (.CLK(clknet_leaf_19_clk_i),
    .D(_00049_),
    .RESET_B(net644),
    .Q(mstream_o[89]));
 sky130_fd_sc_hd__dfrtp_4 _21627_ (.CLK(clknet_leaf_19_clk_i),
    .D(_00050_),
    .RESET_B(net644),
    .Q(mstream_o[90]));
 sky130_fd_sc_hd__dfrtp_4 _21628_ (.CLK(clknet_leaf_19_clk_i),
    .D(_00051_),
    .RESET_B(net644),
    .Q(mstream_o[91]));
 sky130_fd_sc_hd__dfrtp_4 _21629_ (.CLK(clknet_leaf_19_clk_i),
    .D(_00052_),
    .RESET_B(net644),
    .Q(mstream_o[92]));
 sky130_fd_sc_hd__dfrtp_4 _21630_ (.CLK(clknet_leaf_19_clk_i),
    .D(_00053_),
    .RESET_B(net644),
    .Q(mstream_o[93]));
 sky130_fd_sc_hd__dfrtp_4 _21631_ (.CLK(clknet_leaf_19_clk_i),
    .D(_00054_),
    .RESET_B(net644),
    .Q(mstream_o[94]));
 sky130_fd_sc_hd__dfrtp_4 _21632_ (.CLK(clknet_leaf_19_clk_i),
    .D(_00055_),
    .RESET_B(net644),
    .Q(mstream_o[95]));
 sky130_fd_sc_hd__dfrtp_4 _21633_ (.CLK(clknet_leaf_19_clk_i),
    .D(_00056_),
    .RESET_B(net644),
    .Q(mstream_o[96]));
 sky130_fd_sc_hd__dfrtp_4 _21634_ (.CLK(clknet_leaf_19_clk_i),
    .D(net905),
    .RESET_B(net644),
    .Q(mstream_o[97]));
 sky130_fd_sc_hd__dfrtp_4 _21635_ (.CLK(clknet_leaf_19_clk_i),
    .D(net886),
    .RESET_B(net643),
    .Q(mstream_o[98]));
 sky130_fd_sc_hd__dfrtp_4 _21636_ (.CLK(clknet_leaf_18_clk_i),
    .D(net903),
    .RESET_B(net643),
    .Q(mstream_o[99]));
 sky130_fd_sc_hd__dfrtp_4 _21637_ (.CLK(clknet_leaf_18_clk_i),
    .D(_00060_),
    .RESET_B(net643),
    .Q(mstream_o[100]));
 sky130_fd_sc_hd__dfrtp_4 _21638_ (.CLK(clknet_leaf_19_clk_i),
    .D(_00061_),
    .RESET_B(net643),
    .Q(mstream_o[101]));
 sky130_fd_sc_hd__dfrtp_4 _21639_ (.CLK(clknet_leaf_18_clk_i),
    .D(_00062_),
    .RESET_B(net643),
    .Q(mstream_o[102]));
 sky130_fd_sc_hd__dfrtp_4 _21640_ (.CLK(clknet_leaf_18_clk_i),
    .D(net956),
    .RESET_B(net643),
    .Q(mstream_o[103]));
 sky130_fd_sc_hd__dfrtp_4 _21641_ (.CLK(clknet_leaf_18_clk_i),
    .D(net933),
    .RESET_B(net643),
    .Q(mstream_o[104]));
 sky130_fd_sc_hd__dfrtp_4 _21642_ (.CLK(clknet_leaf_18_clk_i),
    .D(_00065_),
    .RESET_B(net643),
    .Q(mstream_o[105]));
 sky130_fd_sc_hd__dfrtp_4 _21643_ (.CLK(clknet_leaf_18_clk_i),
    .D(net946),
    .RESET_B(net643),
    .Q(mstream_o[106]));
 sky130_fd_sc_hd__dfrtp_4 _21644_ (.CLK(clknet_leaf_18_clk_i),
    .D(net935),
    .RESET_B(net643),
    .Q(mstream_o[107]));
 sky130_fd_sc_hd__dfrtp_4 _21645_ (.CLK(clknet_leaf_18_clk_i),
    .D(_00068_),
    .RESET_B(net643),
    .Q(mstream_o[108]));
 sky130_fd_sc_hd__dfrtp_4 _21646_ (.CLK(clknet_leaf_18_clk_i),
    .D(_00069_),
    .RESET_B(net643),
    .Q(mstream_o[109]));
 sky130_fd_sc_hd__dfrtp_4 _21647_ (.CLK(clknet_leaf_18_clk_i),
    .D(net953),
    .RESET_B(net643),
    .Q(mstream_o[110]));
 sky130_fd_sc_hd__dfrtp_4 _21648_ (.CLK(clknet_leaf_18_clk_i),
    .D(_00071_),
    .RESET_B(net643),
    .Q(mstream_o[111]));
 sky130_fd_sc_hd__dfrtp_4 _21649_ (.CLK(clknet_leaf_18_clk_i),
    .D(_00072_),
    .RESET_B(net643),
    .Q(mstream_o[112]));
 sky130_fd_sc_hd__dfrtp_4 _21650_ (.CLK(clknet_leaf_18_clk_i),
    .D(net930),
    .RESET_B(net643),
    .Q(mstream_o[113]));
 sky130_fd_sc_hd__dfrtp_4 _21651_ (.CLK(clknet_leaf_13_clk_i),
    .D(_00074_),
    .RESET_B(net646),
    .Q(mstream_o[115]));
 sky130_fd_sc_hd__dfxtp_1 _21652_ (.CLK(clknet_leaf_26_clk_i),
    .D(_00075_),
    .Q(\tx[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21653_ (.CLK(clknet_leaf_26_clk_i),
    .D(_00076_),
    .Q(\tx[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21654_ (.CLK(clknet_leaf_26_clk_i),
    .D(_00077_),
    .Q(\tx[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21655_ (.CLK(clknet_leaf_26_clk_i),
    .D(_00078_),
    .Q(\tx[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21656_ (.CLK(clknet_leaf_25_clk_i),
    .D(_00079_),
    .Q(\tx[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21657_ (.CLK(clknet_leaf_25_clk_i),
    .D(_00080_),
    .Q(\tx[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21658_ (.CLK(clknet_leaf_25_clk_i),
    .D(_00081_),
    .Q(\tx[6] ));
 sky130_fd_sc_hd__dfxtp_1 _21659_ (.CLK(clknet_leaf_25_clk_i),
    .D(_00082_),
    .Q(\tx[7] ));
 sky130_fd_sc_hd__dfxtp_1 _21660_ (.CLK(clknet_leaf_25_clk_i),
    .D(_00083_),
    .Q(\tx[8] ));
 sky130_fd_sc_hd__dfxtp_1 _21661_ (.CLK(clknet_leaf_25_clk_i),
    .D(_00084_),
    .Q(\tx[9] ));
 sky130_fd_sc_hd__dfxtp_1 _21662_ (.CLK(clknet_leaf_25_clk_i),
    .D(_00085_),
    .Q(\tx[10] ));
 sky130_fd_sc_hd__dfxtp_1 _21663_ (.CLK(clknet_leaf_24_clk_i),
    .D(_00086_),
    .Q(\tx[11] ));
 sky130_fd_sc_hd__dfxtp_1 _21664_ (.CLK(clknet_leaf_24_clk_i),
    .D(_00087_),
    .Q(\tx[12] ));
 sky130_fd_sc_hd__dfxtp_1 _21665_ (.CLK(clknet_leaf_24_clk_i),
    .D(_00088_),
    .Q(\tx[13] ));
 sky130_fd_sc_hd__dfxtp_1 _21666_ (.CLK(clknet_leaf_24_clk_i),
    .D(_00089_),
    .Q(\tx[14] ));
 sky130_fd_sc_hd__dfxtp_1 _21667_ (.CLK(clknet_leaf_24_clk_i),
    .D(_00090_),
    .Q(\tx[15] ));
 sky130_fd_sc_hd__dfxtp_1 _21668_ (.CLK(clknet_leaf_24_clk_i),
    .D(_00091_),
    .Q(\tx[16] ));
 sky130_fd_sc_hd__dfxtp_1 _21669_ (.CLK(clknet_leaf_24_clk_i),
    .D(_00092_),
    .Q(\tx[17] ));
 sky130_fd_sc_hd__dfxtp_1 _21670_ (.CLK(clknet_leaf_20_clk_i),
    .D(_00093_),
    .Q(\tx[18] ));
 sky130_fd_sc_hd__dfxtp_1 _21671_ (.CLK(clknet_leaf_24_clk_i),
    .D(_00094_),
    .Q(\tx[19] ));
 sky130_fd_sc_hd__dfxtp_1 _21672_ (.CLK(clknet_leaf_20_clk_i),
    .D(_00095_),
    .Q(\tx[20] ));
 sky130_fd_sc_hd__dfxtp_1 _21673_ (.CLK(clknet_leaf_20_clk_i),
    .D(_00096_),
    .Q(\tx[21] ));
 sky130_fd_sc_hd__dfxtp_1 _21674_ (.CLK(clknet_leaf_20_clk_i),
    .D(_00097_),
    .Q(\tx[22] ));
 sky130_fd_sc_hd__dfxtp_1 _21675_ (.CLK(clknet_leaf_20_clk_i),
    .D(_00098_),
    .Q(\tx[23] ));
 sky130_fd_sc_hd__dfxtp_1 _21676_ (.CLK(clknet_leaf_19_clk_i),
    .D(_00099_),
    .Q(\tx[24] ));
 sky130_fd_sc_hd__dfxtp_1 _21677_ (.CLK(clknet_leaf_19_clk_i),
    .D(_00100_),
    .Q(\tx[25] ));
 sky130_fd_sc_hd__dfxtp_1 _21678_ (.CLK(clknet_leaf_20_clk_i),
    .D(_00101_),
    .Q(\tx[26] ));
 sky130_fd_sc_hd__dfxtp_1 _21679_ (.CLK(clknet_leaf_19_clk_i),
    .D(_00102_),
    .Q(\tx[27] ));
 sky130_fd_sc_hd__dfxtp_1 _21680_ (.CLK(clknet_leaf_19_clk_i),
    .D(_00103_),
    .Q(\tx[28] ));
 sky130_fd_sc_hd__dfxtp_1 _21681_ (.CLK(clknet_leaf_19_clk_i),
    .D(_00104_),
    .Q(\tx[29] ));
 sky130_fd_sc_hd__dfxtp_1 _21682_ (.CLK(clknet_leaf_19_clk_i),
    .D(_00105_),
    .Q(\tx[30] ));
 sky130_fd_sc_hd__dfxtp_1 _21683_ (.CLK(clknet_leaf_20_clk_i),
    .D(_00106_),
    .Q(\tx[31] ));
 sky130_fd_sc_hd__dfxtp_1 _21684_ (.CLK(clknet_leaf_35_clk_i),
    .D(_00107_),
    .Q(\depth[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21685_ (.CLK(clknet_leaf_35_clk_i),
    .D(_00108_),
    .Q(\depth[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21686_ (.CLK(clknet_leaf_35_clk_i),
    .D(_00109_),
    .Q(\depth[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21687_ (.CLK(clknet_leaf_35_clk_i),
    .D(_00110_),
    .Q(\depth[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21688_ (.CLK(clknet_leaf_35_clk_i),
    .D(_00111_),
    .Q(\depth[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21689_ (.CLK(clknet_leaf_34_clk_i),
    .D(_00112_),
    .Q(\depth[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21690_ (.CLK(clknet_leaf_34_clk_i),
    .D(_00113_),
    .Q(\depth[6] ));
 sky130_fd_sc_hd__dfxtp_1 _21691_ (.CLK(clknet_leaf_34_clk_i),
    .D(_00114_),
    .Q(\depth[7] ));
 sky130_fd_sc_hd__dfxtp_1 _21692_ (.CLK(clknet_leaf_34_clk_i),
    .D(_00115_),
    .Q(\depth[8] ));
 sky130_fd_sc_hd__dfxtp_1 _21693_ (.CLK(clknet_leaf_34_clk_i),
    .D(_00116_),
    .Q(\depth[9] ));
 sky130_fd_sc_hd__dfxtp_1 _21694_ (.CLK(clknet_leaf_34_clk_i),
    .D(_00117_),
    .Q(\depth[10] ));
 sky130_fd_sc_hd__dfxtp_1 _21695_ (.CLK(clknet_leaf_34_clk_i),
    .D(_00118_),
    .Q(\depth[11] ));
 sky130_fd_sc_hd__dfxtp_1 _21696_ (.CLK(clknet_leaf_34_clk_i),
    .D(_00119_),
    .Q(\depth[12] ));
 sky130_fd_sc_hd__dfxtp_1 _21697_ (.CLK(clknet_leaf_34_clk_i),
    .D(_00120_),
    .Q(\depth[13] ));
 sky130_fd_sc_hd__dfxtp_1 _21698_ (.CLK(clknet_leaf_34_clk_i),
    .D(_00121_),
    .Q(\depth[14] ));
 sky130_fd_sc_hd__dfxtp_1 _21699_ (.CLK(clknet_leaf_33_clk_i),
    .D(_00122_),
    .Q(\depth[15] ));
 sky130_fd_sc_hd__dfxtp_1 _21700_ (.CLK(clknet_leaf_34_clk_i),
    .D(_00123_),
    .Q(\depth[16] ));
 sky130_fd_sc_hd__dfxtp_1 _21701_ (.CLK(clknet_leaf_33_clk_i),
    .D(_00124_),
    .Q(\depth[17] ));
 sky130_fd_sc_hd__dfxtp_1 _21702_ (.CLK(clknet_leaf_33_clk_i),
    .D(_00125_),
    .Q(\depth[18] ));
 sky130_fd_sc_hd__dfxtp_1 _21703_ (.CLK(clknet_leaf_33_clk_i),
    .D(_00126_),
    .Q(\depth[19] ));
 sky130_fd_sc_hd__dfxtp_1 _21704_ (.CLK(clknet_leaf_33_clk_i),
    .D(_00127_),
    .Q(\depth[20] ));
 sky130_fd_sc_hd__dfxtp_1 _21705_ (.CLK(clknet_leaf_33_clk_i),
    .D(_00128_),
    .Q(\depth[21] ));
 sky130_fd_sc_hd__dfxtp_1 _21706_ (.CLK(clknet_leaf_33_clk_i),
    .D(_00129_),
    .Q(\depth[22] ));
 sky130_fd_sc_hd__dfxtp_1 _21707_ (.CLK(clknet_leaf_33_clk_i),
    .D(_00130_),
    .Q(\depth[23] ));
 sky130_fd_sc_hd__dfxtp_1 _21708_ (.CLK(clknet_leaf_33_clk_i),
    .D(_00131_),
    .Q(\depth[24] ));
 sky130_fd_sc_hd__dfxtp_1 _21709_ (.CLK(clknet_leaf_33_clk_i),
    .D(_00132_),
    .Q(\depth[25] ));
 sky130_fd_sc_hd__dfxtp_1 _21710_ (.CLK(clknet_leaf_32_clk_i),
    .D(_00133_),
    .Q(\depth[26] ));
 sky130_fd_sc_hd__dfxtp_1 _21711_ (.CLK(clknet_leaf_32_clk_i),
    .D(_00134_),
    .Q(\depth[27] ));
 sky130_fd_sc_hd__dfxtp_1 _21712_ (.CLK(clknet_leaf_32_clk_i),
    .D(_00135_),
    .Q(\depth[28] ));
 sky130_fd_sc_hd__dfxtp_1 _21713_ (.CLK(clknet_leaf_32_clk_i),
    .D(_00136_),
    .Q(\depth[29] ));
 sky130_fd_sc_hd__dfxtp_1 _21714_ (.CLK(clknet_leaf_32_clk_i),
    .D(_00137_),
    .Q(\depth[30] ));
 sky130_fd_sc_hd__dfxtp_1 _21715_ (.CLK(clknet_leaf_32_clk_i),
    .D(_00138_),
    .Q(\depth[31] ));
 sky130_fd_sc_hd__dfstp_4 _21716_ (.CLK(clknet_leaf_18_clk_i),
    .D(_00001_),
    .SET_B(net645),
    .Q(sstream_o));
 sky130_fd_sc_hd__dfrtp_4 _21717_ (.CLK(clknet_leaf_25_clk_i),
    .D(net648),
    .RESET_B(net641),
    .Q(\state[1] ));
 sky130_fd_sc_hd__dfrtp_4 _21718_ (.CLK(clknet_leaf_43_clk_i),
    .D(net587),
    .RESET_B(net646),
    .Q(\state[2] ));
 sky130_fd_sc_hd__dfrtp_1 _21719_ (.CLK(clknet_leaf_1_clk_i),
    .D(net647),
    .RESET_B(net646),
    .Q(\state[3] ));
 sky130_fd_sc_hd__dfrtp_4 _21720_ (.CLK(clknet_leaf_25_clk_i),
    .D(net596),
    .RESET_B(net642),
    .Q(\state[4] ));
 sky130_fd_sc_hd__dfrtp_1 _21721_ (.CLK(clknet_leaf_1_clk_i),
    .D(_00000_),
    .RESET_B(net646),
    .Q(\state[5] ));
 sky130_fd_sc_hd__dfrtp_4 _21722_ (.CLK(clknet_leaf_18_clk_i),
    .D(_00002_),
    .RESET_B(net644),
    .Q(mstream_o[114]));
 sky130_fd_sc_hd__dfrtp_1 _21723_ (.CLK(clknet_leaf_37_clk_i),
    .D(net610),
    .RESET_B(net639),
    .Q(\state[7] ));
 sky130_fd_sc_hd__dfrtp_1 _21724_ (.CLK(clknet_leaf_43_clk_i),
    .D(net601),
    .RESET_B(net646),
    .Q(\state[8] ));
 sky130_fd_sc_hd__dfrtp_4 _21725_ (.CLK(clknet_leaf_23_clk_i),
    .D(net599),
    .RESET_B(net645),
    .Q(\state[9] ));
 sky130_fd_sc_hd__dfxtp_1 _21726_ (.CLK(clknet_leaf_2_clk_i),
    .D(_00139_),
    .Q(\mul0.a[0] ));
 sky130_fd_sc_hd__dfxtp_2 _21727_ (.CLK(clknet_leaf_2_clk_i),
    .D(_00140_),
    .Q(\mul0.a[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21728_ (.CLK(clknet_leaf_1_clk_i),
    .D(_00141_),
    .Q(\mul0.a[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21729_ (.CLK(clknet_leaf_2_clk_i),
    .D(_00142_),
    .Q(\mul0.a[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21730_ (.CLK(clknet_leaf_3_clk_i),
    .D(_00143_),
    .Q(\mul0.a[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21731_ (.CLK(clknet_leaf_3_clk_i),
    .D(_00144_),
    .Q(\mul0.a[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21732_ (.CLK(clknet_leaf_5_clk_i),
    .D(_00145_),
    .Q(\mul0.a[6] ));
 sky130_fd_sc_hd__dfxtp_4 _21733_ (.CLK(clknet_leaf_5_clk_i),
    .D(_00146_),
    .Q(\mul0.a[7] ));
 sky130_fd_sc_hd__dfxtp_4 _21734_ (.CLK(clknet_leaf_5_clk_i),
    .D(_00147_),
    .Q(\mul0.a[8] ));
 sky130_fd_sc_hd__dfxtp_4 _21735_ (.CLK(clknet_leaf_5_clk_i),
    .D(_00148_),
    .Q(\mul0.a[9] ));
 sky130_fd_sc_hd__dfxtp_1 _21736_ (.CLK(clknet_leaf_5_clk_i),
    .D(_00149_),
    .Q(\mul0.a[10] ));
 sky130_fd_sc_hd__dfxtp_2 _21737_ (.CLK(clknet_leaf_5_clk_i),
    .D(_00150_),
    .Q(\mul0.a[11] ));
 sky130_fd_sc_hd__dfxtp_2 _21738_ (.CLK(clknet_leaf_5_clk_i),
    .D(_00151_),
    .Q(\mul0.a[12] ));
 sky130_fd_sc_hd__dfxtp_1 _21739_ (.CLK(clknet_leaf_5_clk_i),
    .D(_00152_),
    .Q(\mul0.a[13] ));
 sky130_fd_sc_hd__dfxtp_4 _21740_ (.CLK(clknet_leaf_4_clk_i),
    .D(_00153_),
    .Q(\mul0.a[14] ));
 sky130_fd_sc_hd__dfxtp_4 _21741_ (.CLK(clknet_leaf_4_clk_i),
    .D(_00154_),
    .Q(\mul0.a[15] ));
 sky130_fd_sc_hd__dfxtp_4 _21742_ (.CLK(clknet_leaf_9_clk_i),
    .D(_00155_),
    .Q(\mul0.a[16] ));
 sky130_fd_sc_hd__dfxtp_4 _21743_ (.CLK(clknet_leaf_4_clk_i),
    .D(_00156_),
    .Q(\mul0.a[17] ));
 sky130_fd_sc_hd__dfxtp_2 _21744_ (.CLK(clknet_leaf_9_clk_i),
    .D(_00157_),
    .Q(\mul0.a[18] ));
 sky130_fd_sc_hd__dfxtp_2 _21745_ (.CLK(clknet_leaf_9_clk_i),
    .D(_00158_),
    .Q(\mul0.a[19] ));
 sky130_fd_sc_hd__dfxtp_2 _21746_ (.CLK(clknet_leaf_9_clk_i),
    .D(_00159_),
    .Q(\mul0.a[20] ));
 sky130_fd_sc_hd__dfxtp_4 _21747_ (.CLK(clknet_leaf_9_clk_i),
    .D(_00160_),
    .Q(\mul0.a[21] ));
 sky130_fd_sc_hd__dfxtp_4 _21748_ (.CLK(clknet_leaf_9_clk_i),
    .D(_00161_),
    .Q(\mul0.a[22] ));
 sky130_fd_sc_hd__dfxtp_1 _21749_ (.CLK(clknet_leaf_11_clk_i),
    .D(_00162_),
    .Q(\mul0.a[23] ));
 sky130_fd_sc_hd__dfxtp_1 _21750_ (.CLK(clknet_leaf_11_clk_i),
    .D(_00163_),
    .Q(\mul0.a[24] ));
 sky130_fd_sc_hd__dfxtp_1 _21751_ (.CLK(clknet_leaf_11_clk_i),
    .D(_00164_),
    .Q(\mul0.a[25] ));
 sky130_fd_sc_hd__dfxtp_1 _21752_ (.CLK(clknet_leaf_12_clk_i),
    .D(_00165_),
    .Q(\mul0.a[26] ));
 sky130_fd_sc_hd__dfxtp_2 _21753_ (.CLK(clknet_leaf_12_clk_i),
    .D(_00166_),
    .Q(\mul0.a[27] ));
 sky130_fd_sc_hd__dfxtp_2 _21754_ (.CLK(clknet_leaf_12_clk_i),
    .D(_00167_),
    .Q(\mul0.a[28] ));
 sky130_fd_sc_hd__dfxtp_4 _21755_ (.CLK(clknet_leaf_13_clk_i),
    .D(_00168_),
    .Q(\mul0.a[29] ));
 sky130_fd_sc_hd__dfxtp_1 _21756_ (.CLK(clknet_leaf_13_clk_i),
    .D(_00169_),
    .Q(\mul0.a[30] ));
 sky130_fd_sc_hd__dfxtp_2 _21757_ (.CLK(clknet_leaf_13_clk_i),
    .D(_00170_),
    .Q(\mul0.a[31] ));
 sky130_fd_sc_hd__dfxtp_1 _21758_ (.CLK(clknet_leaf_2_clk_i),
    .D(_00171_),
    .Q(\mul0.b[0] ));
 sky130_fd_sc_hd__dfxtp_4 _21759_ (.CLK(clknet_leaf_2_clk_i),
    .D(_00172_),
    .Q(\mul0.b[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21760_ (.CLK(clknet_leaf_44_clk_i),
    .D(_00173_),
    .Q(\mul0.b[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21761_ (.CLK(clknet_leaf_1_clk_i),
    .D(_00174_),
    .Q(\mul0.b[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21762_ (.CLK(clknet_leaf_44_clk_i),
    .D(_00175_),
    .Q(\mul0.b[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21763_ (.CLK(clknet_leaf_44_clk_i),
    .D(_00176_),
    .Q(\mul0.b[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21764_ (.CLK(clknet_leaf_0_clk_i),
    .D(_00177_),
    .Q(\mul0.b[6] ));
 sky130_fd_sc_hd__dfxtp_4 _21765_ (.CLK(clknet_leaf_0_clk_i),
    .D(_00178_),
    .Q(\mul0.b[7] ));
 sky130_fd_sc_hd__dfxtp_4 _21766_ (.CLK(clknet_leaf_0_clk_i),
    .D(_00179_),
    .Q(\mul0.b[8] ));
 sky130_fd_sc_hd__dfxtp_1 _21767_ (.CLK(clknet_leaf_0_clk_i),
    .D(_00180_),
    .Q(\mul0.b[9] ));
 sky130_fd_sc_hd__dfxtp_4 _21768_ (.CLK(clknet_leaf_40_clk_i),
    .D(_00181_),
    .Q(\mul0.b[10] ));
 sky130_fd_sc_hd__dfxtp_4 _21769_ (.CLK(clknet_leaf_40_clk_i),
    .D(_00182_),
    .Q(\mul0.b[11] ));
 sky130_fd_sc_hd__dfxtp_2 _21770_ (.CLK(clknet_leaf_40_clk_i),
    .D(_00183_),
    .Q(\mul0.b[12] ));
 sky130_fd_sc_hd__dfxtp_2 _21771_ (.CLK(clknet_leaf_40_clk_i),
    .D(_00184_),
    .Q(\mul0.b[13] ));
 sky130_fd_sc_hd__dfxtp_1 _21772_ (.CLK(clknet_leaf_40_clk_i),
    .D(_00185_),
    .Q(\mul0.b[14] ));
 sky130_fd_sc_hd__dfxtp_2 _21773_ (.CLK(clknet_leaf_40_clk_i),
    .D(_00186_),
    .Q(\mul0.b[15] ));
 sky130_fd_sc_hd__dfxtp_1 _21774_ (.CLK(clknet_leaf_40_clk_i),
    .D(_00187_),
    .Q(\mul0.b[16] ));
 sky130_fd_sc_hd__dfxtp_2 _21775_ (.CLK(clknet_leaf_6_clk_i),
    .D(_00188_),
    .Q(\mul0.b[17] ));
 sky130_fd_sc_hd__dfxtp_4 _21776_ (.CLK(clknet_2_0__leaf_clk_i),
    .D(_00189_),
    .Q(\mul0.b[18] ));
 sky130_fd_sc_hd__dfxtp_2 _21777_ (.CLK(clknet_leaf_6_clk_i),
    .D(_00190_),
    .Q(\mul0.b[19] ));
 sky130_fd_sc_hd__dfxtp_1 _21778_ (.CLK(clknet_leaf_7_clk_i),
    .D(_00191_),
    .Q(\mul0.b[20] ));
 sky130_fd_sc_hd__dfxtp_1 _21779_ (.CLK(clknet_leaf_40_clk_i),
    .D(_00192_),
    .Q(\mul0.b[21] ));
 sky130_fd_sc_hd__dfxtp_1 _21780_ (.CLK(clknet_leaf_6_clk_i),
    .D(_00193_),
    .Q(\mul0.b[22] ));
 sky130_fd_sc_hd__dfxtp_2 _21781_ (.CLK(clknet_leaf_14_clk_i),
    .D(_00194_),
    .Q(\mul0.b[23] ));
 sky130_fd_sc_hd__dfxtp_1 _21782_ (.CLK(clknet_leaf_14_clk_i),
    .D(_00195_),
    .Q(\mul0.b[24] ));
 sky130_fd_sc_hd__dfxtp_1 _21783_ (.CLK(clknet_leaf_14_clk_i),
    .D(_00196_),
    .Q(\mul0.b[25] ));
 sky130_fd_sc_hd__dfxtp_2 _21784_ (.CLK(clknet_leaf_14_clk_i),
    .D(_00197_),
    .Q(\mul0.b[26] ));
 sky130_fd_sc_hd__dfxtp_1 _21785_ (.CLK(clknet_leaf_16_clk_i),
    .D(_00198_),
    .Q(\mul0.b[27] ));
 sky130_fd_sc_hd__dfxtp_1 _21786_ (.CLK(clknet_leaf_16_clk_i),
    .D(_00199_),
    .Q(\mul0.b[28] ));
 sky130_fd_sc_hd__dfxtp_2 _21787_ (.CLK(clknet_leaf_16_clk_i),
    .D(_00200_),
    .Q(\mul0.b[29] ));
 sky130_fd_sc_hd__dfxtp_2 _21788_ (.CLK(clknet_leaf_16_clk_i),
    .D(_00201_),
    .Q(\mul0.b[30] ));
 sky130_fd_sc_hd__dfxtp_4 _21789_ (.CLK(clknet_leaf_40_clk_i),
    .D(_00202_),
    .Q(\mul0.b[31] ));
 sky130_fd_sc_hd__dfxtp_1 _21790_ (.CLK(clknet_leaf_44_clk_i),
    .D(_00203_),
    .Q(\mul1.a[0] ));
 sky130_fd_sc_hd__dfxtp_4 _21791_ (.CLK(clknet_leaf_1_clk_i),
    .D(_00204_),
    .Q(\mul1.a[1] ));
 sky130_fd_sc_hd__dfxtp_4 _21792_ (.CLK(clknet_leaf_1_clk_i),
    .D(_00205_),
    .Q(\mul1.a[2] ));
 sky130_fd_sc_hd__dfxtp_4 _21793_ (.CLK(clknet_leaf_2_clk_i),
    .D(_00206_),
    .Q(\mul1.a[3] ));
 sky130_fd_sc_hd__dfxtp_4 _21794_ (.CLK(clknet_leaf_2_clk_i),
    .D(_00207_),
    .Q(\mul1.a[4] ));
 sky130_fd_sc_hd__dfxtp_4 _21795_ (.CLK(clknet_leaf_3_clk_i),
    .D(_00208_),
    .Q(\mul1.a[5] ));
 sky130_fd_sc_hd__dfxtp_4 _21796_ (.CLK(clknet_leaf_5_clk_i),
    .D(_00209_),
    .Q(\mul1.a[6] ));
 sky130_fd_sc_hd__dfxtp_1 _21797_ (.CLK(clknet_leaf_5_clk_i),
    .D(_00210_),
    .Q(\mul1.a[7] ));
 sky130_fd_sc_hd__dfxtp_2 _21798_ (.CLK(clknet_leaf_5_clk_i),
    .D(_00211_),
    .Q(\mul1.a[8] ));
 sky130_fd_sc_hd__dfxtp_4 _21799_ (.CLK(clknet_leaf_5_clk_i),
    .D(_00212_),
    .Q(\mul1.a[9] ));
 sky130_fd_sc_hd__dfxtp_4 _21800_ (.CLK(clknet_leaf_5_clk_i),
    .D(_00213_),
    .Q(\mul1.a[10] ));
 sky130_fd_sc_hd__dfxtp_1 _21801_ (.CLK(clknet_leaf_5_clk_i),
    .D(_00214_),
    .Q(\mul1.a[11] ));
 sky130_fd_sc_hd__dfxtp_4 _21802_ (.CLK(clknet_leaf_5_clk_i),
    .D(_00215_),
    .Q(\mul1.a[12] ));
 sky130_fd_sc_hd__dfxtp_2 _21803_ (.CLK(clknet_leaf_5_clk_i),
    .D(_00216_),
    .Q(\mul1.a[13] ));
 sky130_fd_sc_hd__dfxtp_1 _21804_ (.CLK(clknet_leaf_4_clk_i),
    .D(_00217_),
    .Q(\mul1.a[14] ));
 sky130_fd_sc_hd__dfxtp_1 _21805_ (.CLK(clknet_leaf_4_clk_i),
    .D(_00218_),
    .Q(\mul1.a[15] ));
 sky130_fd_sc_hd__dfxtp_1 _21806_ (.CLK(clknet_2_1__leaf_clk_i),
    .D(_00219_),
    .Q(\mul1.a[16] ));
 sky130_fd_sc_hd__dfxtp_2 _21807_ (.CLK(clknet_leaf_6_clk_i),
    .D(_00220_),
    .Q(\mul1.a[17] ));
 sky130_fd_sc_hd__dfxtp_1 _21808_ (.CLK(clknet_leaf_6_clk_i),
    .D(_00221_),
    .Q(\mul1.a[18] ));
 sky130_fd_sc_hd__dfxtp_1 _21809_ (.CLK(clknet_leaf_6_clk_i),
    .D(_00222_),
    .Q(\mul1.a[19] ));
 sky130_fd_sc_hd__dfxtp_1 _21810_ (.CLK(clknet_leaf_7_clk_i),
    .D(_00223_),
    .Q(\mul1.a[20] ));
 sky130_fd_sc_hd__dfxtp_1 _21811_ (.CLK(clknet_leaf_7_clk_i),
    .D(_00224_),
    .Q(\mul1.a[21] ));
 sky130_fd_sc_hd__dfxtp_1 _21812_ (.CLK(clknet_leaf_7_clk_i),
    .D(_00225_),
    .Q(\mul1.a[22] ));
 sky130_fd_sc_hd__dfxtp_1 _21813_ (.CLK(clknet_leaf_7_clk_i),
    .D(_00226_),
    .Q(\mul1.a[23] ));
 sky130_fd_sc_hd__dfxtp_1 _21814_ (.CLK(clknet_leaf_7_clk_i),
    .D(_00227_),
    .Q(\mul1.a[24] ));
 sky130_fd_sc_hd__dfxtp_4 _21815_ (.CLK(clknet_leaf_15_clk_i),
    .D(_00228_),
    .Q(\mul1.a[25] ));
 sky130_fd_sc_hd__dfxtp_4 _21816_ (.CLK(clknet_leaf_7_clk_i),
    .D(_00229_),
    .Q(\mul1.a[26] ));
 sky130_fd_sc_hd__dfxtp_2 _21817_ (.CLK(clknet_leaf_15_clk_i),
    .D(_00230_),
    .Q(\mul1.a[27] ));
 sky130_fd_sc_hd__dfxtp_1 _21818_ (.CLK(clknet_leaf_14_clk_i),
    .D(_00231_),
    .Q(\mul1.a[28] ));
 sky130_fd_sc_hd__dfxtp_2 _21819_ (.CLK(clknet_leaf_14_clk_i),
    .D(_00232_),
    .Q(\mul1.a[29] ));
 sky130_fd_sc_hd__dfxtp_2 _21820_ (.CLK(clknet_leaf_14_clk_i),
    .D(_00233_),
    .Q(\mul1.a[30] ));
 sky130_fd_sc_hd__dfxtp_1 _21821_ (.CLK(clknet_leaf_14_clk_i),
    .D(_00234_),
    .Q(\mul1.a[31] ));
 sky130_fd_sc_hd__dfxtp_2 _21822_ (.CLK(clknet_2_0__leaf_clk_i),
    .D(_00235_),
    .Q(\mul1.b[0] ));
 sky130_fd_sc_hd__dfxtp_2 _21823_ (.CLK(clknet_leaf_41_clk_i),
    .D(_00236_),
    .Q(\mul1.b[1] ));
 sky130_fd_sc_hd__dfxtp_4 _21824_ (.CLK(clknet_leaf_41_clk_i),
    .D(_00237_),
    .Q(\mul1.b[2] ));
 sky130_fd_sc_hd__dfxtp_4 _21825_ (.CLK(clknet_leaf_41_clk_i),
    .D(_00238_),
    .Q(\mul1.b[3] ));
 sky130_fd_sc_hd__dfxtp_2 _21826_ (.CLK(clknet_leaf_41_clk_i),
    .D(_00239_),
    .Q(\mul1.b[4] ));
 sky130_fd_sc_hd__dfxtp_2 _21827_ (.CLK(clknet_leaf_41_clk_i),
    .D(_00240_),
    .Q(\mul1.b[5] ));
 sky130_fd_sc_hd__dfxtp_2 _21828_ (.CLK(clknet_leaf_41_clk_i),
    .D(_00241_),
    .Q(\mul1.b[6] ));
 sky130_fd_sc_hd__dfxtp_2 _21829_ (.CLK(clknet_leaf_41_clk_i),
    .D(_00242_),
    .Q(\mul1.b[7] ));
 sky130_fd_sc_hd__dfxtp_4 _21830_ (.CLK(clknet_leaf_38_clk_i),
    .D(_00243_),
    .Q(\mul1.b[8] ));
 sky130_fd_sc_hd__dfxtp_2 _21831_ (.CLK(clknet_leaf_38_clk_i),
    .D(_00244_),
    .Q(\mul1.b[9] ));
 sky130_fd_sc_hd__dfxtp_2 _21832_ (.CLK(clknet_leaf_38_clk_i),
    .D(_00245_),
    .Q(\mul1.b[10] ));
 sky130_fd_sc_hd__dfxtp_4 _21833_ (.CLK(clknet_leaf_38_clk_i),
    .D(_00246_),
    .Q(\mul1.b[11] ));
 sky130_fd_sc_hd__dfxtp_1 _21834_ (.CLK(clknet_leaf_38_clk_i),
    .D(_00247_),
    .Q(\mul1.b[12] ));
 sky130_fd_sc_hd__dfxtp_1 _21835_ (.CLK(clknet_leaf_38_clk_i),
    .D(_00248_),
    .Q(\mul1.b[13] ));
 sky130_fd_sc_hd__dfxtp_1 _21836_ (.CLK(clknet_leaf_38_clk_i),
    .D(_00249_),
    .Q(\mul1.b[14] ));
 sky130_fd_sc_hd__dfxtp_1 _21837_ (.CLK(clknet_leaf_38_clk_i),
    .D(_00250_),
    .Q(\mul1.b[15] ));
 sky130_fd_sc_hd__dfxtp_1 _21838_ (.CLK(clknet_leaf_37_clk_i),
    .D(_00251_),
    .Q(\mul1.b[16] ));
 sky130_fd_sc_hd__dfxtp_4 _21839_ (.CLK(clknet_leaf_37_clk_i),
    .D(_00252_),
    .Q(\mul1.b[17] ));
 sky130_fd_sc_hd__dfxtp_1 _21840_ (.CLK(clknet_leaf_37_clk_i),
    .D(_00253_),
    .Q(\mul1.b[18] ));
 sky130_fd_sc_hd__dfxtp_4 _21841_ (.CLK(clknet_leaf_37_clk_i),
    .D(_00254_),
    .Q(\mul1.b[19] ));
 sky130_fd_sc_hd__dfxtp_4 _21842_ (.CLK(clknet_leaf_37_clk_i),
    .D(_00255_),
    .Q(\mul1.b[20] ));
 sky130_fd_sc_hd__dfxtp_2 _21843_ (.CLK(clknet_leaf_37_clk_i),
    .D(_00256_),
    .Q(\mul1.b[21] ));
 sky130_fd_sc_hd__dfxtp_2 _21844_ (.CLK(clknet_leaf_37_clk_i),
    .D(_00257_),
    .Q(\mul1.b[22] ));
 sky130_fd_sc_hd__dfxtp_1 _21845_ (.CLK(clknet_leaf_37_clk_i),
    .D(_00258_),
    .Q(\mul1.b[23] ));
 sky130_fd_sc_hd__dfxtp_1 _21846_ (.CLK(clknet_leaf_36_clk_i),
    .D(_00259_),
    .Q(\mul1.b[24] ));
 sky130_fd_sc_hd__dfxtp_4 _21847_ (.CLK(clknet_leaf_36_clk_i),
    .D(_00260_),
    .Q(\mul1.b[25] ));
 sky130_fd_sc_hd__dfxtp_2 _21848_ (.CLK(clknet_leaf_36_clk_i),
    .D(_00261_),
    .Q(\mul1.b[26] ));
 sky130_fd_sc_hd__dfxtp_1 _21849_ (.CLK(clknet_leaf_36_clk_i),
    .D(_00262_),
    .Q(\mul1.b[27] ));
 sky130_fd_sc_hd__dfxtp_1 _21850_ (.CLK(clknet_leaf_36_clk_i),
    .D(_00263_),
    .Q(\mul1.b[28] ));
 sky130_fd_sc_hd__dfxtp_1 _21851_ (.CLK(clknet_leaf_36_clk_i),
    .D(_00264_),
    .Q(\mul1.b[29] ));
 sky130_fd_sc_hd__dfxtp_1 _21852_ (.CLK(clknet_leaf_36_clk_i),
    .D(_00265_),
    .Q(\mul1.b[30] ));
 sky130_fd_sc_hd__dfxtp_4 _21853_ (.CLK(clknet_leaf_36_clk_i),
    .D(_00266_),
    .Q(\mul1.b[31] ));
 sky130_fd_sc_hd__dfxtp_1 _21854_ (.CLK(clknet_leaf_31_clk_i),
    .D(_00267_),
    .Q(\add0.a_i[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21855_ (.CLK(clknet_leaf_27_clk_i),
    .D(_00268_),
    .Q(\add0.a_i[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21856_ (.CLK(clknet_leaf_26_clk_i),
    .D(net760),
    .Q(\add0.a_i[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21857_ (.CLK(clknet_leaf_27_clk_i),
    .D(net721),
    .Q(\add0.a_i[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21858_ (.CLK(clknet_leaf_28_clk_i),
    .D(_00271_),
    .Q(\add0.a_i[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21859_ (.CLK(clknet_leaf_27_clk_i),
    .D(_00272_),
    .Q(\add0.a_i[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21860_ (.CLK(clknet_leaf_29_clk_i),
    .D(_00273_),
    .Q(\add0.a_i[6] ));
 sky130_fd_sc_hd__dfxtp_1 _21861_ (.CLK(clknet_leaf_29_clk_i),
    .D(net754),
    .Q(\add0.a_i[7] ));
 sky130_fd_sc_hd__dfxtp_1 _21862_ (.CLK(clknet_leaf_29_clk_i),
    .D(_00275_),
    .Q(\add0.a_i[8] ));
 sky130_fd_sc_hd__dfxtp_1 _21863_ (.CLK(clknet_leaf_29_clk_i),
    .D(_00276_),
    .Q(\add0.a_i[9] ));
 sky130_fd_sc_hd__dfxtp_1 _21864_ (.CLK(clknet_leaf_29_clk_i),
    .D(_00277_),
    .Q(\add0.a_i[10] ));
 sky130_fd_sc_hd__dfxtp_1 _21865_ (.CLK(clknet_leaf_30_clk_i),
    .D(_00278_),
    .Q(\add0.a_i[11] ));
 sky130_fd_sc_hd__dfxtp_1 _21866_ (.CLK(clknet_leaf_30_clk_i),
    .D(net676),
    .Q(\add0.a_i[12] ));
 sky130_fd_sc_hd__dfxtp_1 _21867_ (.CLK(clknet_leaf_22_clk_i),
    .D(_00280_),
    .Q(\add0.a_i[13] ));
 sky130_fd_sc_hd__dfxtp_1 _21868_ (.CLK(clknet_leaf_22_clk_i),
    .D(net787),
    .Q(\add0.a_i[14] ));
 sky130_fd_sc_hd__dfxtp_1 _21869_ (.CLK(clknet_leaf_22_clk_i),
    .D(_00282_),
    .Q(\add0.a_i[15] ));
 sky130_fd_sc_hd__dfxtp_1 _21870_ (.CLK(clknet_leaf_25_clk_i),
    .D(_00283_),
    .Q(\add0.a_i[16] ));
 sky130_fd_sc_hd__dfxtp_1 _21871_ (.CLK(clknet_leaf_25_clk_i),
    .D(_00284_),
    .Q(\add0.a_i[17] ));
 sky130_fd_sc_hd__dfxtp_1 _21872_ (.CLK(clknet_leaf_23_clk_i),
    .D(net730),
    .Q(\add0.a_i[18] ));
 sky130_fd_sc_hd__dfxtp_1 _21873_ (.CLK(clknet_leaf_23_clk_i),
    .D(net749),
    .Q(\add0.a_i[19] ));
 sky130_fd_sc_hd__dfxtp_1 _21874_ (.CLK(clknet_leaf_24_clk_i),
    .D(_00287_),
    .Q(\add0.a_i[20] ));
 sky130_fd_sc_hd__dfxtp_1 _21875_ (.CLK(clknet_leaf_20_clk_i),
    .D(_00288_),
    .Q(\add0.a_i[21] ));
 sky130_fd_sc_hd__dfxtp_1 _21876_ (.CLK(clknet_leaf_21_clk_i),
    .D(net756),
    .Q(\add0.a_i[22] ));
 sky130_fd_sc_hd__dfxtp_1 _21877_ (.CLK(clknet_leaf_22_clk_i),
    .D(_00290_),
    .Q(\add0.a_i[23] ));
 sky130_fd_sc_hd__dfxtp_1 _21878_ (.CLK(clknet_leaf_21_clk_i),
    .D(_00291_),
    .Q(\add0.a_i[24] ));
 sky130_fd_sc_hd__dfxtp_2 _21879_ (.CLK(clknet_leaf_21_clk_i),
    .D(_00292_),
    .Q(\add0.a_i[25] ));
 sky130_fd_sc_hd__dfxtp_1 _21880_ (.CLK(clknet_leaf_21_clk_i),
    .D(_00293_),
    .Q(\add0.a_i[26] ));
 sky130_fd_sc_hd__dfxtp_1 _21881_ (.CLK(clknet_leaf_21_clk_i),
    .D(net683),
    .Q(\add0.a_i[27] ));
 sky130_fd_sc_hd__dfxtp_1 _21882_ (.CLK(clknet_leaf_17_clk_i),
    .D(_00295_),
    .Q(\add0.a_i[28] ));
 sky130_fd_sc_hd__dfxtp_1 _21883_ (.CLK(clknet_leaf_17_clk_i),
    .D(net775),
    .Q(\add0.a_i[29] ));
 sky130_fd_sc_hd__dfxtp_1 _21884_ (.CLK(clknet_leaf_30_clk_i),
    .D(net739),
    .Q(\add0.a_i[30] ));
 sky130_fd_sc_hd__dfxtp_1 _21885_ (.CLK(clknet_leaf_21_clk_i),
    .D(_00298_),
    .Q(\add0.a_i[31] ));
 sky130_fd_sc_hd__dfxtp_1 _21886_ (.CLK(clknet_leaf_28_clk_i),
    .D(_00299_),
    .Q(\add0.b_i[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21887_ (.CLK(clknet_leaf_31_clk_i),
    .D(_00300_),
    .Q(\add0.b_i[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21888_ (.CLK(clknet_leaf_26_clk_i),
    .D(net781),
    .Q(\add0.b_i[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21889_ (.CLK(clknet_leaf_27_clk_i),
    .D(net737),
    .Q(\add0.b_i[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21890_ (.CLK(clknet_leaf_28_clk_i),
    .D(_00303_),
    .Q(\add0.b_i[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21891_ (.CLK(clknet_leaf_27_clk_i),
    .D(_00304_),
    .Q(\add0.b_i[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21892_ (.CLK(clknet_leaf_28_clk_i),
    .D(_00305_),
    .Q(\add0.b_i[6] ));
 sky130_fd_sc_hd__dfxtp_1 _21893_ (.CLK(clknet_leaf_29_clk_i),
    .D(net751),
    .Q(\add0.b_i[7] ));
 sky130_fd_sc_hd__dfxtp_1 _21894_ (.CLK(clknet_leaf_23_clk_i),
    .D(_00307_),
    .Q(\add0.b_i[8] ));
 sky130_fd_sc_hd__dfxtp_1 _21895_ (.CLK(clknet_leaf_29_clk_i),
    .D(_00308_),
    .Q(\add0.b_i[9] ));
 sky130_fd_sc_hd__dfxtp_1 _21896_ (.CLK(clknet_leaf_29_clk_i),
    .D(net681),
    .Q(\add0.b_i[10] ));
 sky130_fd_sc_hd__dfxtp_1 _21897_ (.CLK(clknet_leaf_29_clk_i),
    .D(_00310_),
    .Q(\add0.b_i[11] ));
 sky130_fd_sc_hd__dfxtp_1 _21898_ (.CLK(clknet_leaf_30_clk_i),
    .D(net669),
    .Q(\add0.b_i[12] ));
 sky130_fd_sc_hd__dfxtp_1 _21899_ (.CLK(clknet_leaf_22_clk_i),
    .D(_00312_),
    .Q(\add0.b_i[13] ));
 sky130_fd_sc_hd__dfxtp_1 _21900_ (.CLK(clknet_leaf_22_clk_i),
    .D(net744),
    .Q(\add0.b_i[14] ));
 sky130_fd_sc_hd__dfxtp_1 _21901_ (.CLK(clknet_leaf_22_clk_i),
    .D(_00314_),
    .Q(\add0.b_i[15] ));
 sky130_fd_sc_hd__dfxtp_1 _21902_ (.CLK(clknet_leaf_25_clk_i),
    .D(net899),
    .Q(\add0.b_i[16] ));
 sky130_fd_sc_hd__dfxtp_1 _21903_ (.CLK(clknet_leaf_23_clk_i),
    .D(net864),
    .Q(\add0.b_i[17] ));
 sky130_fd_sc_hd__dfxtp_1 _21904_ (.CLK(clknet_leaf_23_clk_i),
    .D(net784),
    .Q(\add0.b_i[18] ));
 sky130_fd_sc_hd__dfxtp_1 _21905_ (.CLK(clknet_leaf_23_clk_i),
    .D(net773),
    .Q(\add0.b_i[19] ));
 sky130_fd_sc_hd__dfxtp_1 _21906_ (.CLK(clknet_leaf_24_clk_i),
    .D(_00319_),
    .Q(\add0.b_i[20] ));
 sky130_fd_sc_hd__dfxtp_1 _21907_ (.CLK(clknet_leaf_20_clk_i),
    .D(_00320_),
    .Q(\add0.b_i[21] ));
 sky130_fd_sc_hd__dfxtp_1 _21908_ (.CLK(clknet_leaf_21_clk_i),
    .D(net805),
    .Q(\add0.b_i[22] ));
 sky130_fd_sc_hd__dfxtp_1 _21909_ (.CLK(clknet_leaf_22_clk_i),
    .D(_00322_),
    .Q(\add0.b_i[23] ));
 sky130_fd_sc_hd__dfxtp_1 _21910_ (.CLK(clknet_leaf_21_clk_i),
    .D(_00323_),
    .Q(\add0.b_i[24] ));
 sky130_fd_sc_hd__dfxtp_2 _21911_ (.CLK(clknet_leaf_21_clk_i),
    .D(_00324_),
    .Q(\add0.b_i[25] ));
 sky130_fd_sc_hd__dfxtp_1 _21912_ (.CLK(clknet_leaf_21_clk_i),
    .D(_00325_),
    .Q(\add0.b_i[26] ));
 sky130_fd_sc_hd__dfxtp_1 _21913_ (.CLK(clknet_leaf_21_clk_i),
    .D(_00326_),
    .Q(\add0.b_i[27] ));
 sky130_fd_sc_hd__dfxtp_1 _21914_ (.CLK(clknet_leaf_17_clk_i),
    .D(_00327_),
    .Q(\add0.b_i[28] ));
 sky130_fd_sc_hd__dfxtp_1 _21915_ (.CLK(clknet_leaf_17_clk_i),
    .D(net793),
    .Q(\add0.b_i[29] ));
 sky130_fd_sc_hd__dfxtp_1 _21916_ (.CLK(clknet_leaf_30_clk_i),
    .D(net818),
    .Q(\add0.b_i[30] ));
 sky130_fd_sc_hd__dfxtp_1 _21917_ (.CLK(clknet_leaf_30_clk_i),
    .D(_00330_),
    .Q(\add0.b_i[31] ));
 sky130_fd_sc_hd__dfxtp_1 _21918_ (.CLK(clknet_leaf_28_clk_i),
    .D(_00331_),
    .Q(\temp[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21919_ (.CLK(clknet_leaf_31_clk_i),
    .D(_00332_),
    .Q(\temp[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21920_ (.CLK(clknet_leaf_27_clk_i),
    .D(_00333_),
    .Q(\temp[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21921_ (.CLK(clknet_leaf_27_clk_i),
    .D(_00334_),
    .Q(\temp[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21922_ (.CLK(clknet_leaf_28_clk_i),
    .D(_00335_),
    .Q(\temp[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21923_ (.CLK(clknet_leaf_27_clk_i),
    .D(_00336_),
    .Q(\temp[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21924_ (.CLK(clknet_leaf_28_clk_i),
    .D(_00337_),
    .Q(\temp[6] ));
 sky130_fd_sc_hd__dfxtp_1 _21925_ (.CLK(clknet_leaf_29_clk_i),
    .D(_00338_),
    .Q(\temp[7] ));
 sky130_fd_sc_hd__dfxtp_1 _21926_ (.CLK(clknet_leaf_28_clk_i),
    .D(_00339_),
    .Q(\temp[8] ));
 sky130_fd_sc_hd__dfxtp_1 _21927_ (.CLK(clknet_leaf_29_clk_i),
    .D(_00340_),
    .Q(\temp[9] ));
 sky130_fd_sc_hd__dfxtp_1 _21928_ (.CLK(clknet_leaf_29_clk_i),
    .D(_00341_),
    .Q(\temp[10] ));
 sky130_fd_sc_hd__dfxtp_1 _21929_ (.CLK(clknet_leaf_29_clk_i),
    .D(_00342_),
    .Q(\temp[11] ));
 sky130_fd_sc_hd__dfxtp_1 _21930_ (.CLK(clknet_leaf_30_clk_i),
    .D(_00343_),
    .Q(\temp[12] ));
 sky130_fd_sc_hd__dfxtp_1 _21931_ (.CLK(clknet_leaf_22_clk_i),
    .D(_00344_),
    .Q(\temp[13] ));
 sky130_fd_sc_hd__dfxtp_1 _21932_ (.CLK(clknet_leaf_29_clk_i),
    .D(_00345_),
    .Q(\temp[14] ));
 sky130_fd_sc_hd__dfxtp_1 _21933_ (.CLK(clknet_leaf_22_clk_i),
    .D(_00346_),
    .Q(\temp[15] ));
 sky130_fd_sc_hd__dfxtp_1 _21934_ (.CLK(clknet_leaf_25_clk_i),
    .D(_00347_),
    .Q(\temp[16] ));
 sky130_fd_sc_hd__dfxtp_1 _21935_ (.CLK(clknet_leaf_23_clk_i),
    .D(_00348_),
    .Q(\temp[17] ));
 sky130_fd_sc_hd__dfxtp_1 _21936_ (.CLK(clknet_leaf_23_clk_i),
    .D(_00349_),
    .Q(\temp[18] ));
 sky130_fd_sc_hd__dfxtp_1 _21937_ (.CLK(clknet_leaf_22_clk_i),
    .D(_00350_),
    .Q(\temp[19] ));
 sky130_fd_sc_hd__dfxtp_1 _21938_ (.CLK(clknet_leaf_23_clk_i),
    .D(_00351_),
    .Q(\temp[20] ));
 sky130_fd_sc_hd__dfxtp_1 _21939_ (.CLK(clknet_leaf_20_clk_i),
    .D(_00352_),
    .Q(\temp[21] ));
 sky130_fd_sc_hd__dfxtp_1 _21940_ (.CLK(clknet_leaf_22_clk_i),
    .D(_00353_),
    .Q(\temp[22] ));
 sky130_fd_sc_hd__dfxtp_1 _21941_ (.CLK(clknet_leaf_22_clk_i),
    .D(_00354_),
    .Q(\temp[23] ));
 sky130_fd_sc_hd__dfxtp_1 _21942_ (.CLK(clknet_leaf_22_clk_i),
    .D(_00355_),
    .Q(\temp[24] ));
 sky130_fd_sc_hd__dfxtp_1 _21943_ (.CLK(clknet_leaf_21_clk_i),
    .D(_00356_),
    .Q(\temp[25] ));
 sky130_fd_sc_hd__dfxtp_1 _21944_ (.CLK(clknet_leaf_21_clk_i),
    .D(_00357_),
    .Q(\temp[26] ));
 sky130_fd_sc_hd__dfxtp_1 _21945_ (.CLK(clknet_leaf_21_clk_i),
    .D(_00358_),
    .Q(\temp[27] ));
 sky130_fd_sc_hd__dfxtp_1 _21946_ (.CLK(clknet_leaf_17_clk_i),
    .D(_00359_),
    .Q(\temp[28] ));
 sky130_fd_sc_hd__dfxtp_1 _21947_ (.CLK(clknet_leaf_17_clk_i),
    .D(_00360_),
    .Q(\temp[29] ));
 sky130_fd_sc_hd__dfxtp_1 _21948_ (.CLK(clknet_leaf_30_clk_i),
    .D(_00361_),
    .Q(\temp[30] ));
 sky130_fd_sc_hd__dfxtp_1 _21949_ (.CLK(clknet_leaf_17_clk_i),
    .D(_00362_),
    .Q(\temp[31] ));
 sky130_fd_sc_hd__dfxtp_1 _21950_ (.CLK(clknet_leaf_44_clk_i),
    .D(_00363_),
    .Q(\in_data[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21951_ (.CLK(clknet_leaf_44_clk_i),
    .D(_00364_),
    .Q(\in_data[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21952_ (.CLK(clknet_leaf_44_clk_i),
    .D(_00365_),
    .Q(\in_data[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21953_ (.CLK(clknet_leaf_44_clk_i),
    .D(_00366_),
    .Q(\in_data[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21954_ (.CLK(clknet_leaf_44_clk_i),
    .D(_00367_),
    .Q(\in_data[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21955_ (.CLK(clknet_leaf_44_clk_i),
    .D(_00368_),
    .Q(\in_data[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21956_ (.CLK(clknet_leaf_44_clk_i),
    .D(_00369_),
    .Q(\in_data[6] ));
 sky130_fd_sc_hd__dfxtp_1 _21957_ (.CLK(clknet_leaf_44_clk_i),
    .D(_00370_),
    .Q(\in_data[7] ));
 sky130_fd_sc_hd__dfxtp_1 _21958_ (.CLK(clknet_leaf_44_clk_i),
    .D(_00371_),
    .Q(\in_data[8] ));
 sky130_fd_sc_hd__dfxtp_1 _21959_ (.CLK(clknet_leaf_44_clk_i),
    .D(_00372_),
    .Q(\in_data[9] ));
 sky130_fd_sc_hd__dfxtp_1 _21960_ (.CLK(clknet_leaf_44_clk_i),
    .D(_00373_),
    .Q(\in_data[10] ));
 sky130_fd_sc_hd__dfxtp_1 _21961_ (.CLK(clknet_leaf_44_clk_i),
    .D(_00374_),
    .Q(\in_data[11] ));
 sky130_fd_sc_hd__dfxtp_1 _21962_ (.CLK(clknet_leaf_44_clk_i),
    .D(_00375_),
    .Q(\in_data[12] ));
 sky130_fd_sc_hd__dfxtp_1 _21963_ (.CLK(clknet_leaf_44_clk_i),
    .D(_00376_),
    .Q(\in_data[13] ));
 sky130_fd_sc_hd__dfxtp_1 _21964_ (.CLK(clknet_leaf_1_clk_i),
    .D(_00377_),
    .Q(\in_data[14] ));
 sky130_fd_sc_hd__dfxtp_1 _21965_ (.CLK(clknet_leaf_1_clk_i),
    .D(_00378_),
    .Q(\in_data[15] ));
 sky130_fd_sc_hd__dfxtp_1 _21966_ (.CLK(clknet_leaf_1_clk_i),
    .D(_00379_),
    .Q(\in_data[16] ));
 sky130_fd_sc_hd__dfxtp_1 _21967_ (.CLK(clknet_leaf_1_clk_i),
    .D(_00380_),
    .Q(\in_data[17] ));
 sky130_fd_sc_hd__dfxtp_1 _21968_ (.CLK(clknet_leaf_1_clk_i),
    .D(_00381_),
    .Q(\in_data[18] ));
 sky130_fd_sc_hd__dfxtp_1 _21969_ (.CLK(clknet_leaf_1_clk_i),
    .D(_00382_),
    .Q(\in_data[19] ));
 sky130_fd_sc_hd__dfxtp_1 _21970_ (.CLK(clknet_leaf_1_clk_i),
    .D(_00383_),
    .Q(\in_data[20] ));
 sky130_fd_sc_hd__dfxtp_1 _21971_ (.CLK(clknet_leaf_1_clk_i),
    .D(_00384_),
    .Q(\in_data[21] ));
 sky130_fd_sc_hd__dfxtp_1 _21972_ (.CLK(clknet_leaf_1_clk_i),
    .D(_00385_),
    .Q(\in_data[22] ));
 sky130_fd_sc_hd__dfxtp_1 _21973_ (.CLK(clknet_leaf_2_clk_i),
    .D(_00386_),
    .Q(\in_data[23] ));
 sky130_fd_sc_hd__dfxtp_1 _21974_ (.CLK(clknet_leaf_1_clk_i),
    .D(_00387_),
    .Q(\in_data[24] ));
 sky130_fd_sc_hd__dfxtp_1 _21975_ (.CLK(clknet_leaf_2_clk_i),
    .D(_00388_),
    .Q(\in_data[25] ));
 sky130_fd_sc_hd__dfxtp_1 _21976_ (.CLK(clknet_leaf_10_clk_i),
    .D(_00389_),
    .Q(\in_data[26] ));
 sky130_fd_sc_hd__dfxtp_1 _21977_ (.CLK(clknet_leaf_4_clk_i),
    .D(_00390_),
    .Q(\in_data[27] ));
 sky130_fd_sc_hd__dfxtp_1 _21978_ (.CLK(clknet_leaf_9_clk_i),
    .D(_00391_),
    .Q(\in_data[28] ));
 sky130_fd_sc_hd__dfxtp_1 _21979_ (.CLK(clknet_leaf_10_clk_i),
    .D(_00392_),
    .Q(\in_data[29] ));
 sky130_fd_sc_hd__dfxtp_1 _21980_ (.CLK(clknet_leaf_10_clk_i),
    .D(_00393_),
    .Q(\in_data[30] ));
 sky130_fd_sc_hd__dfxtp_1 _21981_ (.CLK(clknet_leaf_10_clk_i),
    .D(_00394_),
    .Q(\in_data[31] ));
 sky130_fd_sc_hd__dfxtp_1 _21982_ (.CLK(clknet_leaf_2_clk_i),
    .D(_00395_),
    .Q(\in_data[32] ));
 sky130_fd_sc_hd__dfxtp_1 _21983_ (.CLK(clknet_leaf_2_clk_i),
    .D(_00396_),
    .Q(\in_data[33] ));
 sky130_fd_sc_hd__dfxtp_1 _21984_ (.CLK(clknet_leaf_2_clk_i),
    .D(_00397_),
    .Q(\in_data[34] ));
 sky130_fd_sc_hd__dfxtp_1 _21985_ (.CLK(clknet_leaf_3_clk_i),
    .D(_00398_),
    .Q(\in_data[35] ));
 sky130_fd_sc_hd__dfxtp_1 _21986_ (.CLK(clknet_leaf_3_clk_i),
    .D(_00399_),
    .Q(\in_data[36] ));
 sky130_fd_sc_hd__dfxtp_1 _21987_ (.CLK(clknet_leaf_3_clk_i),
    .D(_00400_),
    .Q(\in_data[37] ));
 sky130_fd_sc_hd__dfxtp_1 _21988_ (.CLK(clknet_leaf_3_clk_i),
    .D(_00401_),
    .Q(\in_data[38] ));
 sky130_fd_sc_hd__dfxtp_1 _21989_ (.CLK(clknet_leaf_3_clk_i),
    .D(_00402_),
    .Q(\in_data[39] ));
 sky130_fd_sc_hd__dfxtp_1 _21990_ (.CLK(clknet_leaf_3_clk_i),
    .D(_00403_),
    .Q(\in_data[40] ));
 sky130_fd_sc_hd__dfxtp_1 _21991_ (.CLK(clknet_leaf_3_clk_i),
    .D(_00404_),
    .Q(\in_data[41] ));
 sky130_fd_sc_hd__dfxtp_1 _21992_ (.CLK(clknet_leaf_3_clk_i),
    .D(_00405_),
    .Q(\in_data[42] ));
 sky130_fd_sc_hd__dfxtp_1 _21993_ (.CLK(clknet_leaf_3_clk_i),
    .D(_00406_),
    .Q(\in_data[43] ));
 sky130_fd_sc_hd__dfxtp_1 _21994_ (.CLK(clknet_leaf_4_clk_i),
    .D(_00407_),
    .Q(\in_data[44] ));
 sky130_fd_sc_hd__dfxtp_1 _21995_ (.CLK(clknet_leaf_4_clk_i),
    .D(_00408_),
    .Q(\in_data[45] ));
 sky130_fd_sc_hd__dfxtp_1 _21996_ (.CLK(clknet_leaf_4_clk_i),
    .D(_00409_),
    .Q(\in_data[46] ));
 sky130_fd_sc_hd__dfxtp_1 _21997_ (.CLK(clknet_leaf_4_clk_i),
    .D(_00410_),
    .Q(\in_data[47] ));
 sky130_fd_sc_hd__dfxtp_1 _21998_ (.CLK(clknet_leaf_4_clk_i),
    .D(_00411_),
    .Q(\in_data[48] ));
 sky130_fd_sc_hd__dfxtp_1 _21999_ (.CLK(clknet_leaf_9_clk_i),
    .D(_00412_),
    .Q(\in_data[49] ));
 sky130_fd_sc_hd__dfxtp_1 _22000_ (.CLK(clknet_leaf_9_clk_i),
    .D(_00413_),
    .Q(\in_data[50] ));
 sky130_fd_sc_hd__dfxtp_1 _22001_ (.CLK(clknet_leaf_9_clk_i),
    .D(_00414_),
    .Q(\in_data[51] ));
 sky130_fd_sc_hd__dfxtp_1 _22002_ (.CLK(clknet_leaf_9_clk_i),
    .D(_00415_),
    .Q(\in_data[52] ));
 sky130_fd_sc_hd__dfxtp_1 _22003_ (.CLK(clknet_leaf_9_clk_i),
    .D(_00416_),
    .Q(\in_data[53] ));
 sky130_fd_sc_hd__dfxtp_1 _22004_ (.CLK(clknet_leaf_9_clk_i),
    .D(_00417_),
    .Q(\in_data[54] ));
 sky130_fd_sc_hd__dfxtp_1 _22005_ (.CLK(clknet_leaf_9_clk_i),
    .D(_00418_),
    .Q(\in_data[55] ));
 sky130_fd_sc_hd__dfxtp_1 _22006_ (.CLK(clknet_leaf_10_clk_i),
    .D(_00419_),
    .Q(\in_data[56] ));
 sky130_fd_sc_hd__dfxtp_1 _22007_ (.CLK(clknet_leaf_10_clk_i),
    .D(_00420_),
    .Q(\in_data[57] ));
 sky130_fd_sc_hd__dfxtp_1 _22008_ (.CLK(clknet_leaf_10_clk_i),
    .D(_00421_),
    .Q(\in_data[58] ));
 sky130_fd_sc_hd__dfxtp_1 _22009_ (.CLK(clknet_leaf_10_clk_i),
    .D(_00422_),
    .Q(\in_data[59] ));
 sky130_fd_sc_hd__dfxtp_1 _22010_ (.CLK(clknet_leaf_10_clk_i),
    .D(_00423_),
    .Q(\in_data[60] ));
 sky130_fd_sc_hd__dfxtp_1 _22011_ (.CLK(clknet_leaf_10_clk_i),
    .D(_00424_),
    .Q(\in_data[61] ));
 sky130_fd_sc_hd__dfxtp_1 _22012_ (.CLK(clknet_leaf_10_clk_i),
    .D(_00425_),
    .Q(\in_data[62] ));
 sky130_fd_sc_hd__dfxtp_1 _22013_ (.CLK(clknet_leaf_10_clk_i),
    .D(_00426_),
    .Q(\in_data[63] ));
 sky130_fd_sc_hd__dfxtp_1 _22014_ (.CLK(clknet_leaf_2_clk_i),
    .D(_00427_),
    .Q(\in_data[64] ));
 sky130_fd_sc_hd__dfxtp_1 _22015_ (.CLK(clknet_leaf_2_clk_i),
    .D(_00428_),
    .Q(\in_data[65] ));
 sky130_fd_sc_hd__dfxtp_1 _22016_ (.CLK(clknet_leaf_2_clk_i),
    .D(_00429_),
    .Q(\in_data[66] ));
 sky130_fd_sc_hd__dfxtp_1 _22017_ (.CLK(clknet_leaf_3_clk_i),
    .D(_00430_),
    .Q(\in_data[67] ));
 sky130_fd_sc_hd__dfxtp_1 _22018_ (.CLK(clknet_leaf_3_clk_i),
    .D(_00431_),
    .Q(\in_data[68] ));
 sky130_fd_sc_hd__dfxtp_1 _22019_ (.CLK(clknet_leaf_3_clk_i),
    .D(_00432_),
    .Q(\in_data[69] ));
 sky130_fd_sc_hd__dfxtp_1 _22020_ (.CLK(clknet_leaf_3_clk_i),
    .D(_00433_),
    .Q(\in_data[70] ));
 sky130_fd_sc_hd__dfxtp_1 _22021_ (.CLK(clknet_leaf_4_clk_i),
    .D(_00434_),
    .Q(\in_data[71] ));
 sky130_fd_sc_hd__dfxtp_1 _22022_ (.CLK(clknet_leaf_11_clk_i),
    .D(_00435_),
    .Q(\in_data[72] ));
 sky130_fd_sc_hd__dfxtp_1 _22023_ (.CLK(clknet_leaf_11_clk_i),
    .D(_00436_),
    .Q(\in_data[73] ));
 sky130_fd_sc_hd__dfxtp_1 _22024_ (.CLK(clknet_leaf_11_clk_i),
    .D(_00437_),
    .Q(\in_data[74] ));
 sky130_fd_sc_hd__dfxtp_1 _22025_ (.CLK(clknet_leaf_11_clk_i),
    .D(_00438_),
    .Q(\in_data[75] ));
 sky130_fd_sc_hd__dfxtp_1 _22026_ (.CLK(clknet_leaf_11_clk_i),
    .D(_00439_),
    .Q(\in_data[76] ));
 sky130_fd_sc_hd__dfxtp_1 _22027_ (.CLK(clknet_leaf_11_clk_i),
    .D(_00440_),
    .Q(\in_data[77] ));
 sky130_fd_sc_hd__dfxtp_1 _22028_ (.CLK(clknet_leaf_11_clk_i),
    .D(_00441_),
    .Q(\in_data[78] ));
 sky130_fd_sc_hd__dfxtp_1 _22029_ (.CLK(clknet_leaf_11_clk_i),
    .D(_00442_),
    .Q(\in_data[79] ));
 sky130_fd_sc_hd__dfxtp_1 _22030_ (.CLK(clknet_leaf_11_clk_i),
    .D(_00443_),
    .Q(\in_data[80] ));
 sky130_fd_sc_hd__dfxtp_1 _22031_ (.CLK(clknet_leaf_11_clk_i),
    .D(_00444_),
    .Q(\in_data[81] ));
 sky130_fd_sc_hd__dfxtp_1 _22032_ (.CLK(clknet_leaf_11_clk_i),
    .D(_00445_),
    .Q(\in_data[82] ));
 sky130_fd_sc_hd__dfxtp_1 _22033_ (.CLK(clknet_leaf_11_clk_i),
    .D(_00446_),
    .Q(\in_data[83] ));
 sky130_fd_sc_hd__dfxtp_1 _22034_ (.CLK(clknet_leaf_11_clk_i),
    .D(_00447_),
    .Q(\in_data[84] ));
 sky130_fd_sc_hd__dfxtp_1 _22035_ (.CLK(clknet_leaf_11_clk_i),
    .D(_00448_),
    .Q(\in_data[85] ));
 sky130_fd_sc_hd__dfxtp_1 _22036_ (.CLK(clknet_leaf_11_clk_i),
    .D(_00449_),
    .Q(\in_data[86] ));
 sky130_fd_sc_hd__dfxtp_1 _22037_ (.CLK(clknet_leaf_12_clk_i),
    .D(_00450_),
    .Q(\in_data[87] ));
 sky130_fd_sc_hd__dfxtp_1 _22038_ (.CLK(clknet_leaf_11_clk_i),
    .D(_00451_),
    .Q(\in_data[88] ));
 sky130_fd_sc_hd__dfxtp_1 _22039_ (.CLK(clknet_leaf_12_clk_i),
    .D(_00452_),
    .Q(\in_data[89] ));
 sky130_fd_sc_hd__dfxtp_1 _22040_ (.CLK(clknet_leaf_12_clk_i),
    .D(_00453_),
    .Q(\in_data[90] ));
 sky130_fd_sc_hd__dfxtp_1 _22041_ (.CLK(clknet_leaf_12_clk_i),
    .D(_00454_),
    .Q(\in_data[91] ));
 sky130_fd_sc_hd__dfxtp_1 _22042_ (.CLK(clknet_leaf_12_clk_i),
    .D(_00455_),
    .Q(\in_data[92] ));
 sky130_fd_sc_hd__dfxtp_1 _22043_ (.CLK(clknet_leaf_12_clk_i),
    .D(_00456_),
    .Q(\in_data[93] ));
 sky130_fd_sc_hd__dfxtp_1 _22044_ (.CLK(clknet_leaf_12_clk_i),
    .D(_00457_),
    .Q(\in_data[94] ));
 sky130_fd_sc_hd__dfxtp_1 _22045_ (.CLK(clknet_leaf_12_clk_i),
    .D(_00458_),
    .Q(\in_data[95] ));
 sky130_fd_sc_hd__dfxtp_4 _22046_ (.CLK(clknet_leaf_12_clk_i),
    .D(_00459_),
    .Q(\in_data[96] ));
 sky130_fd_sc_hd__dfxtp_4 _22047_ (.CLK(clknet_leaf_12_clk_i),
    .D(_00460_),
    .Q(\in_data[97] ));
 sky130_fd_sc_hd__dfxtp_4 _22048_ (.CLK(clknet_leaf_12_clk_i),
    .D(_00461_),
    .Q(\in_data[98] ));
 sky130_fd_sc_hd__dfxtp_4 _22049_ (.CLK(clknet_leaf_12_clk_i),
    .D(_00462_),
    .Q(\in_data[99] ));
 sky130_fd_sc_hd__dfxtp_4 _22050_ (.CLK(clknet_leaf_13_clk_i),
    .D(_00463_),
    .Q(\in_data[100] ));
 sky130_fd_sc_hd__dfxtp_4 _22051_ (.CLK(clknet_leaf_13_clk_i),
    .D(_00464_),
    .Q(\in_data[101] ));
 sky130_fd_sc_hd__dfxtp_4 _22052_ (.CLK(clknet_leaf_13_clk_i),
    .D(_00465_),
    .Q(\in_data[102] ));
 sky130_fd_sc_hd__dfxtp_4 _22053_ (.CLK(clknet_leaf_13_clk_i),
    .D(_00466_),
    .Q(\in_data[103] ));
 sky130_fd_sc_hd__dfxtp_4 _22054_ (.CLK(clknet_leaf_13_clk_i),
    .D(_00467_),
    .Q(\in_data[104] ));
 sky130_fd_sc_hd__dfxtp_4 _22055_ (.CLK(clknet_leaf_13_clk_i),
    .D(_00468_),
    .Q(\in_data[105] ));
 sky130_fd_sc_hd__dfxtp_4 _22056_ (.CLK(clknet_leaf_13_clk_i),
    .D(_00469_),
    .Q(\in_data[106] ));
 sky130_fd_sc_hd__dfxtp_4 _22057_ (.CLK(clknet_leaf_13_clk_i),
    .D(_00470_),
    .Q(\in_data[107] ));
 sky130_fd_sc_hd__dfxtp_4 _22058_ (.CLK(clknet_leaf_13_clk_i),
    .D(_00471_),
    .Q(\in_data[108] ));
 sky130_fd_sc_hd__dfxtp_4 _22059_ (.CLK(clknet_leaf_13_clk_i),
    .D(_00472_),
    .Q(\in_data[109] ));
 sky130_fd_sc_hd__dfxtp_4 _22060_ (.CLK(clknet_leaf_13_clk_i),
    .D(_00473_),
    .Q(\in_data[110] ));
 sky130_fd_sc_hd__dfxtp_4 _22061_ (.CLK(clknet_leaf_13_clk_i),
    .D(_00474_),
    .Q(\in_data[111] ));
 sky130_fd_sc_hd__dfxtp_4 _22062_ (.CLK(clknet_leaf_13_clk_i),
    .D(_00475_),
    .Q(\in_data[112] ));
 sky130_fd_sc_hd__dfxtp_4 _22063_ (.CLK(clknet_leaf_13_clk_i),
    .D(_00476_),
    .Q(\in_data[113] ));
 sky130_fd_sc_hd__dfrtp_4 _22064_ (.CLK(clknet_leaf_35_clk_i),
    .D(_00477_),
    .RESET_B(net639),
    .Q(mstream_o[0]));
 sky130_fd_sc_hd__dfrtp_4 _22065_ (.CLK(clknet_leaf_35_clk_i),
    .D(_00478_),
    .RESET_B(net639),
    .Q(mstream_o[1]));
 sky130_fd_sc_hd__dfrtp_4 _22066_ (.CLK(clknet_leaf_35_clk_i),
    .D(_00479_),
    .RESET_B(net639),
    .Q(mstream_o[2]));
 sky130_fd_sc_hd__dfrtp_4 _22067_ (.CLK(clknet_leaf_35_clk_i),
    .D(_00480_),
    .RESET_B(net639),
    .Q(mstream_o[3]));
 sky130_fd_sc_hd__dfrtp_4 _22068_ (.CLK(clknet_leaf_35_clk_i),
    .D(_00481_),
    .RESET_B(net639),
    .Q(mstream_o[4]));
 sky130_fd_sc_hd__dfrtp_4 _22069_ (.CLK(clknet_leaf_35_clk_i),
    .D(_00482_),
    .RESET_B(net639),
    .Q(mstream_o[5]));
 sky130_fd_sc_hd__dfrtp_4 _22070_ (.CLK(clknet_leaf_34_clk_i),
    .D(_00483_),
    .RESET_B(net639),
    .Q(mstream_o[6]));
 sky130_fd_sc_hd__dfrtp_4 _22071_ (.CLK(clknet_leaf_34_clk_i),
    .D(_00484_),
    .RESET_B(net639),
    .Q(mstream_o[7]));
 sky130_fd_sc_hd__dfrtp_4 _22072_ (.CLK(clknet_leaf_34_clk_i),
    .D(_00485_),
    .RESET_B(net639),
    .Q(mstream_o[8]));
 sky130_fd_sc_hd__dfrtp_4 _22073_ (.CLK(clknet_leaf_34_clk_i),
    .D(_00486_),
    .RESET_B(net639),
    .Q(mstream_o[9]));
 sky130_fd_sc_hd__dfrtp_4 _22074_ (.CLK(clknet_leaf_34_clk_i),
    .D(_00487_),
    .RESET_B(net639),
    .Q(mstream_o[10]));
 sky130_fd_sc_hd__dfrtp_4 _22075_ (.CLK(clknet_leaf_34_clk_i),
    .D(_00488_),
    .RESET_B(net636),
    .Q(mstream_o[11]));
 sky130_fd_sc_hd__dfrtp_4 _22076_ (.CLK(clknet_leaf_34_clk_i),
    .D(_00489_),
    .RESET_B(net636),
    .Q(mstream_o[12]));
 sky130_fd_sc_hd__dfrtp_4 _22077_ (.CLK(clknet_leaf_34_clk_i),
    .D(_00490_),
    .RESET_B(net636),
    .Q(mstream_o[13]));
 sky130_fd_sc_hd__dfrtp_4 _22078_ (.CLK(clknet_leaf_34_clk_i),
    .D(_00491_),
    .RESET_B(net636),
    .Q(mstream_o[14]));
 sky130_fd_sc_hd__dfrtp_4 _22079_ (.CLK(clknet_leaf_33_clk_i),
    .D(_00492_),
    .RESET_B(net636),
    .Q(mstream_o[15]));
 sky130_fd_sc_hd__dfrtp_4 _22080_ (.CLK(clknet_leaf_34_clk_i),
    .D(_00493_),
    .RESET_B(net636),
    .Q(mstream_o[16]));
 sky130_fd_sc_hd__dfrtp_4 _22081_ (.CLK(clknet_leaf_33_clk_i),
    .D(_00494_),
    .RESET_B(net636),
    .Q(mstream_o[17]));
 sky130_fd_sc_hd__dfrtp_4 _22082_ (.CLK(clknet_leaf_33_clk_i),
    .D(_00495_),
    .RESET_B(net636),
    .Q(mstream_o[18]));
 sky130_fd_sc_hd__dfrtp_4 _22083_ (.CLK(clknet_leaf_33_clk_i),
    .D(_00496_),
    .RESET_B(net636),
    .Q(mstream_o[19]));
 sky130_fd_sc_hd__dfrtp_4 _22084_ (.CLK(clknet_leaf_33_clk_i),
    .D(_00497_),
    .RESET_B(net636),
    .Q(mstream_o[20]));
 sky130_fd_sc_hd__dfrtp_4 _22085_ (.CLK(clknet_leaf_33_clk_i),
    .D(_00498_),
    .RESET_B(net636),
    .Q(mstream_o[21]));
 sky130_fd_sc_hd__dfrtp_4 _22086_ (.CLK(clknet_leaf_33_clk_i),
    .D(_00499_),
    .RESET_B(net636),
    .Q(mstream_o[22]));
 sky130_fd_sc_hd__dfrtp_4 _22087_ (.CLK(clknet_leaf_33_clk_i),
    .D(_00500_),
    .RESET_B(net636),
    .Q(mstream_o[23]));
 sky130_fd_sc_hd__dfrtp_4 _22088_ (.CLK(clknet_leaf_33_clk_i),
    .D(_00501_),
    .RESET_B(net636),
    .Q(mstream_o[24]));
 sky130_fd_sc_hd__dfrtp_4 _22089_ (.CLK(clknet_leaf_33_clk_i),
    .D(_00502_),
    .RESET_B(net636),
    .Q(mstream_o[25]));
 sky130_fd_sc_hd__dfrtp_4 _22090_ (.CLK(clknet_leaf_32_clk_i),
    .D(_00503_),
    .RESET_B(net637),
    .Q(mstream_o[26]));
 sky130_fd_sc_hd__dfrtp_4 _22091_ (.CLK(clknet_leaf_32_clk_i),
    .D(_00504_),
    .RESET_B(net637),
    .Q(mstream_o[27]));
 sky130_fd_sc_hd__dfrtp_4 _22092_ (.CLK(clknet_leaf_33_clk_i),
    .D(_00505_),
    .RESET_B(net638),
    .Q(mstream_o[28]));
 sky130_fd_sc_hd__dfrtp_4 _22093_ (.CLK(clknet_leaf_32_clk_i),
    .D(_00506_),
    .RESET_B(net637),
    .Q(mstream_o[29]));
 sky130_fd_sc_hd__dfrtp_4 _22094_ (.CLK(clknet_leaf_32_clk_i),
    .D(_00507_),
    .RESET_B(net637),
    .Q(mstream_o[30]));
 sky130_fd_sc_hd__dfrtp_4 _22095_ (.CLK(clknet_leaf_32_clk_i),
    .D(_00508_),
    .RESET_B(net637),
    .Q(mstream_o[31]));
 sky130_fd_sc_hd__dfrtp_4 _22096_ (.CLK(clknet_leaf_33_clk_i),
    .D(_00509_),
    .RESET_B(net636),
    .Q(mstream_o[32]));
 sky130_fd_sc_hd__dfrtp_4 _22097_ (.CLK(clknet_leaf_32_clk_i),
    .D(_00510_),
    .RESET_B(net637),
    .Q(mstream_o[33]));
 sky130_fd_sc_hd__dfrtp_4 _22098_ (.CLK(clknet_leaf_32_clk_i),
    .D(_00511_),
    .RESET_B(net637),
    .Q(mstream_o[34]));
 sky130_fd_sc_hd__dfrtp_4 _22099_ (.CLK(clknet_leaf_32_clk_i),
    .D(_00512_),
    .RESET_B(net637),
    .Q(mstream_o[35]));
 sky130_fd_sc_hd__dfrtp_4 _22100_ (.CLK(clknet_leaf_32_clk_i),
    .D(_00513_),
    .RESET_B(net637),
    .Q(mstream_o[36]));
 sky130_fd_sc_hd__dfrtp_4 _22101_ (.CLK(clknet_leaf_32_clk_i),
    .D(_00514_),
    .RESET_B(net637),
    .Q(mstream_o[37]));
 sky130_fd_sc_hd__dfrtp_4 _22102_ (.CLK(clknet_leaf_32_clk_i),
    .D(_00515_),
    .RESET_B(net638),
    .Q(mstream_o[38]));
 sky130_fd_sc_hd__dfrtp_4 _22103_ (.CLK(clknet_leaf_32_clk_i),
    .D(_00516_),
    .RESET_B(net637),
    .Q(mstream_o[39]));
 sky130_fd_sc_hd__dfrtp_4 _22104_ (.CLK(clknet_leaf_32_clk_i),
    .D(_00517_),
    .RESET_B(net637),
    .Q(mstream_o[40]));
 sky130_fd_sc_hd__dfrtp_4 _22105_ (.CLK(clknet_leaf_32_clk_i),
    .D(_00518_),
    .RESET_B(net638),
    .Q(mstream_o[41]));
 sky130_fd_sc_hd__dfrtp_4 _22106_ (.CLK(clknet_leaf_31_clk_i),
    .D(_00519_),
    .RESET_B(net638),
    .Q(mstream_o[42]));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk_i (.A(clk_i),
    .X(clknet_0_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_0__f_clk_i (.A(clknet_0_clk_i),
    .X(clknet_2_0__leaf_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_1__f_clk_i (.A(clknet_0_clk_i),
    .X(clknet_2_1__leaf_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_2__f_clk_i (.A(clknet_0_clk_i),
    .X(clknet_2_2__leaf_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_3__f_clk_i (.A(clknet_0_clk_i),
    .X(clknet_2_3__leaf_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_0_clk_i (.A(clknet_2_0__leaf_clk_i),
    .X(clknet_leaf_0_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_10_clk_i (.A(clknet_2_1__leaf_clk_i),
    .X(clknet_leaf_10_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_11_clk_i (.A(clknet_2_1__leaf_clk_i),
    .X(clknet_leaf_11_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_12_clk_i (.A(clknet_2_1__leaf_clk_i),
    .X(clknet_leaf_12_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_13_clk_i (.A(clknet_2_1__leaf_clk_i),
    .X(clknet_leaf_13_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_14_clk_i (.A(clknet_2_1__leaf_clk_i),
    .X(clknet_leaf_14_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_15_clk_i (.A(clknet_2_1__leaf_clk_i),
    .X(clknet_leaf_15_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_16_clk_i (.A(clknet_2_3__leaf_clk_i),
    .X(clknet_leaf_16_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_17_clk_i (.A(clknet_2_3__leaf_clk_i),
    .X(clknet_leaf_17_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_18_clk_i (.A(clknet_2_3__leaf_clk_i),
    .X(clknet_leaf_18_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_19_clk_i (.A(clknet_2_3__leaf_clk_i),
    .X(clknet_leaf_19_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_1_clk_i (.A(clknet_2_0__leaf_clk_i),
    .X(clknet_leaf_1_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_20_clk_i (.A(clknet_2_3__leaf_clk_i),
    .X(clknet_leaf_20_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_21_clk_i (.A(clknet_2_3__leaf_clk_i),
    .X(clknet_leaf_21_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_22_clk_i (.A(clknet_2_3__leaf_clk_i),
    .X(clknet_leaf_22_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_23_clk_i (.A(clknet_2_3__leaf_clk_i),
    .X(clknet_leaf_23_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_24_clk_i (.A(clknet_2_3__leaf_clk_i),
    .X(clknet_leaf_24_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_25_clk_i (.A(clknet_2_3__leaf_clk_i),
    .X(clknet_leaf_25_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_26_clk_i (.A(clknet_2_3__leaf_clk_i),
    .X(clknet_leaf_26_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_27_clk_i (.A(clknet_2_3__leaf_clk_i),
    .X(clknet_leaf_27_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_28_clk_i (.A(clknet_2_2__leaf_clk_i),
    .X(clknet_leaf_28_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_29_clk_i (.A(clknet_2_2__leaf_clk_i),
    .X(clknet_leaf_29_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_2_clk_i (.A(clknet_2_0__leaf_clk_i),
    .X(clknet_leaf_2_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_30_clk_i (.A(clknet_2_3__leaf_clk_i),
    .X(clknet_leaf_30_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_31_clk_i (.A(clknet_2_2__leaf_clk_i),
    .X(clknet_leaf_31_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_32_clk_i (.A(clknet_2_2__leaf_clk_i),
    .X(clknet_leaf_32_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_33_clk_i (.A(clknet_2_2__leaf_clk_i),
    .X(clknet_leaf_33_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_34_clk_i (.A(clknet_2_2__leaf_clk_i),
    .X(clknet_leaf_34_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_35_clk_i (.A(clknet_2_2__leaf_clk_i),
    .X(clknet_leaf_35_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_36_clk_i (.A(clknet_2_2__leaf_clk_i),
    .X(clknet_leaf_36_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_37_clk_i (.A(clknet_2_2__leaf_clk_i),
    .X(clknet_leaf_37_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_38_clk_i (.A(clknet_2_2__leaf_clk_i),
    .X(clknet_leaf_38_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_3_clk_i (.A(clknet_2_0__leaf_clk_i),
    .X(clknet_leaf_3_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_40_clk_i (.A(clknet_2_0__leaf_clk_i),
    .X(clknet_leaf_40_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_41_clk_i (.A(clknet_2_0__leaf_clk_i),
    .X(clknet_leaf_41_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_43_clk_i (.A(clknet_2_0__leaf_clk_i),
    .X(clknet_leaf_43_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_44_clk_i (.A(clknet_2_0__leaf_clk_i),
    .X(clknet_leaf_44_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_4_clk_i (.A(clknet_2_1__leaf_clk_i),
    .X(clknet_leaf_4_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_5_clk_i (.A(clknet_2_1__leaf_clk_i),
    .X(clknet_leaf_5_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_6_clk_i (.A(clknet_2_1__leaf_clk_i),
    .X(clknet_leaf_6_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_7_clk_i (.A(clknet_2_1__leaf_clk_i),
    .X(clknet_leaf_7_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_9_clk_i (.A(clknet_2_1__leaf_clk_i),
    .X(clknet_leaf_9_clk_i));
 sky130_fd_sc_hd__clkbuf_8 fanout1 (.A(net2),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_8 fanout10 (.A(_03050_),
    .X(net10));
 sky130_fd_sc_hd__buf_4 fanout100 (.A(net101),
    .X(net100));
 sky130_fd_sc_hd__clkbuf_8 fanout101 (.A(\mul1.b[20] ),
    .X(net101));
 sky130_fd_sc_hd__buf_6 fanout102 (.A(\mul1.b[19] ),
    .X(net102));
 sky130_fd_sc_hd__buf_4 fanout103 (.A(net106),
    .X(net103));
 sky130_fd_sc_hd__buf_2 fanout104 (.A(net106),
    .X(net104));
 sky130_fd_sc_hd__buf_4 fanout105 (.A(net106),
    .X(net105));
 sky130_fd_sc_hd__clkbuf_4 fanout106 (.A(\mul1.b[19] ),
    .X(net106));
 sky130_fd_sc_hd__clkbuf_8 fanout107 (.A(net112),
    .X(net107));
 sky130_fd_sc_hd__buf_4 fanout108 (.A(net111),
    .X(net108));
 sky130_fd_sc_hd__buf_2 fanout109 (.A(net111),
    .X(net109));
 sky130_fd_sc_hd__clkbuf_8 fanout11 (.A(net13),
    .X(net11));
 sky130_fd_sc_hd__buf_4 fanout110 (.A(net111),
    .X(net110));
 sky130_fd_sc_hd__clkbuf_4 fanout111 (.A(net112),
    .X(net111));
 sky130_fd_sc_hd__buf_4 fanout112 (.A(\mul1.b[18] ),
    .X(net112));
 sky130_fd_sc_hd__buf_4 fanout113 (.A(net114),
    .X(net113));
 sky130_fd_sc_hd__clkbuf_8 fanout114 (.A(\mul1.b[17] ),
    .X(net114));
 sky130_fd_sc_hd__buf_4 fanout115 (.A(net116),
    .X(net115));
 sky130_fd_sc_hd__buf_6 fanout116 (.A(\mul1.b[17] ),
    .X(net116));
 sky130_fd_sc_hd__buf_4 fanout117 (.A(net118),
    .X(net117));
 sky130_fd_sc_hd__clkbuf_8 fanout118 (.A(net121),
    .X(net118));
 sky130_fd_sc_hd__buf_4 fanout119 (.A(net120),
    .X(net119));
 sky130_fd_sc_hd__buf_6 fanout12 (.A(net13),
    .X(net12));
 sky130_fd_sc_hd__buf_6 fanout120 (.A(net121),
    .X(net120));
 sky130_fd_sc_hd__buf_4 fanout121 (.A(\mul1.b[16] ),
    .X(net121));
 sky130_fd_sc_hd__buf_4 fanout122 (.A(net123),
    .X(net122));
 sky130_fd_sc_hd__clkbuf_8 fanout123 (.A(net126),
    .X(net123));
 sky130_fd_sc_hd__buf_4 fanout124 (.A(net125),
    .X(net124));
 sky130_fd_sc_hd__buf_8 fanout125 (.A(net126),
    .X(net125));
 sky130_fd_sc_hd__buf_4 fanout126 (.A(\mul1.b[15] ),
    .X(net126));
 sky130_fd_sc_hd__clkbuf_8 fanout127 (.A(net128),
    .X(net127));
 sky130_fd_sc_hd__clkbuf_8 fanout128 (.A(\mul1.b[14] ),
    .X(net128));
 sky130_fd_sc_hd__clkbuf_8 fanout129 (.A(net130),
    .X(net129));
 sky130_fd_sc_hd__buf_6 fanout13 (.A(_02920_),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_8 fanout130 (.A(\mul1.b[14] ),
    .X(net130));
 sky130_fd_sc_hd__buf_4 fanout131 (.A(net132),
    .X(net131));
 sky130_fd_sc_hd__buf_4 fanout132 (.A(net135),
    .X(net132));
 sky130_fd_sc_hd__clkbuf_8 fanout133 (.A(net135),
    .X(net133));
 sky130_fd_sc_hd__buf_4 fanout134 (.A(net135),
    .X(net134));
 sky130_fd_sc_hd__buf_4 fanout135 (.A(\mul1.b[13] ),
    .X(net135));
 sky130_fd_sc_hd__buf_4 fanout136 (.A(net137),
    .X(net136));
 sky130_fd_sc_hd__clkbuf_8 fanout137 (.A(\mul1.b[12] ),
    .X(net137));
 sky130_fd_sc_hd__clkbuf_8 fanout138 (.A(net140),
    .X(net138));
 sky130_fd_sc_hd__buf_4 fanout139 (.A(net140),
    .X(net139));
 sky130_fd_sc_hd__clkbuf_8 fanout14 (.A(net16),
    .X(net14));
 sky130_fd_sc_hd__buf_4 fanout140 (.A(\mul1.b[12] ),
    .X(net140));
 sky130_fd_sc_hd__buf_4 fanout141 (.A(net142),
    .X(net141));
 sky130_fd_sc_hd__clkbuf_4 fanout142 (.A(\mul1.b[11] ),
    .X(net142));
 sky130_fd_sc_hd__clkbuf_8 fanout143 (.A(net144),
    .X(net143));
 sky130_fd_sc_hd__clkbuf_8 fanout144 (.A(\mul1.b[11] ),
    .X(net144));
 sky130_fd_sc_hd__buf_4 fanout145 (.A(net146),
    .X(net145));
 sky130_fd_sc_hd__buf_2 fanout146 (.A(\mul1.b[10] ),
    .X(net146));
 sky130_fd_sc_hd__clkbuf_8 fanout147 (.A(net149),
    .X(net147));
 sky130_fd_sc_hd__buf_6 fanout148 (.A(net149),
    .X(net148));
 sky130_fd_sc_hd__clkbuf_4 fanout149 (.A(\mul1.b[10] ),
    .X(net149));
 sky130_fd_sc_hd__clkbuf_4 fanout15 (.A(net16),
    .X(net15));
 sky130_fd_sc_hd__buf_4 fanout150 (.A(net151),
    .X(net150));
 sky130_fd_sc_hd__buf_2 fanout151 (.A(\mul1.b[9] ),
    .X(net151));
 sky130_fd_sc_hd__buf_4 fanout152 (.A(net154),
    .X(net152));
 sky130_fd_sc_hd__buf_6 fanout153 (.A(net154),
    .X(net153));
 sky130_fd_sc_hd__buf_4 fanout154 (.A(\mul1.b[9] ),
    .X(net154));
 sky130_fd_sc_hd__clkbuf_8 fanout155 (.A(\mul1.b[8] ),
    .X(net155));
 sky130_fd_sc_hd__clkbuf_8 fanout156 (.A(net158),
    .X(net156));
 sky130_fd_sc_hd__clkbuf_8 fanout157 (.A(net158),
    .X(net157));
 sky130_fd_sc_hd__buf_6 fanout158 (.A(\mul1.b[8] ),
    .X(net158));
 sky130_fd_sc_hd__buf_4 fanout159 (.A(net160),
    .X(net159));
 sky130_fd_sc_hd__clkbuf_4 fanout160 (.A(\mul1.b[7] ),
    .X(net160));
 sky130_fd_sc_hd__clkbuf_8 fanout161 (.A(net164),
    .X(net161));
 sky130_fd_sc_hd__clkbuf_8 fanout162 (.A(net164),
    .X(net162));
 sky130_fd_sc_hd__clkbuf_4 fanout163 (.A(net164),
    .X(net163));
 sky130_fd_sc_hd__clkbuf_4 fanout164 (.A(\mul1.b[7] ),
    .X(net164));
 sky130_fd_sc_hd__buf_4 fanout165 (.A(net166),
    .X(net165));
 sky130_fd_sc_hd__clkbuf_4 fanout166 (.A(\mul1.b[6] ),
    .X(net166));
 sky130_fd_sc_hd__clkbuf_8 fanout167 (.A(net170),
    .X(net167));
 sky130_fd_sc_hd__clkbuf_4 fanout168 (.A(net170),
    .X(net168));
 sky130_fd_sc_hd__buf_4 fanout169 (.A(net170),
    .X(net169));
 sky130_fd_sc_hd__buf_4 fanout17 (.A(net19),
    .X(net17));
 sky130_fd_sc_hd__buf_4 fanout170 (.A(\mul1.b[6] ),
    .X(net170));
 sky130_fd_sc_hd__buf_4 fanout171 (.A(net172),
    .X(net171));
 sky130_fd_sc_hd__buf_2 fanout172 (.A(\mul1.b[5] ),
    .X(net172));
 sky130_fd_sc_hd__buf_4 fanout173 (.A(net174),
    .X(net173));
 sky130_fd_sc_hd__buf_4 fanout174 (.A(net175),
    .X(net174));
 sky130_fd_sc_hd__clkbuf_4 fanout175 (.A(\mul1.b[5] ),
    .X(net175));
 sky130_fd_sc_hd__buf_4 fanout176 (.A(net177),
    .X(net176));
 sky130_fd_sc_hd__clkbuf_4 fanout177 (.A(\mul1.b[4] ),
    .X(net177));
 sky130_fd_sc_hd__buf_4 fanout178 (.A(net180),
    .X(net178));
 sky130_fd_sc_hd__buf_4 fanout179 (.A(net180),
    .X(net179));
 sky130_fd_sc_hd__clkbuf_4 fanout18 (.A(net19),
    .X(net18));
 sky130_fd_sc_hd__buf_4 fanout180 (.A(\mul1.b[4] ),
    .X(net180));
 sky130_fd_sc_hd__buf_4 fanout181 (.A(net182),
    .X(net181));
 sky130_fd_sc_hd__clkbuf_2 fanout182 (.A(\mul1.b[3] ),
    .X(net182));
 sky130_fd_sc_hd__buf_4 fanout183 (.A(net185),
    .X(net183));
 sky130_fd_sc_hd__buf_4 fanout184 (.A(net185),
    .X(net184));
 sky130_fd_sc_hd__buf_4 fanout185 (.A(\mul1.b[3] ),
    .X(net185));
 sky130_fd_sc_hd__buf_4 fanout186 (.A(\mul1.b[2] ),
    .X(net186));
 sky130_fd_sc_hd__buf_4 fanout187 (.A(\mul1.b[2] ),
    .X(net187));
 sky130_fd_sc_hd__buf_4 fanout188 (.A(net189),
    .X(net188));
 sky130_fd_sc_hd__buf_4 fanout189 (.A(\mul1.b[1] ),
    .X(net189));
 sky130_fd_sc_hd__buf_4 fanout19 (.A(_02823_),
    .X(net19));
 sky130_fd_sc_hd__buf_4 fanout190 (.A(net191),
    .X(net190));
 sky130_fd_sc_hd__clkbuf_4 fanout191 (.A(net192),
    .X(net191));
 sky130_fd_sc_hd__clkbuf_4 fanout192 (.A(\mul1.b[1] ),
    .X(net192));
 sky130_fd_sc_hd__buf_4 fanout193 (.A(net194),
    .X(net193));
 sky130_fd_sc_hd__buf_4 fanout194 (.A(net973),
    .X(net194));
 sky130_fd_sc_hd__buf_4 fanout195 (.A(net196),
    .X(net195));
 sky130_fd_sc_hd__buf_4 fanout196 (.A(\mul1.a[30] ),
    .X(net196));
 sky130_fd_sc_hd__buf_4 fanout197 (.A(net198),
    .X(net197));
 sky130_fd_sc_hd__clkbuf_8 fanout198 (.A(\mul1.a[29] ),
    .X(net198));
 sky130_fd_sc_hd__buf_4 fanout199 (.A(net201),
    .X(net199));
 sky130_fd_sc_hd__buf_4 fanout2 (.A(_03055_),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_8 fanout20 (.A(_02823_),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_4 fanout200 (.A(net201),
    .X(net200));
 sky130_fd_sc_hd__clkbuf_8 fanout201 (.A(\mul1.a[28] ),
    .X(net201));
 sky130_fd_sc_hd__clkbuf_8 fanout202 (.A(\mul1.a[27] ),
    .X(net202));
 sky130_fd_sc_hd__buf_4 fanout203 (.A(\mul1.a[27] ),
    .X(net203));
 sky130_fd_sc_hd__buf_4 fanout204 (.A(\mul1.a[27] ),
    .X(net204));
 sky130_fd_sc_hd__clkbuf_8 fanout205 (.A(net206),
    .X(net205));
 sky130_fd_sc_hd__buf_4 fanout206 (.A(\mul1.a[26] ),
    .X(net206));
 sky130_fd_sc_hd__buf_4 fanout207 (.A(\mul1.a[26] ),
    .X(net207));
 sky130_fd_sc_hd__clkbuf_8 fanout208 (.A(net209),
    .X(net208));
 sky130_fd_sc_hd__buf_4 fanout209 (.A(\mul1.a[25] ),
    .X(net209));
 sky130_fd_sc_hd__clkbuf_4 fanout21 (.A(_02823_),
    .X(net21));
 sky130_fd_sc_hd__buf_4 fanout210 (.A(\mul1.a[25] ),
    .X(net210));
 sky130_fd_sc_hd__clkbuf_8 fanout211 (.A(net212),
    .X(net211));
 sky130_fd_sc_hd__buf_4 fanout212 (.A(net214),
    .X(net212));
 sky130_fd_sc_hd__buf_4 fanout213 (.A(net214),
    .X(net213));
 sky130_fd_sc_hd__clkbuf_4 fanout214 (.A(net978),
    .X(net214));
 sky130_fd_sc_hd__clkbuf_8 fanout215 (.A(net216),
    .X(net215));
 sky130_fd_sc_hd__buf_4 fanout216 (.A(net218),
    .X(net216));
 sky130_fd_sc_hd__buf_4 fanout217 (.A(net218),
    .X(net217));
 sky130_fd_sc_hd__buf_4 fanout218 (.A(net969),
    .X(net218));
 sky130_fd_sc_hd__buf_4 fanout219 (.A(net221),
    .X(net219));
 sky130_fd_sc_hd__buf_4 fanout22 (.A(net23),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_4 fanout220 (.A(net221),
    .X(net220));
 sky130_fd_sc_hd__buf_2 fanout221 (.A(net223),
    .X(net221));
 sky130_fd_sc_hd__buf_4 fanout222 (.A(net223),
    .X(net222));
 sky130_fd_sc_hd__clkbuf_4 fanout223 (.A(net974),
    .X(net223));
 sky130_fd_sc_hd__buf_4 fanout224 (.A(net225),
    .X(net224));
 sky130_fd_sc_hd__buf_4 fanout225 (.A(net227),
    .X(net225));
 sky130_fd_sc_hd__buf_4 fanout226 (.A(net227),
    .X(net226));
 sky130_fd_sc_hd__clkbuf_8 fanout227 (.A(net970),
    .X(net227));
 sky130_fd_sc_hd__buf_4 fanout228 (.A(net229),
    .X(net228));
 sky130_fd_sc_hd__clkbuf_4 fanout229 (.A(net231),
    .X(net229));
 sky130_fd_sc_hd__buf_4 fanout23 (.A(_02757_),
    .X(net23));
 sky130_fd_sc_hd__buf_4 fanout230 (.A(net231),
    .X(net230));
 sky130_fd_sc_hd__clkbuf_4 fanout231 (.A(net232),
    .X(net231));
 sky130_fd_sc_hd__buf_4 fanout232 (.A(net977),
    .X(net232));
 sky130_fd_sc_hd__buf_4 fanout233 (.A(net235),
    .X(net233));
 sky130_fd_sc_hd__buf_2 fanout234 (.A(net235),
    .X(net234));
 sky130_fd_sc_hd__buf_4 fanout235 (.A(\mul1.a[19] ),
    .X(net235));
 sky130_fd_sc_hd__buf_4 fanout236 (.A(net237),
    .X(net236));
 sky130_fd_sc_hd__buf_2 fanout237 (.A(\mul1.a[19] ),
    .X(net237));
 sky130_fd_sc_hd__buf_4 fanout238 (.A(net240),
    .X(net238));
 sky130_fd_sc_hd__clkbuf_4 fanout239 (.A(net240),
    .X(net239));
 sky130_fd_sc_hd__clkbuf_8 fanout24 (.A(net25),
    .X(net24));
 sky130_fd_sc_hd__buf_4 fanout240 (.A(\mul1.a[18] ),
    .X(net240));
 sky130_fd_sc_hd__buf_4 fanout241 (.A(net242),
    .X(net241));
 sky130_fd_sc_hd__clkbuf_4 fanout242 (.A(\mul1.a[18] ),
    .X(net242));
 sky130_fd_sc_hd__buf_4 fanout243 (.A(net244),
    .X(net243));
 sky130_fd_sc_hd__clkbuf_4 fanout244 (.A(\mul1.a[17] ),
    .X(net244));
 sky130_fd_sc_hd__buf_4 fanout245 (.A(net246),
    .X(net245));
 sky130_fd_sc_hd__buf_2 fanout246 (.A(\mul1.a[17] ),
    .X(net246));
 sky130_fd_sc_hd__buf_4 fanout247 (.A(\mul1.a[17] ),
    .X(net247));
 sky130_fd_sc_hd__buf_4 fanout248 (.A(net249),
    .X(net248));
 sky130_fd_sc_hd__clkbuf_4 fanout249 (.A(net251),
    .X(net249));
 sky130_fd_sc_hd__buf_6 fanout25 (.A(net26),
    .X(net25));
 sky130_fd_sc_hd__buf_4 fanout250 (.A(net251),
    .X(net250));
 sky130_fd_sc_hd__buf_6 fanout251 (.A(net252),
    .X(net251));
 sky130_fd_sc_hd__buf_4 fanout252 (.A(net976),
    .X(net252));
 sky130_fd_sc_hd__buf_4 fanout253 (.A(net257),
    .X(net253));
 sky130_fd_sc_hd__clkbuf_2 fanout254 (.A(net257),
    .X(net254));
 sky130_fd_sc_hd__buf_4 fanout255 (.A(net256),
    .X(net255));
 sky130_fd_sc_hd__clkbuf_8 fanout256 (.A(net257),
    .X(net256));
 sky130_fd_sc_hd__buf_8 fanout257 (.A(net968),
    .X(net257));
 sky130_fd_sc_hd__clkbuf_8 fanout258 (.A(\mul1.a[13] ),
    .X(net258));
 sky130_fd_sc_hd__buf_4 fanout259 (.A(net260),
    .X(net259));
 sky130_fd_sc_hd__buf_8 fanout26 (.A(_02756_),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_4 fanout260 (.A(net262),
    .X(net260));
 sky130_fd_sc_hd__buf_4 fanout261 (.A(net262),
    .X(net261));
 sky130_fd_sc_hd__buf_4 fanout262 (.A(\mul1.a[13] ),
    .X(net262));
 sky130_fd_sc_hd__clkbuf_8 fanout263 (.A(\mul1.a[12] ),
    .X(net263));
 sky130_fd_sc_hd__buf_4 fanout264 (.A(net266),
    .X(net264));
 sky130_fd_sc_hd__buf_4 fanout265 (.A(net266),
    .X(net265));
 sky130_fd_sc_hd__clkbuf_4 fanout266 (.A(net267),
    .X(net266));
 sky130_fd_sc_hd__clkbuf_4 fanout267 (.A(\mul1.a[12] ),
    .X(net267));
 sky130_fd_sc_hd__clkbuf_8 fanout268 (.A(net272),
    .X(net268));
 sky130_fd_sc_hd__buf_4 fanout269 (.A(net270),
    .X(net269));
 sky130_fd_sc_hd__buf_6 fanout27 (.A(_02756_),
    .X(net27));
 sky130_fd_sc_hd__buf_4 fanout270 (.A(net271),
    .X(net270));
 sky130_fd_sc_hd__buf_4 fanout271 (.A(net272),
    .X(net271));
 sky130_fd_sc_hd__buf_4 fanout272 (.A(\mul1.a[11] ),
    .X(net272));
 sky130_fd_sc_hd__clkbuf_8 fanout273 (.A(\mul1.a[10] ),
    .X(net273));
 sky130_fd_sc_hd__buf_2 fanout274 (.A(\mul1.a[10] ),
    .X(net274));
 sky130_fd_sc_hd__clkbuf_8 fanout275 (.A(net276),
    .X(net275));
 sky130_fd_sc_hd__buf_4 fanout276 (.A(net277),
    .X(net276));
 sky130_fd_sc_hd__buf_4 fanout277 (.A(\mul1.a[10] ),
    .X(net277));
 sky130_fd_sc_hd__clkbuf_8 fanout278 (.A(\mul1.a[9] ),
    .X(net278));
 sky130_fd_sc_hd__clkbuf_4 fanout279 (.A(\mul1.a[9] ),
    .X(net279));
 sky130_fd_sc_hd__buf_4 fanout28 (.A(net29),
    .X(net28));
 sky130_fd_sc_hd__clkbuf_8 fanout280 (.A(net281),
    .X(net280));
 sky130_fd_sc_hd__buf_4 fanout281 (.A(net282),
    .X(net281));
 sky130_fd_sc_hd__buf_4 fanout282 (.A(\mul1.a[9] ),
    .X(net282));
 sky130_fd_sc_hd__buf_4 fanout283 (.A(net284),
    .X(net283));
 sky130_fd_sc_hd__clkbuf_8 fanout284 (.A(\mul1.a[8] ),
    .X(net284));
 sky130_fd_sc_hd__buf_4 fanout285 (.A(net286),
    .X(net285));
 sky130_fd_sc_hd__buf_4 fanout286 (.A(net287),
    .X(net286));
 sky130_fd_sc_hd__buf_4 fanout287 (.A(\mul1.a[8] ),
    .X(net287));
 sky130_fd_sc_hd__buf_4 fanout288 (.A(net289),
    .X(net288));
 sky130_fd_sc_hd__buf_6 fanout289 (.A(net292),
    .X(net289));
 sky130_fd_sc_hd__clkbuf_8 fanout29 (.A(_02755_),
    .X(net29));
 sky130_fd_sc_hd__clkbuf_8 fanout290 (.A(net292),
    .X(net290));
 sky130_fd_sc_hd__clkbuf_4 fanout291 (.A(net292),
    .X(net291));
 sky130_fd_sc_hd__buf_8 fanout292 (.A(\mul1.a[7] ),
    .X(net292));
 sky130_fd_sc_hd__clkbuf_8 fanout293 (.A(net294),
    .X(net293));
 sky130_fd_sc_hd__clkbuf_4 fanout294 (.A(net295),
    .X(net294));
 sky130_fd_sc_hd__clkbuf_8 fanout295 (.A(\mul1.a[6] ),
    .X(net295));
 sky130_fd_sc_hd__clkbuf_8 fanout296 (.A(\mul1.a[6] ),
    .X(net296));
 sky130_fd_sc_hd__clkbuf_4 fanout297 (.A(\mul1.a[6] ),
    .X(net297));
 sky130_fd_sc_hd__clkbuf_8 fanout298 (.A(net299),
    .X(net298));
 sky130_fd_sc_hd__clkbuf_4 fanout299 (.A(net300),
    .X(net299));
 sky130_fd_sc_hd__clkbuf_8 fanout3 (.A(_03055_),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_8 fanout30 (.A(net31),
    .X(net30));
 sky130_fd_sc_hd__buf_4 fanout300 (.A(\mul1.a[5] ),
    .X(net300));
 sky130_fd_sc_hd__clkbuf_8 fanout301 (.A(\mul1.a[5] ),
    .X(net301));
 sky130_fd_sc_hd__buf_2 fanout302 (.A(\mul1.a[5] ),
    .X(net302));
 sky130_fd_sc_hd__buf_4 fanout303 (.A(net304),
    .X(net303));
 sky130_fd_sc_hd__clkbuf_4 fanout304 (.A(net305),
    .X(net304));
 sky130_fd_sc_hd__clkbuf_8 fanout305 (.A(\mul1.a[4] ),
    .X(net305));
 sky130_fd_sc_hd__buf_4 fanout306 (.A(net307),
    .X(net306));
 sky130_fd_sc_hd__buf_4 fanout307 (.A(\mul1.a[4] ),
    .X(net307));
 sky130_fd_sc_hd__buf_4 fanout308 (.A(net309),
    .X(net308));
 sky130_fd_sc_hd__buf_4 fanout309 (.A(net310),
    .X(net309));
 sky130_fd_sc_hd__clkbuf_8 fanout31 (.A(net38),
    .X(net31));
 sky130_fd_sc_hd__clkbuf_8 fanout310 (.A(\mul1.a[3] ),
    .X(net310));
 sky130_fd_sc_hd__buf_4 fanout311 (.A(net312),
    .X(net311));
 sky130_fd_sc_hd__buf_4 fanout312 (.A(\mul1.a[3] ),
    .X(net312));
 sky130_fd_sc_hd__buf_4 fanout313 (.A(net314),
    .X(net313));
 sky130_fd_sc_hd__clkbuf_4 fanout314 (.A(\mul1.a[2] ),
    .X(net314));
 sky130_fd_sc_hd__buf_4 fanout315 (.A(\mul1.a[2] ),
    .X(net315));
 sky130_fd_sc_hd__buf_4 fanout316 (.A(net317),
    .X(net316));
 sky130_fd_sc_hd__buf_4 fanout317 (.A(\mul1.a[2] ),
    .X(net317));
 sky130_fd_sc_hd__buf_4 fanout318 (.A(net320),
    .X(net318));
 sky130_fd_sc_hd__buf_4 fanout319 (.A(net320),
    .X(net319));
 sky130_fd_sc_hd__clkbuf_8 fanout32 (.A(net33),
    .X(net32));
 sky130_fd_sc_hd__clkbuf_8 fanout320 (.A(\mul1.a[1] ),
    .X(net320));
 sky130_fd_sc_hd__clkbuf_8 fanout321 (.A(\mul1.a[1] ),
    .X(net321));
 sky130_fd_sc_hd__buf_4 fanout322 (.A(net325),
    .X(net322));
 sky130_fd_sc_hd__buf_4 fanout323 (.A(net325),
    .X(net323));
 sky130_fd_sc_hd__clkbuf_8 fanout324 (.A(net325),
    .X(net324));
 sky130_fd_sc_hd__buf_6 fanout325 (.A(\mul1.a[0] ),
    .X(net325));
 sky130_fd_sc_hd__clkbuf_8 fanout326 (.A(\mul0.b[31] ),
    .X(net326));
 sky130_fd_sc_hd__clkbuf_4 fanout327 (.A(net328),
    .X(net327));
 sky130_fd_sc_hd__clkbuf_8 fanout328 (.A(\mul0.b[30] ),
    .X(net328));
 sky130_fd_sc_hd__buf_4 fanout329 (.A(net330),
    .X(net329));
 sky130_fd_sc_hd__clkbuf_8 fanout33 (.A(net38),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_8 fanout330 (.A(\mul0.b[29] ),
    .X(net330));
 sky130_fd_sc_hd__buf_4 fanout331 (.A(net332),
    .X(net331));
 sky130_fd_sc_hd__buf_4 fanout332 (.A(net333),
    .X(net332));
 sky130_fd_sc_hd__buf_4 fanout333 (.A(\mul0.b[28] ),
    .X(net333));
 sky130_fd_sc_hd__buf_4 fanout334 (.A(net335),
    .X(net334));
 sky130_fd_sc_hd__buf_4 fanout335 (.A(net336),
    .X(net335));
 sky130_fd_sc_hd__clkbuf_8 fanout336 (.A(\mul0.b[27] ),
    .X(net336));
 sky130_fd_sc_hd__buf_4 fanout337 (.A(\mul0.b[26] ),
    .X(net337));
 sky130_fd_sc_hd__buf_4 fanout338 (.A(net339),
    .X(net338));
 sky130_fd_sc_hd__clkbuf_4 fanout339 (.A(\mul0.b[26] ),
    .X(net339));
 sky130_fd_sc_hd__clkbuf_8 fanout34 (.A(net38),
    .X(net34));
 sky130_fd_sc_hd__buf_4 fanout340 (.A(net341),
    .X(net340));
 sky130_fd_sc_hd__clkbuf_4 fanout341 (.A(\mul0.b[25] ),
    .X(net341));
 sky130_fd_sc_hd__buf_4 fanout342 (.A(net343),
    .X(net342));
 sky130_fd_sc_hd__clkbuf_4 fanout343 (.A(\mul0.b[25] ),
    .X(net343));
 sky130_fd_sc_hd__buf_4 fanout344 (.A(net345),
    .X(net344));
 sky130_fd_sc_hd__clkbuf_4 fanout345 (.A(\mul0.b[24] ),
    .X(net345));
 sky130_fd_sc_hd__buf_4 fanout346 (.A(net347),
    .X(net346));
 sky130_fd_sc_hd__clkbuf_4 fanout347 (.A(\mul0.b[24] ),
    .X(net347));
 sky130_fd_sc_hd__clkbuf_8 fanout348 (.A(\mul0.b[23] ),
    .X(net348));
 sky130_fd_sc_hd__buf_4 fanout349 (.A(net351),
    .X(net349));
 sky130_fd_sc_hd__clkbuf_4 fanout35 (.A(net38),
    .X(net35));
 sky130_fd_sc_hd__buf_2 fanout350 (.A(net351),
    .X(net350));
 sky130_fd_sc_hd__clkbuf_4 fanout351 (.A(\mul0.b[23] ),
    .X(net351));
 sky130_fd_sc_hd__buf_4 fanout352 (.A(net354),
    .X(net352));
 sky130_fd_sc_hd__buf_4 fanout353 (.A(net354),
    .X(net353));
 sky130_fd_sc_hd__clkbuf_8 fanout354 (.A(net355),
    .X(net354));
 sky130_fd_sc_hd__clkbuf_8 fanout355 (.A(net972),
    .X(net355));
 sky130_fd_sc_hd__buf_6 fanout356 (.A(net360),
    .X(net356));
 sky130_fd_sc_hd__buf_4 fanout357 (.A(net359),
    .X(net357));
 sky130_fd_sc_hd__buf_2 fanout358 (.A(net359),
    .X(net358));
 sky130_fd_sc_hd__clkbuf_4 fanout359 (.A(net360),
    .X(net359));
 sky130_fd_sc_hd__clkbuf_8 fanout36 (.A(net38),
    .X(net36));
 sky130_fd_sc_hd__buf_6 fanout360 (.A(net979),
    .X(net360));
 sky130_fd_sc_hd__clkbuf_4 fanout361 (.A(net362),
    .X(net361));
 sky130_fd_sc_hd__buf_4 fanout362 (.A(net363),
    .X(net362));
 sky130_fd_sc_hd__buf_4 fanout363 (.A(\mul0.b[20] ),
    .X(net363));
 sky130_fd_sc_hd__clkbuf_8 fanout364 (.A(\mul0.b[20] ),
    .X(net364));
 sky130_fd_sc_hd__buf_4 fanout365 (.A(\mul0.b[19] ),
    .X(net365));
 sky130_fd_sc_hd__buf_4 fanout366 (.A(net367),
    .X(net366));
 sky130_fd_sc_hd__clkbuf_4 fanout367 (.A(net369),
    .X(net367));
 sky130_fd_sc_hd__buf_4 fanout368 (.A(net369),
    .X(net368));
 sky130_fd_sc_hd__buf_2 fanout369 (.A(\mul0.b[19] ),
    .X(net369));
 sky130_fd_sc_hd__clkbuf_4 fanout37 (.A(net38),
    .X(net37));
 sky130_fd_sc_hd__buf_4 fanout370 (.A(net371),
    .X(net370));
 sky130_fd_sc_hd__clkbuf_4 fanout371 (.A(\mul0.b[17] ),
    .X(net371));
 sky130_fd_sc_hd__buf_4 fanout372 (.A(\mul0.b[17] ),
    .X(net372));
 sky130_fd_sc_hd__buf_2 fanout373 (.A(\mul0.b[17] ),
    .X(net373));
 sky130_fd_sc_hd__clkbuf_8 fanout374 (.A(\mul0.b[17] ),
    .X(net374));
 sky130_fd_sc_hd__buf_4 fanout375 (.A(net380),
    .X(net375));
 sky130_fd_sc_hd__clkbuf_4 fanout376 (.A(net380),
    .X(net376));
 sky130_fd_sc_hd__buf_4 fanout377 (.A(net380),
    .X(net377));
 sky130_fd_sc_hd__buf_4 fanout378 (.A(net379),
    .X(net378));
 sky130_fd_sc_hd__buf_2 fanout379 (.A(net380),
    .X(net379));
 sky130_fd_sc_hd__buf_4 fanout38 (.A(_02559_),
    .X(net38));
 sky130_fd_sc_hd__buf_4 fanout380 (.A(\mul0.b[16] ),
    .X(net380));
 sky130_fd_sc_hd__buf_4 fanout381 (.A(\mul0.b[15] ),
    .X(net381));
 sky130_fd_sc_hd__clkbuf_4 fanout382 (.A(\mul0.b[15] ),
    .X(net382));
 sky130_fd_sc_hd__clkbuf_8 fanout383 (.A(net385),
    .X(net383));
 sky130_fd_sc_hd__buf_4 fanout384 (.A(net385),
    .X(net384));
 sky130_fd_sc_hd__buf_4 fanout385 (.A(\mul0.b[15] ),
    .X(net385));
 sky130_fd_sc_hd__clkbuf_8 fanout386 (.A(net389),
    .X(net386));
 sky130_fd_sc_hd__buf_4 fanout387 (.A(net389),
    .X(net387));
 sky130_fd_sc_hd__clkbuf_8 fanout388 (.A(net389),
    .X(net388));
 sky130_fd_sc_hd__buf_6 fanout389 (.A(\mul0.b[14] ),
    .X(net389));
 sky130_fd_sc_hd__buf_4 fanout39 (.A(net40),
    .X(net39));
 sky130_fd_sc_hd__buf_4 fanout390 (.A(\mul0.b[13] ),
    .X(net390));
 sky130_fd_sc_hd__clkbuf_4 fanout391 (.A(\mul0.b[13] ),
    .X(net391));
 sky130_fd_sc_hd__clkbuf_8 fanout392 (.A(net394),
    .X(net392));
 sky130_fd_sc_hd__clkbuf_8 fanout393 (.A(net394),
    .X(net393));
 sky130_fd_sc_hd__clkbuf_4 fanout394 (.A(\mul0.b[13] ),
    .X(net394));
 sky130_fd_sc_hd__buf_4 fanout395 (.A(net396),
    .X(net395));
 sky130_fd_sc_hd__buf_4 fanout396 (.A(\mul0.b[12] ),
    .X(net396));
 sky130_fd_sc_hd__buf_4 fanout397 (.A(net399),
    .X(net397));
 sky130_fd_sc_hd__clkbuf_8 fanout398 (.A(net399),
    .X(net398));
 sky130_fd_sc_hd__buf_2 fanout399 (.A(\mul0.b[12] ),
    .X(net399));
 sky130_fd_sc_hd__clkbuf_8 fanout4 (.A(_03055_),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_8 fanout40 (.A(_02499_),
    .X(net40));
 sky130_fd_sc_hd__buf_4 fanout400 (.A(net401),
    .X(net400));
 sky130_fd_sc_hd__buf_4 fanout401 (.A(\mul0.b[11] ),
    .X(net401));
 sky130_fd_sc_hd__clkbuf_8 fanout402 (.A(net403),
    .X(net402));
 sky130_fd_sc_hd__clkbuf_8 fanout403 (.A(\mul0.b[11] ),
    .X(net403));
 sky130_fd_sc_hd__buf_4 fanout404 (.A(net405),
    .X(net404));
 sky130_fd_sc_hd__clkbuf_8 fanout405 (.A(\mul0.b[10] ),
    .X(net405));
 sky130_fd_sc_hd__clkbuf_8 fanout406 (.A(net407),
    .X(net406));
 sky130_fd_sc_hd__buf_6 fanout407 (.A(\mul0.b[10] ),
    .X(net407));
 sky130_fd_sc_hd__buf_4 fanout408 (.A(net412),
    .X(net408));
 sky130_fd_sc_hd__buf_4 fanout409 (.A(net412),
    .X(net409));
 sky130_fd_sc_hd__clkbuf_8 fanout41 (.A(_02498_),
    .X(net41));
 sky130_fd_sc_hd__clkbuf_8 fanout410 (.A(net411),
    .X(net410));
 sky130_fd_sc_hd__clkbuf_8 fanout411 (.A(net412),
    .X(net411));
 sky130_fd_sc_hd__clkbuf_8 fanout412 (.A(\mul0.b[9] ),
    .X(net412));
 sky130_fd_sc_hd__buf_4 fanout413 (.A(net414),
    .X(net413));
 sky130_fd_sc_hd__clkbuf_8 fanout414 (.A(\mul0.b[8] ),
    .X(net414));
 sky130_fd_sc_hd__clkbuf_8 fanout415 (.A(net416),
    .X(net415));
 sky130_fd_sc_hd__clkbuf_8 fanout416 (.A(\mul0.b[8] ),
    .X(net416));
 sky130_fd_sc_hd__buf_4 fanout417 (.A(net418),
    .X(net417));
 sky130_fd_sc_hd__clkbuf_8 fanout418 (.A(\mul0.b[7] ),
    .X(net418));
 sky130_fd_sc_hd__clkbuf_8 fanout419 (.A(net420),
    .X(net419));
 sky130_fd_sc_hd__clkbuf_4 fanout42 (.A(_02498_),
    .X(net42));
 sky130_fd_sc_hd__clkbuf_8 fanout420 (.A(\mul0.b[7] ),
    .X(net420));
 sky130_fd_sc_hd__buf_4 fanout421 (.A(net422),
    .X(net421));
 sky130_fd_sc_hd__clkbuf_8 fanout422 (.A(net425),
    .X(net422));
 sky130_fd_sc_hd__clkbuf_8 fanout423 (.A(net424),
    .X(net423));
 sky130_fd_sc_hd__buf_6 fanout424 (.A(net425),
    .X(net424));
 sky130_fd_sc_hd__buf_4 fanout425 (.A(\mul0.b[6] ),
    .X(net425));
 sky130_fd_sc_hd__buf_4 fanout426 (.A(net427),
    .X(net426));
 sky130_fd_sc_hd__buf_4 fanout427 (.A(\mul0.b[5] ),
    .X(net427));
 sky130_fd_sc_hd__buf_4 fanout428 (.A(net429),
    .X(net428));
 sky130_fd_sc_hd__buf_4 fanout429 (.A(\mul0.b[5] ),
    .X(net429));
 sky130_fd_sc_hd__clkbuf_8 fanout43 (.A(_03051_),
    .X(net43));
 sky130_fd_sc_hd__buf_4 fanout430 (.A(net431),
    .X(net430));
 sky130_fd_sc_hd__clkbuf_4 fanout431 (.A(net432),
    .X(net431));
 sky130_fd_sc_hd__buf_4 fanout432 (.A(\mul0.b[4] ),
    .X(net432));
 sky130_fd_sc_hd__buf_4 fanout433 (.A(net434),
    .X(net433));
 sky130_fd_sc_hd__buf_4 fanout434 (.A(\mul0.b[4] ),
    .X(net434));
 sky130_fd_sc_hd__buf_4 fanout435 (.A(net436),
    .X(net435));
 sky130_fd_sc_hd__buf_4 fanout436 (.A(net437),
    .X(net436));
 sky130_fd_sc_hd__buf_4 fanout437 (.A(\mul0.b[3] ),
    .X(net437));
 sky130_fd_sc_hd__buf_4 fanout438 (.A(net439),
    .X(net438));
 sky130_fd_sc_hd__buf_4 fanout439 (.A(\mul0.b[3] ),
    .X(net439));
 sky130_fd_sc_hd__buf_2 fanout44 (.A(_03051_),
    .X(net44));
 sky130_fd_sc_hd__buf_4 fanout440 (.A(net442),
    .X(net440));
 sky130_fd_sc_hd__buf_2 fanout441 (.A(net442),
    .X(net441));
 sky130_fd_sc_hd__clkbuf_8 fanout442 (.A(\mul0.b[2] ),
    .X(net442));
 sky130_fd_sc_hd__buf_4 fanout443 (.A(net444),
    .X(net443));
 sky130_fd_sc_hd__buf_4 fanout444 (.A(net445),
    .X(net444));
 sky130_fd_sc_hd__buf_2 fanout445 (.A(net446),
    .X(net445));
 sky130_fd_sc_hd__clkbuf_4 fanout446 (.A(\mul0.b[1] ),
    .X(net446));
 sky130_fd_sc_hd__buf_4 fanout447 (.A(\mul0.b[1] ),
    .X(net447));
 sky130_fd_sc_hd__buf_4 fanout448 (.A(net449),
    .X(net448));
 sky130_fd_sc_hd__buf_4 fanout449 (.A(net450),
    .X(net449));
 sky130_fd_sc_hd__buf_4 fanout45 (.A(net46),
    .X(net45));
 sky130_fd_sc_hd__buf_2 fanout450 (.A(net452),
    .X(net450));
 sky130_fd_sc_hd__buf_4 fanout451 (.A(net452),
    .X(net451));
 sky130_fd_sc_hd__clkbuf_8 fanout452 (.A(\mul0.b[0] ),
    .X(net452));
 sky130_fd_sc_hd__clkbuf_8 fanout453 (.A(\mul0.a[31] ),
    .X(net453));
 sky130_fd_sc_hd__clkbuf_4 fanout454 (.A(\mul0.a[31] ),
    .X(net454));
 sky130_fd_sc_hd__buf_4 fanout455 (.A(net456),
    .X(net455));
 sky130_fd_sc_hd__clkbuf_8 fanout456 (.A(net457),
    .X(net456));
 sky130_fd_sc_hd__clkbuf_4 fanout457 (.A(net966),
    .X(net457));
 sky130_fd_sc_hd__buf_4 fanout458 (.A(\mul0.a[29] ),
    .X(net458));
 sky130_fd_sc_hd__buf_4 fanout459 (.A(\mul0.a[29] ),
    .X(net459));
 sky130_fd_sc_hd__clkbuf_8 fanout46 (.A(net49),
    .X(net46));
 sky130_fd_sc_hd__buf_4 fanout460 (.A(net462),
    .X(net460));
 sky130_fd_sc_hd__buf_4 fanout461 (.A(net462),
    .X(net461));
 sky130_fd_sc_hd__clkbuf_8 fanout462 (.A(\mul0.a[28] ),
    .X(net462));
 sky130_fd_sc_hd__clkbuf_8 fanout463 (.A(\mul0.a[27] ),
    .X(net463));
 sky130_fd_sc_hd__clkbuf_4 fanout464 (.A(\mul0.a[27] ),
    .X(net464));
 sky130_fd_sc_hd__clkbuf_8 fanout465 (.A(\mul0.a[27] ),
    .X(net465));
 sky130_fd_sc_hd__clkbuf_8 fanout466 (.A(net469),
    .X(net466));
 sky130_fd_sc_hd__clkbuf_4 fanout467 (.A(net469),
    .X(net467));
 sky130_fd_sc_hd__buf_4 fanout468 (.A(net469),
    .X(net468));
 sky130_fd_sc_hd__buf_4 fanout469 (.A(\mul0.a[26] ),
    .X(net469));
 sky130_fd_sc_hd__buf_4 fanout47 (.A(net49),
    .X(net47));
 sky130_fd_sc_hd__clkbuf_8 fanout470 (.A(net473),
    .X(net470));
 sky130_fd_sc_hd__clkbuf_8 fanout471 (.A(net473),
    .X(net471));
 sky130_fd_sc_hd__buf_2 fanout472 (.A(net473),
    .X(net472));
 sky130_fd_sc_hd__buf_4 fanout473 (.A(\mul0.a[25] ),
    .X(net473));
 sky130_fd_sc_hd__buf_4 fanout474 (.A(net477),
    .X(net474));
 sky130_fd_sc_hd__clkbuf_8 fanout475 (.A(net477),
    .X(net475));
 sky130_fd_sc_hd__clkbuf_4 fanout476 (.A(net477),
    .X(net476));
 sky130_fd_sc_hd__buf_4 fanout477 (.A(\mul0.a[24] ),
    .X(net477));
 sky130_fd_sc_hd__buf_4 fanout478 (.A(net481),
    .X(net478));
 sky130_fd_sc_hd__clkbuf_8 fanout479 (.A(net481),
    .X(net479));
 sky130_fd_sc_hd__buf_4 fanout48 (.A(net49),
    .X(net48));
 sky130_fd_sc_hd__clkbuf_4 fanout480 (.A(net481),
    .X(net480));
 sky130_fd_sc_hd__buf_4 fanout481 (.A(\mul0.a[23] ),
    .X(net481));
 sky130_fd_sc_hd__clkbuf_8 fanout482 (.A(\mul0.a[22] ),
    .X(net482));
 sky130_fd_sc_hd__buf_4 fanout483 (.A(\mul0.a[22] ),
    .X(net483));
 sky130_fd_sc_hd__buf_4 fanout484 (.A(\mul0.a[22] ),
    .X(net484));
 sky130_fd_sc_hd__clkbuf_4 fanout485 (.A(\mul0.a[22] ),
    .X(net485));
 sky130_fd_sc_hd__clkbuf_8 fanout486 (.A(\mul0.a[21] ),
    .X(net486));
 sky130_fd_sc_hd__clkbuf_4 fanout487 (.A(\mul0.a[21] ),
    .X(net487));
 sky130_fd_sc_hd__buf_4 fanout488 (.A(\mul0.a[21] ),
    .X(net488));
 sky130_fd_sc_hd__clkbuf_4 fanout489 (.A(\mul0.a[21] ),
    .X(net489));
 sky130_fd_sc_hd__clkbuf_4 fanout49 (.A(_02754_),
    .X(net49));
 sky130_fd_sc_hd__clkbuf_8 fanout490 (.A(\mul0.a[20] ),
    .X(net490));
 sky130_fd_sc_hd__buf_4 fanout491 (.A(\mul0.a[20] ),
    .X(net491));
 sky130_fd_sc_hd__buf_4 fanout492 (.A(net493),
    .X(net492));
 sky130_fd_sc_hd__buf_4 fanout493 (.A(\mul0.a[20] ),
    .X(net493));
 sky130_fd_sc_hd__clkbuf_8 fanout494 (.A(\mul0.a[19] ),
    .X(net494));
 sky130_fd_sc_hd__buf_4 fanout495 (.A(\mul0.a[19] ),
    .X(net495));
 sky130_fd_sc_hd__buf_4 fanout496 (.A(net497),
    .X(net496));
 sky130_fd_sc_hd__buf_4 fanout497 (.A(\mul0.a[19] ),
    .X(net497));
 sky130_fd_sc_hd__buf_4 fanout498 (.A(net499),
    .X(net498));
 sky130_fd_sc_hd__clkbuf_8 fanout499 (.A(\mul0.a[18] ),
    .X(net499));
 sky130_fd_sc_hd__clkbuf_8 fanout5 (.A(net6),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_8 fanout50 (.A(_02753_),
    .X(net50));
 sky130_fd_sc_hd__buf_4 fanout500 (.A(net501),
    .X(net500));
 sky130_fd_sc_hd__buf_2 fanout501 (.A(net502),
    .X(net501));
 sky130_fd_sc_hd__clkbuf_4 fanout502 (.A(\mul0.a[18] ),
    .X(net502));
 sky130_fd_sc_hd__buf_4 fanout503 (.A(\mul0.a[17] ),
    .X(net503));
 sky130_fd_sc_hd__buf_4 fanout504 (.A(\mul0.a[17] ),
    .X(net504));
 sky130_fd_sc_hd__buf_4 fanout505 (.A(net506),
    .X(net505));
 sky130_fd_sc_hd__buf_4 fanout506 (.A(\mul0.a[17] ),
    .X(net506));
 sky130_fd_sc_hd__buf_4 fanout507 (.A(net508),
    .X(net507));
 sky130_fd_sc_hd__clkbuf_8 fanout508 (.A(\mul0.a[16] ),
    .X(net508));
 sky130_fd_sc_hd__buf_4 fanout509 (.A(net510),
    .X(net509));
 sky130_fd_sc_hd__buf_4 fanout51 (.A(_02753_),
    .X(net51));
 sky130_fd_sc_hd__buf_4 fanout510 (.A(\mul0.a[16] ),
    .X(net510));
 sky130_fd_sc_hd__clkbuf_8 fanout511 (.A(net512),
    .X(net511));
 sky130_fd_sc_hd__clkbuf_8 fanout512 (.A(\mul0.a[15] ),
    .X(net512));
 sky130_fd_sc_hd__buf_4 fanout513 (.A(\mul0.a[15] ),
    .X(net513));
 sky130_fd_sc_hd__buf_4 fanout514 (.A(\mul0.a[15] ),
    .X(net514));
 sky130_fd_sc_hd__buf_4 fanout515 (.A(net516),
    .X(net515));
 sky130_fd_sc_hd__clkbuf_4 fanout516 (.A(net517),
    .X(net516));
 sky130_fd_sc_hd__buf_4 fanout517 (.A(\mul0.a[14] ),
    .X(net517));
 sky130_fd_sc_hd__clkbuf_4 fanout518 (.A(\mul0.a[14] ),
    .X(net518));
 sky130_fd_sc_hd__buf_4 fanout519 (.A(\mul0.a[14] ),
    .X(net519));
 sky130_fd_sc_hd__clkbuf_8 fanout52 (.A(net53),
    .X(net52));
 sky130_fd_sc_hd__buf_4 fanout520 (.A(net521),
    .X(net520));
 sky130_fd_sc_hd__clkbuf_8 fanout521 (.A(net524),
    .X(net521));
 sky130_fd_sc_hd__buf_4 fanout522 (.A(net523),
    .X(net522));
 sky130_fd_sc_hd__buf_4 fanout523 (.A(net524),
    .X(net523));
 sky130_fd_sc_hd__buf_4 fanout524 (.A(\mul0.a[13] ),
    .X(net524));
 sky130_fd_sc_hd__buf_4 fanout525 (.A(net527),
    .X(net525));
 sky130_fd_sc_hd__clkbuf_2 fanout526 (.A(net527),
    .X(net526));
 sky130_fd_sc_hd__clkbuf_8 fanout527 (.A(\mul0.a[12] ),
    .X(net527));
 sky130_fd_sc_hd__buf_4 fanout528 (.A(net529),
    .X(net528));
 sky130_fd_sc_hd__clkbuf_4 fanout529 (.A(\mul0.a[12] ),
    .X(net529));
 sky130_fd_sc_hd__clkbuf_8 fanout53 (.A(_02752_),
    .X(net53));
 sky130_fd_sc_hd__buf_4 fanout530 (.A(net531),
    .X(net530));
 sky130_fd_sc_hd__clkbuf_4 fanout531 (.A(net532),
    .X(net531));
 sky130_fd_sc_hd__buf_4 fanout532 (.A(\mul0.a[11] ),
    .X(net532));
 sky130_fd_sc_hd__buf_4 fanout533 (.A(\mul0.a[11] ),
    .X(net533));
 sky130_fd_sc_hd__clkbuf_4 fanout534 (.A(\mul0.a[11] ),
    .X(net534));
 sky130_fd_sc_hd__buf_4 fanout535 (.A(net536),
    .X(net535));
 sky130_fd_sc_hd__buf_4 fanout536 (.A(net537),
    .X(net536));
 sky130_fd_sc_hd__buf_4 fanout537 (.A(net539),
    .X(net537));
 sky130_fd_sc_hd__clkbuf_8 fanout538 (.A(net539),
    .X(net538));
 sky130_fd_sc_hd__buf_4 fanout539 (.A(\mul0.a[10] ),
    .X(net539));
 sky130_fd_sc_hd__clkbuf_8 fanout54 (.A(net55),
    .X(net54));
 sky130_fd_sc_hd__buf_4 fanout540 (.A(net541),
    .X(net540));
 sky130_fd_sc_hd__buf_4 fanout541 (.A(net542),
    .X(net541));
 sky130_fd_sc_hd__clkbuf_8 fanout542 (.A(\mul0.a[9] ),
    .X(net542));
 sky130_fd_sc_hd__clkbuf_8 fanout543 (.A(\mul0.a[9] ),
    .X(net543));
 sky130_fd_sc_hd__buf_4 fanout544 (.A(net545),
    .X(net544));
 sky130_fd_sc_hd__clkbuf_8 fanout545 (.A(\mul0.a[8] ),
    .X(net545));
 sky130_fd_sc_hd__clkbuf_8 fanout546 (.A(\mul0.a[8] ),
    .X(net546));
 sky130_fd_sc_hd__clkbuf_8 fanout547 (.A(\mul0.a[8] ),
    .X(net547));
 sky130_fd_sc_hd__buf_4 fanout548 (.A(net549),
    .X(net548));
 sky130_fd_sc_hd__clkbuf_8 fanout549 (.A(net550),
    .X(net549));
 sky130_fd_sc_hd__clkbuf_8 fanout55 (.A(_02736_),
    .X(net55));
 sky130_fd_sc_hd__clkbuf_8 fanout550 (.A(\mul0.a[7] ),
    .X(net550));
 sky130_fd_sc_hd__clkbuf_8 fanout551 (.A(\mul0.a[7] ),
    .X(net551));
 sky130_fd_sc_hd__buf_4 fanout552 (.A(net553),
    .X(net552));
 sky130_fd_sc_hd__clkbuf_8 fanout553 (.A(net554),
    .X(net553));
 sky130_fd_sc_hd__clkbuf_8 fanout554 (.A(net556),
    .X(net554));
 sky130_fd_sc_hd__clkbuf_8 fanout555 (.A(net556),
    .X(net555));
 sky130_fd_sc_hd__buf_4 fanout556 (.A(\mul0.a[6] ),
    .X(net556));
 sky130_fd_sc_hd__buf_4 fanout557 (.A(net558),
    .X(net557));
 sky130_fd_sc_hd__clkbuf_8 fanout558 (.A(\mul0.a[5] ),
    .X(net558));
 sky130_fd_sc_hd__buf_4 fanout559 (.A(net560),
    .X(net559));
 sky130_fd_sc_hd__buf_4 fanout56 (.A(_02568_),
    .X(net56));
 sky130_fd_sc_hd__buf_4 fanout560 (.A(\mul0.a[5] ),
    .X(net560));
 sky130_fd_sc_hd__clkbuf_8 fanout561 (.A(net565),
    .X(net561));
 sky130_fd_sc_hd__buf_4 fanout562 (.A(net563),
    .X(net562));
 sky130_fd_sc_hd__clkbuf_4 fanout563 (.A(net564),
    .X(net563));
 sky130_fd_sc_hd__buf_4 fanout564 (.A(net565),
    .X(net564));
 sky130_fd_sc_hd__clkbuf_4 fanout565 (.A(\mul0.a[4] ),
    .X(net565));
 sky130_fd_sc_hd__buf_4 fanout566 (.A(net570),
    .X(net566));
 sky130_fd_sc_hd__buf_4 fanout567 (.A(net570),
    .X(net567));
 sky130_fd_sc_hd__buf_4 fanout568 (.A(net569),
    .X(net568));
 sky130_fd_sc_hd__clkbuf_4 fanout569 (.A(net570),
    .X(net569));
 sky130_fd_sc_hd__buf_4 fanout57 (.A(_02567_),
    .X(net57));
 sky130_fd_sc_hd__clkbuf_4 fanout570 (.A(\mul0.a[3] ),
    .X(net570));
 sky130_fd_sc_hd__buf_4 fanout571 (.A(net575),
    .X(net571));
 sky130_fd_sc_hd__buf_4 fanout572 (.A(net575),
    .X(net572));
 sky130_fd_sc_hd__buf_4 fanout573 (.A(net574),
    .X(net573));
 sky130_fd_sc_hd__buf_4 fanout574 (.A(net575),
    .X(net574));
 sky130_fd_sc_hd__buf_4 fanout575 (.A(\mul0.a[2] ),
    .X(net575));
 sky130_fd_sc_hd__buf_4 fanout576 (.A(\mul0.a[1] ),
    .X(net576));
 sky130_fd_sc_hd__buf_4 fanout577 (.A(net580),
    .X(net577));
 sky130_fd_sc_hd__buf_4 fanout578 (.A(net580),
    .X(net578));
 sky130_fd_sc_hd__buf_2 fanout579 (.A(net580),
    .X(net579));
 sky130_fd_sc_hd__buf_4 fanout58 (.A(net59),
    .X(net58));
 sky130_fd_sc_hd__buf_4 fanout580 (.A(\mul0.a[1] ),
    .X(net580));
 sky130_fd_sc_hd__buf_4 fanout581 (.A(net582),
    .X(net581));
 sky130_fd_sc_hd__clkbuf_8 fanout582 (.A(net584),
    .X(net582));
 sky130_fd_sc_hd__buf_4 fanout583 (.A(net584),
    .X(net583));
 sky130_fd_sc_hd__buf_4 fanout584 (.A(\mul0.a[0] ),
    .X(net584));
 sky130_fd_sc_hd__buf_4 fanout585 (.A(net586),
    .X(net585));
 sky130_fd_sc_hd__buf_4 fanout586 (.A(net587),
    .X(net586));
 sky130_fd_sc_hd__buf_6 fanout587 (.A(net592),
    .X(net587));
 sky130_fd_sc_hd__buf_4 fanout588 (.A(net592),
    .X(net588));
 sky130_fd_sc_hd__buf_2 fanout589 (.A(net592),
    .X(net589));
 sky130_fd_sc_hd__buf_4 fanout59 (.A(_02561_),
    .X(net59));
 sky130_fd_sc_hd__buf_4 fanout590 (.A(net591),
    .X(net590));
 sky130_fd_sc_hd__buf_4 fanout591 (.A(net592),
    .X(net591));
 sky130_fd_sc_hd__buf_8 fanout592 (.A(\state[8] ),
    .X(net592));
 sky130_fd_sc_hd__buf_4 fanout593 (.A(net598),
    .X(net593));
 sky130_fd_sc_hd__buf_2 fanout594 (.A(net598),
    .X(net594));
 sky130_fd_sc_hd__clkbuf_8 fanout595 (.A(net596),
    .X(net595));
 sky130_fd_sc_hd__buf_4 fanout596 (.A(net597),
    .X(net596));
 sky130_fd_sc_hd__buf_4 fanout597 (.A(net598),
    .X(net597));
 sky130_fd_sc_hd__buf_8 fanout598 (.A(\state[7] ),
    .X(net598));
 sky130_fd_sc_hd__buf_6 fanout599 (.A(net600),
    .X(net599));
 sky130_fd_sc_hd__clkbuf_8 fanout6 (.A(_03794_),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_8 fanout60 (.A(net61),
    .X(net60));
 sky130_fd_sc_hd__clkbuf_8 fanout600 (.A(\state[4] ),
    .X(net600));
 sky130_fd_sc_hd__clkbuf_8 fanout601 (.A(net606),
    .X(net601));
 sky130_fd_sc_hd__buf_4 fanout602 (.A(net606),
    .X(net602));
 sky130_fd_sc_hd__buf_2 fanout603 (.A(net606),
    .X(net603));
 sky130_fd_sc_hd__buf_4 fanout604 (.A(net606),
    .X(net604));
 sky130_fd_sc_hd__buf_2 fanout605 (.A(net606),
    .X(net605));
 sky130_fd_sc_hd__clkbuf_8 fanout606 (.A(\state[3] ),
    .X(net606));
 sky130_fd_sc_hd__clkbuf_8 fanout607 (.A(\state[2] ),
    .X(net607));
 sky130_fd_sc_hd__buf_4 fanout608 (.A(\state[2] ),
    .X(net608));
 sky130_fd_sc_hd__buf_2 fanout609 (.A(\state[2] ),
    .X(net609));
 sky130_fd_sc_hd__buf_6 fanout61 (.A(_02561_),
    .X(net61));
 sky130_fd_sc_hd__buf_4 fanout610 (.A(\state[2] ),
    .X(net610));
 sky130_fd_sc_hd__clkbuf_4 fanout611 (.A(\state[2] ),
    .X(net611));
 sky130_fd_sc_hd__clkbuf_8 fanout612 (.A(net616),
    .X(net612));
 sky130_fd_sc_hd__clkbuf_4 fanout613 (.A(net616),
    .X(net613));
 sky130_fd_sc_hd__clkbuf_8 fanout614 (.A(net616),
    .X(net614));
 sky130_fd_sc_hd__clkbuf_8 fanout615 (.A(net616),
    .X(net615));
 sky130_fd_sc_hd__clkbuf_4 fanout616 (.A(\state[1] ),
    .X(net616));
 sky130_fd_sc_hd__clkbuf_8 fanout617 (.A(\state[1] ),
    .X(net617));
 sky130_fd_sc_hd__clkbuf_4 fanout618 (.A(\state[1] ),
    .X(net618));
 sky130_fd_sc_hd__clkbuf_8 fanout619 (.A(\state[1] ),
    .X(net619));
 sky130_fd_sc_hd__buf_6 fanout62 (.A(\mul1.b[31] ),
    .X(net62));
 sky130_fd_sc_hd__buf_4 fanout620 (.A(\state[1] ),
    .X(net620));
 sky130_fd_sc_hd__buf_4 fanout621 (.A(net622),
    .X(net621));
 sky130_fd_sc_hd__buf_4 fanout622 (.A(\mul1.b[0] ),
    .X(net622));
 sky130_fd_sc_hd__buf_4 fanout623 (.A(net625),
    .X(net623));
 sky130_fd_sc_hd__clkbuf_4 fanout624 (.A(net625),
    .X(net624));
 sky130_fd_sc_hd__buf_4 fanout625 (.A(\mul1.b[0] ),
    .X(net625));
 sky130_fd_sc_hd__clkbuf_8 fanout626 (.A(net629),
    .X(net626));
 sky130_fd_sc_hd__buf_2 fanout627 (.A(net629),
    .X(net627));
 sky130_fd_sc_hd__buf_4 fanout628 (.A(net629),
    .X(net628));
 sky130_fd_sc_hd__clkbuf_8 fanout629 (.A(net630),
    .X(net629));
 sky130_fd_sc_hd__clkbuf_4 fanout63 (.A(net65),
    .X(net63));
 sky130_fd_sc_hd__buf_8 fanout630 (.A(\mul1.a[16] ),
    .X(net630));
 sky130_fd_sc_hd__clkbuf_8 fanout631 (.A(\mul0.b[18] ),
    .X(net631));
 sky130_fd_sc_hd__buf_4 fanout632 (.A(\mul0.b[18] ),
    .X(net632));
 sky130_fd_sc_hd__buf_2 fanout633 (.A(\mul0.b[18] ),
    .X(net633));
 sky130_fd_sc_hd__buf_4 fanout634 (.A(net635),
    .X(net634));
 sky130_fd_sc_hd__clkbuf_4 fanout635 (.A(\mul0.b[18] ),
    .X(net635));
 sky130_fd_sc_hd__clkbuf_8 fanout636 (.A(net638),
    .X(net636));
 sky130_fd_sc_hd__clkbuf_8 fanout637 (.A(net638),
    .X(net637));
 sky130_fd_sc_hd__buf_4 fanout638 (.A(net639),
    .X(net638));
 sky130_fd_sc_hd__clkbuf_8 fanout639 (.A(net646),
    .X(net639));
 sky130_fd_sc_hd__buf_2 fanout64 (.A(net65),
    .X(net64));
 sky130_fd_sc_hd__clkbuf_8 fanout640 (.A(net642),
    .X(net640));
 sky130_fd_sc_hd__clkbuf_8 fanout641 (.A(net642),
    .X(net641));
 sky130_fd_sc_hd__clkbuf_4 fanout642 (.A(net645),
    .X(net642));
 sky130_fd_sc_hd__clkbuf_8 fanout643 (.A(net645),
    .X(net643));
 sky130_fd_sc_hd__clkbuf_8 fanout644 (.A(net645),
    .X(net644));
 sky130_fd_sc_hd__buf_4 fanout645 (.A(net646),
    .X(net645));
 sky130_fd_sc_hd__buf_12 fanout646 (.A(nrst_i),
    .X(net646));
 sky130_fd_sc_hd__buf_4 fanout65 (.A(net967),
    .X(net65));
 sky130_fd_sc_hd__buf_4 fanout66 (.A(net67),
    .X(net66));
 sky130_fd_sc_hd__buf_4 fanout67 (.A(net68),
    .X(net67));
 sky130_fd_sc_hd__clkbuf_4 fanout68 (.A(net971),
    .X(net68));
 sky130_fd_sc_hd__buf_4 fanout69 (.A(net70),
    .X(net69));
 sky130_fd_sc_hd__buf_4 fanout7 (.A(net8),
    .X(net7));
 sky130_fd_sc_hd__buf_4 fanout70 (.A(net71),
    .X(net70));
 sky130_fd_sc_hd__buf_4 fanout71 (.A(net975),
    .X(net71));
 sky130_fd_sc_hd__buf_4 fanout72 (.A(net73),
    .X(net72));
 sky130_fd_sc_hd__buf_4 fanout73 (.A(\mul1.b[27] ),
    .X(net73));
 sky130_fd_sc_hd__clkbuf_8 fanout74 (.A(\mul1.b[27] ),
    .X(net74));
 sky130_fd_sc_hd__buf_4 fanout75 (.A(\mul1.b[26] ),
    .X(net75));
 sky130_fd_sc_hd__buf_4 fanout76 (.A(net77),
    .X(net76));
 sky130_fd_sc_hd__buf_4 fanout77 (.A(\mul1.b[26] ),
    .X(net77));
 sky130_fd_sc_hd__buf_4 fanout78 (.A(\mul1.b[25] ),
    .X(net78));
 sky130_fd_sc_hd__buf_4 fanout79 (.A(net80),
    .X(net79));
 sky130_fd_sc_hd__clkbuf_8 fanout8 (.A(_03053_),
    .X(net8));
 sky130_fd_sc_hd__buf_4 fanout80 (.A(\mul1.b[25] ),
    .X(net80));
 sky130_fd_sc_hd__buf_4 fanout81 (.A(net82),
    .X(net81));
 sky130_fd_sc_hd__clkbuf_4 fanout82 (.A(\mul1.b[24] ),
    .X(net82));
 sky130_fd_sc_hd__buf_4 fanout83 (.A(net84),
    .X(net83));
 sky130_fd_sc_hd__buf_4 fanout84 (.A(\mul1.b[24] ),
    .X(net84));
 sky130_fd_sc_hd__clkbuf_8 fanout85 (.A(net88),
    .X(net85));
 sky130_fd_sc_hd__buf_4 fanout86 (.A(net87),
    .X(net86));
 sky130_fd_sc_hd__buf_4 fanout87 (.A(net88),
    .X(net87));
 sky130_fd_sc_hd__buf_4 fanout88 (.A(\mul1.b[23] ),
    .X(net88));
 sky130_fd_sc_hd__clkbuf_8 fanout89 (.A(net90),
    .X(net89));
 sky130_fd_sc_hd__clkbuf_8 fanout9 (.A(_03057_),
    .X(net9));
 sky130_fd_sc_hd__buf_4 fanout90 (.A(\mul1.b[22] ),
    .X(net90));
 sky130_fd_sc_hd__clkbuf_8 fanout91 (.A(\mul1.b[22] ),
    .X(net91));
 sky130_fd_sc_hd__clkbuf_4 fanout92 (.A(\mul1.b[22] ),
    .X(net92));
 sky130_fd_sc_hd__clkbuf_8 fanout93 (.A(net94),
    .X(net93));
 sky130_fd_sc_hd__buf_4 fanout94 (.A(net96),
    .X(net94));
 sky130_fd_sc_hd__clkbuf_8 fanout95 (.A(net96),
    .X(net95));
 sky130_fd_sc_hd__buf_4 fanout96 (.A(\mul1.b[21] ),
    .X(net96));
 sky130_fd_sc_hd__buf_6 fanout97 (.A(\mul1.b[21] ),
    .X(net97));
 sky130_fd_sc_hd__clkbuf_8 fanout98 (.A(\mul1.b[20] ),
    .X(net98));
 sky130_fd_sc_hd__buf_4 fanout99 (.A(net100),
    .X(net99));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1 (.A(\state[5] ),
    .X(net647));
 sky130_fd_sc_hd__dlygate4sd3_1 hold10 (.A(\tx[14] ),
    .X(net656));
 sky130_fd_sc_hd__dlygate4sd3_1 hold100 (.A(\add0.b_i[28] ),
    .X(net746));
 sky130_fd_sc_hd__dlygate4sd3_1 hold101 (.A(\add0.b_i[23] ),
    .X(net747));
 sky130_fd_sc_hd__dlygate4sd3_1 hold102 (.A(\add0.a_i[19] ),
    .X(net748));
 sky130_fd_sc_hd__dlygate4sd3_1 hold103 (.A(_00286_),
    .X(net749));
 sky130_fd_sc_hd__dlygate4sd3_1 hold104 (.A(\add0.b_i[7] ),
    .X(net750));
 sky130_fd_sc_hd__dlygate4sd3_1 hold105 (.A(_00306_),
    .X(net751));
 sky130_fd_sc_hd__dlygate4sd3_1 hold106 (.A(\depth[15] ),
    .X(net752));
 sky130_fd_sc_hd__dlygate4sd3_1 hold107 (.A(\add0.a_i[7] ),
    .X(net753));
 sky130_fd_sc_hd__dlygate4sd3_1 hold108 (.A(_00274_),
    .X(net754));
 sky130_fd_sc_hd__dlygate4sd3_1 hold109 (.A(\add0.a_i[22] ),
    .X(net755));
 sky130_fd_sc_hd__dlygate4sd3_1 hold11 (.A(\tx[3] ),
    .X(net657));
 sky130_fd_sc_hd__dlygate4sd3_1 hold110 (.A(_00289_),
    .X(net756));
 sky130_fd_sc_hd__dlygate4sd3_1 hold111 (.A(\temp[17] ),
    .X(net757));
 sky130_fd_sc_hd__dlygate4sd3_1 hold112 (.A(\temp[25] ),
    .X(net758));
 sky130_fd_sc_hd__dlygate4sd3_1 hold113 (.A(\add0.a_i[2] ),
    .X(net759));
 sky130_fd_sc_hd__dlygate4sd3_1 hold114 (.A(_00269_),
    .X(net760));
 sky130_fd_sc_hd__dlygate4sd3_1 hold115 (.A(\add0.b_i[13] ),
    .X(net761));
 sky130_fd_sc_hd__dlygate4sd3_1 hold116 (.A(\in_data[54] ),
    .X(net762));
 sky130_fd_sc_hd__dlygate4sd3_1 hold117 (.A(\temp[27] ),
    .X(net763));
 sky130_fd_sc_hd__dlygate4sd3_1 hold118 (.A(\temp[15] ),
    .X(net764));
 sky130_fd_sc_hd__dlygate4sd3_1 hold119 (.A(\in_data[26] ),
    .X(net765));
 sky130_fd_sc_hd__dlygate4sd3_1 hold12 (.A(\depth[26] ),
    .X(net658));
 sky130_fd_sc_hd__dlygate4sd3_1 hold120 (.A(\in_data[30] ),
    .X(net766));
 sky130_fd_sc_hd__dlygate4sd3_1 hold121 (.A(\add0.b_i[31] ),
    .X(net767));
 sky130_fd_sc_hd__dlygate4sd3_1 hold122 (.A(\add0.b_i[9] ),
    .X(net768));
 sky130_fd_sc_hd__dlygate4sd3_1 hold123 (.A(\in_data[44] ),
    .X(net769));
 sky130_fd_sc_hd__dlygate4sd3_1 hold124 (.A(\temp[26] ),
    .X(net770));
 sky130_fd_sc_hd__dlygate4sd3_1 hold125 (.A(\temp[3] ),
    .X(net771));
 sky130_fd_sc_hd__dlygate4sd3_1 hold126 (.A(\add0.b_i[19] ),
    .X(net772));
 sky130_fd_sc_hd__dlygate4sd3_1 hold127 (.A(_00318_),
    .X(net773));
 sky130_fd_sc_hd__dlygate4sd3_1 hold128 (.A(\add0.a_i[29] ),
    .X(net774));
 sky130_fd_sc_hd__dlygate4sd3_1 hold129 (.A(_00296_),
    .X(net775));
 sky130_fd_sc_hd__dlygate4sd3_1 hold13 (.A(\depth[0] ),
    .X(net659));
 sky130_fd_sc_hd__dlygate4sd3_1 hold130 (.A(\in_data[56] ),
    .X(net776));
 sky130_fd_sc_hd__dlygate4sd3_1 hold131 (.A(\in_data[53] ),
    .X(net777));
 sky130_fd_sc_hd__dlygate4sd3_1 hold132 (.A(\temp[1] ),
    .X(net778));
 sky130_fd_sc_hd__dlygate4sd3_1 hold133 (.A(\add0.a_i[13] ),
    .X(net779));
 sky130_fd_sc_hd__dlygate4sd3_1 hold134 (.A(\add0.b_i[2] ),
    .X(net780));
 sky130_fd_sc_hd__dlygate4sd3_1 hold135 (.A(_00301_),
    .X(net781));
 sky130_fd_sc_hd__dlygate4sd3_1 hold136 (.A(\temp[10] ),
    .X(net782));
 sky130_fd_sc_hd__dlygate4sd3_1 hold137 (.A(\add0.b_i[18] ),
    .X(net783));
 sky130_fd_sc_hd__dlygate4sd3_1 hold138 (.A(_00317_),
    .X(net784));
 sky130_fd_sc_hd__dlygate4sd3_1 hold139 (.A(\in_data[37] ),
    .X(net785));
 sky130_fd_sc_hd__dlygate4sd3_1 hold14 (.A(\tx[20] ),
    .X(net660));
 sky130_fd_sc_hd__dlygate4sd3_1 hold140 (.A(\add0.a_i[14] ),
    .X(net786));
 sky130_fd_sc_hd__dlygate4sd3_1 hold141 (.A(_00281_),
    .X(net787));
 sky130_fd_sc_hd__dlygate4sd3_1 hold142 (.A(\in_data[51] ),
    .X(net788));
 sky130_fd_sc_hd__dlygate4sd3_1 hold143 (.A(\tx[2] ),
    .X(net789));
 sky130_fd_sc_hd__dlygate4sd3_1 hold144 (.A(\depth[19] ),
    .X(net790));
 sky130_fd_sc_hd__dlygate4sd3_1 hold145 (.A(\add0.b_i[27] ),
    .X(net791));
 sky130_fd_sc_hd__dlygate4sd3_1 hold146 (.A(\add0.b_i[29] ),
    .X(net792));
 sky130_fd_sc_hd__dlygate4sd3_1 hold147 (.A(_00328_),
    .X(net793));
 sky130_fd_sc_hd__dlygate4sd3_1 hold148 (.A(\in_data[31] ),
    .X(net794));
 sky130_fd_sc_hd__dlygate4sd3_1 hold149 (.A(\in_data[71] ),
    .X(net795));
 sky130_fd_sc_hd__dlygate4sd3_1 hold15 (.A(\depth[5] ),
    .X(net661));
 sky130_fd_sc_hd__dlygate4sd3_1 hold150 (.A(\temp[12] ),
    .X(net796));
 sky130_fd_sc_hd__dlygate4sd3_1 hold151 (.A(\add0.b_i[11] ),
    .X(net797));
 sky130_fd_sc_hd__dlygate4sd3_1 hold152 (.A(\depth[12] ),
    .X(net798));
 sky130_fd_sc_hd__dlygate4sd3_1 hold153 (.A(\in_data[47] ),
    .X(net799));
 sky130_fd_sc_hd__dlygate4sd3_1 hold154 (.A(\in_data[48] ),
    .X(net800));
 sky130_fd_sc_hd__dlygate4sd3_1 hold155 (.A(\temp[7] ),
    .X(net801));
 sky130_fd_sc_hd__dlygate4sd3_1 hold156 (.A(\temp[0] ),
    .X(net802));
 sky130_fd_sc_hd__dlygate4sd3_1 hold157 (.A(\add0.a_i[15] ),
    .X(net803));
 sky130_fd_sc_hd__dlygate4sd3_1 hold158 (.A(\add0.b_i[22] ),
    .X(net804));
 sky130_fd_sc_hd__dlygate4sd3_1 hold159 (.A(_00321_),
    .X(net805));
 sky130_fd_sc_hd__dlygate4sd3_1 hold16 (.A(\depth[6] ),
    .X(net662));
 sky130_fd_sc_hd__dlygate4sd3_1 hold160 (.A(\in_data[32] ),
    .X(net806));
 sky130_fd_sc_hd__dlygate4sd3_1 hold161 (.A(\in_data[59] ),
    .X(net807));
 sky130_fd_sc_hd__dlygate4sd3_1 hold162 (.A(\in_data[50] ),
    .X(net808));
 sky130_fd_sc_hd__dlygate4sd3_1 hold163 (.A(\temp[5] ),
    .X(net809));
 sky130_fd_sc_hd__dlygate4sd3_1 hold164 (.A(\in_data[55] ),
    .X(net810));
 sky130_fd_sc_hd__dlygate4sd3_1 hold165 (.A(\in_data[68] ),
    .X(net811));
 sky130_fd_sc_hd__dlygate4sd3_1 hold166 (.A(\in_data[52] ),
    .X(net812));
 sky130_fd_sc_hd__dlygate4sd3_1 hold167 (.A(\temp[22] ),
    .X(net813));
 sky130_fd_sc_hd__dlygate4sd3_1 hold168 (.A(\depth[22] ),
    .X(net814));
 sky130_fd_sc_hd__dlygate4sd3_1 hold169 (.A(\temp[18] ),
    .X(net815));
 sky130_fd_sc_hd__dlygate4sd3_1 hold17 (.A(\depth[18] ),
    .X(net663));
 sky130_fd_sc_hd__dlygate4sd3_1 hold170 (.A(\in_data[45] ),
    .X(net816));
 sky130_fd_sc_hd__dlygate4sd3_1 hold171 (.A(\add0.b_i[30] ),
    .X(net817));
 sky130_fd_sc_hd__dlygate4sd3_1 hold172 (.A(_00329_),
    .X(net818));
 sky130_fd_sc_hd__dlygate4sd3_1 hold173 (.A(\depth[9] ),
    .X(net819));
 sky130_fd_sc_hd__dlygate4sd3_1 hold174 (.A(\temp[19] ),
    .X(net820));
 sky130_fd_sc_hd__dlygate4sd3_1 hold175 (.A(\in_data[29] ),
    .X(net821));
 sky130_fd_sc_hd__dlygate4sd3_1 hold176 (.A(\in_data[66] ),
    .X(net822));
 sky130_fd_sc_hd__dlygate4sd3_1 hold177 (.A(\in_data[36] ),
    .X(net823));
 sky130_fd_sc_hd__dlygate4sd3_1 hold178 (.A(\in_data[58] ),
    .X(net824));
 sky130_fd_sc_hd__dlygate4sd3_1 hold179 (.A(\in_data[70] ),
    .X(net825));
 sky130_fd_sc_hd__dlygate4sd3_1 hold18 (.A(\tx[22] ),
    .X(net664));
 sky130_fd_sc_hd__dlygate4sd3_1 hold180 (.A(\in_data[61] ),
    .X(net826));
 sky130_fd_sc_hd__dlygate4sd3_1 hold181 (.A(\in_data[60] ),
    .X(net827));
 sky130_fd_sc_hd__dlygate4sd3_1 hold182 (.A(\in_data[39] ),
    .X(net828));
 sky130_fd_sc_hd__dlygate4sd3_1 hold183 (.A(\in_data[40] ),
    .X(net829));
 sky130_fd_sc_hd__dlygate4sd3_1 hold184 (.A(\in_data[49] ),
    .X(net830));
 sky130_fd_sc_hd__dlygate4sd3_1 hold185 (.A(\temp[24] ),
    .X(net831));
 sky130_fd_sc_hd__dlygate4sd3_1 hold186 (.A(\in_data[69] ),
    .X(net832));
 sky130_fd_sc_hd__dlygate4sd3_1 hold187 (.A(\temp[31] ),
    .X(net833));
 sky130_fd_sc_hd__dlygate4sd3_1 hold188 (.A(\add0.b_i[15] ),
    .X(net834));
 sky130_fd_sc_hd__dlygate4sd3_1 hold189 (.A(\temp[29] ),
    .X(net835));
 sky130_fd_sc_hd__dlygate4sd3_1 hold19 (.A(\depth[7] ),
    .X(net665));
 sky130_fd_sc_hd__dlygate4sd3_1 hold190 (.A(\temp[9] ),
    .X(net836));
 sky130_fd_sc_hd__dlygate4sd3_1 hold191 (.A(\temp[14] ),
    .X(net837));
 sky130_fd_sc_hd__dlygate4sd3_1 hold192 (.A(\in_data[67] ),
    .X(net838));
 sky130_fd_sc_hd__dlygate4sd3_1 hold193 (.A(\temp[2] ),
    .X(net839));
 sky130_fd_sc_hd__dlygate4sd3_1 hold194 (.A(\add0.b_i[0] ),
    .X(net840));
 sky130_fd_sc_hd__dlygate4sd3_1 hold195 (.A(\temp[30] ),
    .X(net841));
 sky130_fd_sc_hd__dlygate4sd3_1 hold196 (.A(\in_data[35] ),
    .X(net842));
 sky130_fd_sc_hd__dlygate4sd3_1 hold197 (.A(\in_data[65] ),
    .X(net843));
 sky130_fd_sc_hd__dlygate4sd3_1 hold198 (.A(\in_data[46] ),
    .X(net844));
 sky130_fd_sc_hd__dlygate4sd3_1 hold199 (.A(\in_data[41] ),
    .X(net845));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(\state[9] ),
    .X(net648));
 sky130_fd_sc_hd__dlygate4sd3_1 hold20 (.A(\add0.a_i[21] ),
    .X(net666));
 sky130_fd_sc_hd__dlygate4sd3_1 hold200 (.A(\in_data[64] ),
    .X(net846));
 sky130_fd_sc_hd__dlygate4sd3_1 hold201 (.A(\in_data[62] ),
    .X(net847));
 sky130_fd_sc_hd__dlygate4sd3_1 hold202 (.A(\in_data[63] ),
    .X(net848));
 sky130_fd_sc_hd__dlygate4sd3_1 hold203 (.A(\add0.a_i[4] ),
    .X(net849));
 sky130_fd_sc_hd__dlygate4sd3_1 hold204 (.A(\in_data[38] ),
    .X(net850));
 sky130_fd_sc_hd__dlygate4sd3_1 hold205 (.A(\add0.a_i[20] ),
    .X(net851));
 sky130_fd_sc_hd__dlygate4sd3_1 hold206 (.A(\add0.a_i[1] ),
    .X(net852));
 sky130_fd_sc_hd__dlygate4sd3_1 hold207 (.A(\in_data[57] ),
    .X(net853));
 sky130_fd_sc_hd__dlygate4sd3_1 hold208 (.A(\add0.a_i[26] ),
    .X(net854));
 sky130_fd_sc_hd__dlygate4sd3_1 hold209 (.A(\in_data[34] ),
    .X(net855));
 sky130_fd_sc_hd__dlygate4sd3_1 hold21 (.A(\depth[3] ),
    .X(net667));
 sky130_fd_sc_hd__dlygate4sd3_1 hold210 (.A(\in_data[42] ),
    .X(net856));
 sky130_fd_sc_hd__dlygate4sd3_1 hold211 (.A(\in_data[43] ),
    .X(net857));
 sky130_fd_sc_hd__dlygate4sd3_1 hold212 (.A(\add0.a_i[0] ),
    .X(net858));
 sky130_fd_sc_hd__dlygate4sd3_1 hold213 (.A(\in_data[33] ),
    .X(net859));
 sky130_fd_sc_hd__dlygate4sd3_1 hold214 (.A(\in_data[28] ),
    .X(net860));
 sky130_fd_sc_hd__dlygate4sd3_1 hold215 (.A(\add0.b_i[4] ),
    .X(net861));
 sky130_fd_sc_hd__dlygate4sd3_1 hold216 (.A(\add0.a_i[17] ),
    .X(net862));
 sky130_fd_sc_hd__dlygate4sd3_1 hold217 (.A(\add0.b_i[17] ),
    .X(net863));
 sky130_fd_sc_hd__dlygate4sd3_1 hold218 (.A(_00316_),
    .X(net864));
 sky130_fd_sc_hd__dlygate4sd3_1 hold219 (.A(\add0.a_i[8] ),
    .X(net865));
 sky130_fd_sc_hd__dlygate4sd3_1 hold22 (.A(\add0.b_i[12] ),
    .X(net668));
 sky130_fd_sc_hd__dlygate4sd3_1 hold220 (.A(\in_data[27] ),
    .X(net866));
 sky130_fd_sc_hd__dlygate4sd3_1 hold221 (.A(\add0.a_i[6] ),
    .X(net867));
 sky130_fd_sc_hd__dlygate4sd3_1 hold222 (.A(\in_data[2] ),
    .X(net868));
 sky130_fd_sc_hd__dlygate4sd3_1 hold223 (.A(\add0.b_i[1] ),
    .X(net869));
 sky130_fd_sc_hd__dlygate4sd3_1 hold224 (.A(\in_data[1] ),
    .X(net870));
 sky130_fd_sc_hd__dlygate4sd3_1 hold225 (.A(\in_data[0] ),
    .X(net871));
 sky130_fd_sc_hd__dlygate4sd3_1 hold226 (.A(\add0.b_i[26] ),
    .X(net872));
 sky130_fd_sc_hd__dlygate4sd3_1 hold227 (.A(\add0.a_i[5] ),
    .X(net873));
 sky130_fd_sc_hd__dlygate4sd3_1 hold228 (.A(\in_data[89] ),
    .X(net874));
 sky130_fd_sc_hd__dlygate4sd3_1 hold229 (.A(\add0.b_i[5] ),
    .X(net875));
 sky130_fd_sc_hd__dlygate4sd3_1 hold23 (.A(_00311_),
    .X(net669));
 sky130_fd_sc_hd__dlygate4sd3_1 hold230 (.A(\in_data[3] ),
    .X(net876));
 sky130_fd_sc_hd__dlygate4sd3_1 hold231 (.A(\in_data[6] ),
    .X(net877));
 sky130_fd_sc_hd__dlygate4sd3_1 hold232 (.A(\add0.a_i[31] ),
    .X(net878));
 sky130_fd_sc_hd__dlygate4sd3_1 hold233 (.A(\in_data[87] ),
    .X(net879));
 sky130_fd_sc_hd__dlygate4sd3_1 hold234 (.A(\in_data[96] ),
    .X(net880));
 sky130_fd_sc_hd__dlygate4sd3_1 hold235 (.A(\in_data[84] ),
    .X(net881));
 sky130_fd_sc_hd__dlygate4sd3_1 hold236 (.A(\in_data[93] ),
    .X(net882));
 sky130_fd_sc_hd__dlygate4sd3_1 hold237 (.A(\in_data[94] ),
    .X(net883));
 sky130_fd_sc_hd__dlygate4sd3_1 hold238 (.A(\in_data[91] ),
    .X(net884));
 sky130_fd_sc_hd__buf_4 hold239 (.A(\in_data[98] ),
    .X(net885));
 sky130_fd_sc_hd__dlygate4sd3_1 hold24 (.A(\tx[15] ),
    .X(net670));
 sky130_fd_sc_hd__dlygate4sd3_1 hold240 (.A(_00058_),
    .X(net886));
 sky130_fd_sc_hd__dlygate4sd3_1 hold241 (.A(\mul0.b[23] ),
    .X(net887));
 sky130_fd_sc_hd__dlygate4sd3_1 hold242 (.A(\in_data[9] ),
    .X(net888));
 sky130_fd_sc_hd__dlygate4sd3_1 hold243 (.A(\add0.a_i[16] ),
    .X(net889));
 sky130_fd_sc_hd__dlygate4sd3_1 hold244 (.A(\in_data[11] ),
    .X(net890));
 sky130_fd_sc_hd__dlygate4sd3_1 hold245 (.A(\in_data[92] ),
    .X(net891));
 sky130_fd_sc_hd__dlygate4sd3_1 hold246 (.A(\in_data[83] ),
    .X(net892));
 sky130_fd_sc_hd__dlygate4sd3_1 hold247 (.A(\in_data[101] ),
    .X(net893));
 sky130_fd_sc_hd__dlygate4sd3_1 hold248 (.A(\in_data[8] ),
    .X(net894));
 sky130_fd_sc_hd__dlygate4sd3_1 hold249 (.A(\in_data[4] ),
    .X(net895));
 sky130_fd_sc_hd__dlygate4sd3_1 hold25 (.A(\tx[9] ),
    .X(net671));
 sky130_fd_sc_hd__dlygate4sd3_1 hold250 (.A(\in_data[12] ),
    .X(net896));
 sky130_fd_sc_hd__dlygate4sd3_1 hold251 (.A(\in_data[95] ),
    .X(net897));
 sky130_fd_sc_hd__dlygate4sd3_1 hold252 (.A(\add0.b_i[16] ),
    .X(net898));
 sky130_fd_sc_hd__dlygate4sd3_1 hold253 (.A(_00315_),
    .X(net899));
 sky130_fd_sc_hd__dlygate4sd3_1 hold254 (.A(\in_data[13] ),
    .X(net900));
 sky130_fd_sc_hd__dlygate4sd3_1 hold255 (.A(\in_data[5] ),
    .X(net901));
 sky130_fd_sc_hd__buf_4 hold256 (.A(\in_data[99] ),
    .X(net902));
 sky130_fd_sc_hd__dlygate4sd3_1 hold257 (.A(_00059_),
    .X(net903));
 sky130_fd_sc_hd__buf_4 hold258 (.A(\in_data[97] ),
    .X(net904));
 sky130_fd_sc_hd__dlygate4sd3_1 hold259 (.A(_00057_),
    .X(net905));
 sky130_fd_sc_hd__dlygate4sd3_1 hold26 (.A(\depth[21] ),
    .X(net672));
 sky130_fd_sc_hd__dlygate4sd3_1 hold260 (.A(\in_data[7] ),
    .X(net906));
 sky130_fd_sc_hd__dlygate4sd3_1 hold261 (.A(\in_data[75] ),
    .X(net907));
 sky130_fd_sc_hd__dlygate4sd3_1 hold262 (.A(\in_data[109] ),
    .X(net908));
 sky130_fd_sc_hd__dlygate4sd3_1 hold263 (.A(\add0.a_i[24] ),
    .X(net909));
 sky130_fd_sc_hd__dlygate4sd3_1 hold264 (.A(\mul1.a[29] ),
    .X(net910));
 sky130_fd_sc_hd__dlygate4sd3_1 hold265 (.A(\in_data[15] ),
    .X(net911));
 sky130_fd_sc_hd__dlygate4sd3_1 hold266 (.A(\in_data[14] ),
    .X(net912));
 sky130_fd_sc_hd__dlygate4sd3_1 hold267 (.A(\in_data[20] ),
    .X(net913));
 sky130_fd_sc_hd__dlygate4sd3_1 hold268 (.A(\in_data[111] ),
    .X(net914));
 sky130_fd_sc_hd__dlygate4sd3_1 hold269 (.A(\in_data[79] ),
    .X(net915));
 sky130_fd_sc_hd__dlygate4sd3_1 hold27 (.A(\tx[11] ),
    .X(net673));
 sky130_fd_sc_hd__dlygate4sd3_1 hold270 (.A(\in_data[105] ),
    .X(net916));
 sky130_fd_sc_hd__dlygate4sd3_1 hold271 (.A(\in_data[88] ),
    .X(net917));
 sky130_fd_sc_hd__dlygate4sd3_1 hold272 (.A(\in_data[90] ),
    .X(net918));
 sky130_fd_sc_hd__dlygate4sd3_1 hold273 (.A(\add0.b_i[24] ),
    .X(net919));
 sky130_fd_sc_hd__dlygate4sd3_1 hold274 (.A(\in_data[108] ),
    .X(net920));
 sky130_fd_sc_hd__dlygate4sd3_1 hold275 (.A(\in_data[102] ),
    .X(net921));
 sky130_fd_sc_hd__dlygate4sd3_1 hold276 (.A(\add0.b_i[25] ),
    .X(net922));
 sky130_fd_sc_hd__dlygate4sd3_1 hold277 (.A(\in_data[112] ),
    .X(net923));
 sky130_fd_sc_hd__dlygate4sd3_1 hold278 (.A(\in_data[10] ),
    .X(net924));
 sky130_fd_sc_hd__dlygate4sd3_1 hold279 (.A(\in_data[17] ),
    .X(net925));
 sky130_fd_sc_hd__dlygate4sd3_1 hold28 (.A(\depth[25] ),
    .X(net674));
 sky130_fd_sc_hd__dlygate4sd3_1 hold280 (.A(\in_data[85] ),
    .X(net926));
 sky130_fd_sc_hd__dlygate4sd3_1 hold281 (.A(\in_data[82] ),
    .X(net927));
 sky130_fd_sc_hd__dlygate4sd3_1 hold282 (.A(\in_data[16] ),
    .X(net928));
 sky130_fd_sc_hd__buf_4 hold283 (.A(\in_data[113] ),
    .X(net929));
 sky130_fd_sc_hd__dlygate4sd3_1 hold284 (.A(_00073_),
    .X(net930));
 sky130_fd_sc_hd__dlygate4sd3_1 hold285 (.A(\in_data[80] ),
    .X(net931));
 sky130_fd_sc_hd__buf_4 hold286 (.A(\in_data[104] ),
    .X(net932));
 sky130_fd_sc_hd__dlygate4sd3_1 hold287 (.A(_00064_),
    .X(net933));
 sky130_fd_sc_hd__buf_4 hold288 (.A(\in_data[107] ),
    .X(net934));
 sky130_fd_sc_hd__dlygate4sd3_1 hold289 (.A(_00067_),
    .X(net935));
 sky130_fd_sc_hd__dlygate4sd3_1 hold29 (.A(\add0.a_i[12] ),
    .X(net675));
 sky130_fd_sc_hd__buf_4 hold290 (.A(\in_data[100] ),
    .X(net936));
 sky130_fd_sc_hd__dlygate4sd3_1 hold291 (.A(\in_data[23] ),
    .X(net937));
 sky130_fd_sc_hd__dlygate4sd3_1 hold292 (.A(\in_data[77] ),
    .X(net938));
 sky130_fd_sc_hd__dlygate4sd3_1 hold293 (.A(\in_data[25] ),
    .X(net939));
 sky130_fd_sc_hd__dlygate4sd3_1 hold294 (.A(\mul1.a[30] ),
    .X(net940));
 sky130_fd_sc_hd__dlygate4sd3_1 hold295 (.A(\in_data[18] ),
    .X(net941));
 sky130_fd_sc_hd__dlygate4sd3_1 hold296 (.A(\in_data[24] ),
    .X(net942));
 sky130_fd_sc_hd__dlygate4sd3_1 hold297 (.A(\in_data[22] ),
    .X(net943));
 sky130_fd_sc_hd__dlygate4sd3_1 hold298 (.A(\in_data[72] ),
    .X(net944));
 sky130_fd_sc_hd__buf_4 hold299 (.A(\in_data[106] ),
    .X(net945));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3 (.A(\tx[26] ),
    .X(net649));
 sky130_fd_sc_hd__dlygate4sd3_1 hold30 (.A(_00279_),
    .X(net676));
 sky130_fd_sc_hd__dlygate4sd3_1 hold300 (.A(_00066_),
    .X(net946));
 sky130_fd_sc_hd__dlygate4sd3_1 hold301 (.A(\in_data[19] ),
    .X(net947));
 sky130_fd_sc_hd__dlygate4sd3_1 hold302 (.A(\in_data[21] ),
    .X(net948));
 sky130_fd_sc_hd__dlygate4sd3_1 hold303 (.A(\in_data[76] ),
    .X(net949));
 sky130_fd_sc_hd__dlygate4sd3_1 hold304 (.A(\in_data[78] ),
    .X(net950));
 sky130_fd_sc_hd__dlygate4sd3_1 hold305 (.A(\in_data[86] ),
    .X(net951));
 sky130_fd_sc_hd__buf_4 hold306 (.A(\in_data[110] ),
    .X(net952));
 sky130_fd_sc_hd__dlygate4sd3_1 hold307 (.A(_00070_),
    .X(net953));
 sky130_fd_sc_hd__dlygate4sd3_1 hold308 (.A(\in_data[73] ),
    .X(net954));
 sky130_fd_sc_hd__buf_4 hold309 (.A(\in_data[103] ),
    .X(net955));
 sky130_fd_sc_hd__dlygate4sd3_1 hold31 (.A(\depth[13] ),
    .X(net677));
 sky130_fd_sc_hd__dlygate4sd3_1 hold310 (.A(_00063_),
    .X(net956));
 sky130_fd_sc_hd__dlygate4sd3_1 hold311 (.A(\in_data[81] ),
    .X(net957));
 sky130_fd_sc_hd__dlygate4sd3_1 hold312 (.A(\in_data[77] ),
    .X(net958));
 sky130_fd_sc_hd__dlygate4sd3_1 hold313 (.A(\mul0.a[31] ),
    .X(net959));
 sky130_fd_sc_hd__dlygate4sd3_1 hold314 (.A(\in_data[9] ),
    .X(net960));
 sky130_fd_sc_hd__dlygate4sd3_1 hold315 (.A(\add0.a_i[9] ),
    .X(net961));
 sky130_fd_sc_hd__dlygate4sd3_1 hold316 (.A(\in_data[74] ),
    .X(net962));
 sky130_fd_sc_hd__dlygate4sd3_1 hold317 (.A(\in_data[3] ),
    .X(net963));
 sky130_fd_sc_hd__dlygate4sd3_1 hold318 (.A(\in_data[11] ),
    .X(net964));
 sky130_fd_sc_hd__dlygate4sd3_1 hold319 (.A(\mul0.b[31] ),
    .X(net965));
 sky130_fd_sc_hd__dlygate4sd3_1 hold32 (.A(\depth[17] ),
    .X(net678));
 sky130_fd_sc_hd__dlygate4sd3_1 hold320 (.A(\mul0.a[30] ),
    .X(net966));
 sky130_fd_sc_hd__dlygate4sd3_1 hold321 (.A(\mul1.b[30] ),
    .X(net967));
 sky130_fd_sc_hd__dlygate4sd3_1 hold322 (.A(\mul1.a[14] ),
    .X(net968));
 sky130_fd_sc_hd__dlygate4sd3_1 hold323 (.A(\mul1.a[23] ),
    .X(net969));
 sky130_fd_sc_hd__dlygate4sd3_1 hold324 (.A(\mul1.a[21] ),
    .X(net970));
 sky130_fd_sc_hd__dlygate4sd3_1 hold325 (.A(\mul1.b[29] ),
    .X(net971));
 sky130_fd_sc_hd__dlygate4sd3_1 hold326 (.A(\mul0.b[22] ),
    .X(net972));
 sky130_fd_sc_hd__dlygate4sd3_1 hold327 (.A(\mul1.a[31] ),
    .X(net973));
 sky130_fd_sc_hd__dlygate4sd3_1 hold328 (.A(\mul1.a[22] ),
    .X(net974));
 sky130_fd_sc_hd__dlygate4sd3_1 hold329 (.A(\mul1.b[28] ),
    .X(net975));
 sky130_fd_sc_hd__dlygate4sd3_1 hold33 (.A(\depth[8] ),
    .X(net679));
 sky130_fd_sc_hd__dlygate4sd3_1 hold330 (.A(\mul1.a[15] ),
    .X(net976));
 sky130_fd_sc_hd__dlygate4sd3_1 hold331 (.A(\mul1.a[20] ),
    .X(net977));
 sky130_fd_sc_hd__dlygate4sd3_1 hold332 (.A(\mul1.a[24] ),
    .X(net978));
 sky130_fd_sc_hd__dlygate4sd3_1 hold333 (.A(\mul0.b[21] ),
    .X(net979));
 sky130_fd_sc_hd__dlygate4sd3_1 hold34 (.A(\add0.b_i[10] ),
    .X(net680));
 sky130_fd_sc_hd__dlygate4sd3_1 hold35 (.A(_00309_),
    .X(net681));
 sky130_fd_sc_hd__dlygate4sd3_1 hold36 (.A(\add0.a_i[27] ),
    .X(net682));
 sky130_fd_sc_hd__dlygate4sd3_1 hold37 (.A(_00294_),
    .X(net683));
 sky130_fd_sc_hd__dlygate4sd3_1 hold38 (.A(\temp[21] ),
    .X(net684));
 sky130_fd_sc_hd__dlygate4sd3_1 hold39 (.A(_06693_),
    .X(net685));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4 (.A(\depth[4] ),
    .X(net650));
 sky130_fd_sc_hd__dlygate4sd3_1 hold40 (.A(\tx[8] ),
    .X(net686));
 sky130_fd_sc_hd__dlygate4sd3_1 hold41 (.A(\tx[29] ),
    .X(net687));
 sky130_fd_sc_hd__dlygate4sd3_1 hold42 (.A(\tx[6] ),
    .X(net688));
 sky130_fd_sc_hd__dlygate4sd3_1 hold43 (.A(\depth[24] ),
    .X(net689));
 sky130_fd_sc_hd__dlygate4sd3_1 hold44 (.A(\tx[28] ),
    .X(net690));
 sky130_fd_sc_hd__dlygate4sd3_1 hold45 (.A(\depth[27] ),
    .X(net691));
 sky130_fd_sc_hd__dlygate4sd3_1 hold46 (.A(\tx[30] ),
    .X(net692));
 sky130_fd_sc_hd__dlygate4sd3_1 hold47 (.A(\temp[13] ),
    .X(net693));
 sky130_fd_sc_hd__dlygate4sd3_1 hold48 (.A(\tx[17] ),
    .X(net694));
 sky130_fd_sc_hd__dlygate4sd3_1 hold49 (.A(\depth[11] ),
    .X(net695));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5 (.A(\depth[28] ),
    .X(net651));
 sky130_fd_sc_hd__dlygate4sd3_1 hold50 (.A(\add0.b_i[21] ),
    .X(net696));
 sky130_fd_sc_hd__dlygate4sd3_1 hold51 (.A(\add0.a_i[11] ),
    .X(net697));
 sky130_fd_sc_hd__dlygate4sd3_1 hold52 (.A(\tx[21] ),
    .X(net698));
 sky130_fd_sc_hd__dlygate4sd3_1 hold53 (.A(\depth[30] ),
    .X(net699));
 sky130_fd_sc_hd__dlygate4sd3_1 hold54 (.A(\depth[23] ),
    .X(net700));
 sky130_fd_sc_hd__dlygate4sd3_1 hold55 (.A(\tx[12] ),
    .X(net701));
 sky130_fd_sc_hd__dlygate4sd3_1 hold56 (.A(\tx[27] ),
    .X(net702));
 sky130_fd_sc_hd__dlygate4sd3_1 hold57 (.A(\temp[16] ),
    .X(net703));
 sky130_fd_sc_hd__dlygate4sd3_1 hold58 (.A(\add0.b_i[8] ),
    .X(net704));
 sky130_fd_sc_hd__dlygate4sd3_1 hold59 (.A(\tx[0] ),
    .X(net705));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6 (.A(\tx[31] ),
    .X(net652));
 sky130_fd_sc_hd__dlygate4sd3_1 hold60 (.A(\temp[4] ),
    .X(net706));
 sky130_fd_sc_hd__dlygate4sd3_1 hold61 (.A(\depth[29] ),
    .X(net707));
 sky130_fd_sc_hd__dlygate4sd3_1 hold62 (.A(\tx[25] ),
    .X(net708));
 sky130_fd_sc_hd__dlygate4sd3_1 hold63 (.A(\temp[8] ),
    .X(net709));
 sky130_fd_sc_hd__dlygate4sd3_1 hold64 (.A(\depth[20] ),
    .X(net710));
 sky130_fd_sc_hd__dlygate4sd3_1 hold65 (.A(\tx[5] ),
    .X(net711));
 sky130_fd_sc_hd__dlygate4sd3_1 hold66 (.A(\tx[7] ),
    .X(net712));
 sky130_fd_sc_hd__dlygate4sd3_1 hold67 (.A(\depth[31] ),
    .X(net713));
 sky130_fd_sc_hd__dlygate4sd3_1 hold68 (.A(\tx[16] ),
    .X(net714));
 sky130_fd_sc_hd__dlygate4sd3_1 hold69 (.A(\tx[19] ),
    .X(net715));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7 (.A(\tx[23] ),
    .X(net653));
 sky130_fd_sc_hd__dlygate4sd3_1 hold70 (.A(\tx[18] ),
    .X(net716));
 sky130_fd_sc_hd__dlygate4sd3_1 hold71 (.A(\tx[24] ),
    .X(net717));
 sky130_fd_sc_hd__dlygate4sd3_1 hold72 (.A(\tx[1] ),
    .X(net718));
 sky130_fd_sc_hd__dlygate4sd3_1 hold73 (.A(\depth[16] ),
    .X(net719));
 sky130_fd_sc_hd__dlygate4sd3_1 hold74 (.A(\add0.a_i[3] ),
    .X(net720));
 sky130_fd_sc_hd__dlygate4sd3_1 hold75 (.A(_00270_),
    .X(net721));
 sky130_fd_sc_hd__dlygate4sd3_1 hold76 (.A(\add0.a_i[28] ),
    .X(net722));
 sky130_fd_sc_hd__dlygate4sd3_1 hold77 (.A(\temp[28] ),
    .X(net723));
 sky130_fd_sc_hd__dlygate4sd3_1 hold78 (.A(\add0.a_i[25] ),
    .X(net724));
 sky130_fd_sc_hd__dlygate4sd3_1 hold79 (.A(\add0.a_i[23] ),
    .X(net725));
 sky130_fd_sc_hd__dlygate4sd3_1 hold8 (.A(\depth[14] ),
    .X(net654));
 sky130_fd_sc_hd__dlygate4sd3_1 hold80 (.A(\add0.b_i[6] ),
    .X(net726));
 sky130_fd_sc_hd__dlygate4sd3_1 hold81 (.A(\tx[10] ),
    .X(net727));
 sky130_fd_sc_hd__dlygate4sd3_1 hold82 (.A(\depth[10] ),
    .X(net728));
 sky130_fd_sc_hd__dlygate4sd3_1 hold83 (.A(\add0.a_i[18] ),
    .X(net729));
 sky130_fd_sc_hd__dlygate4sd3_1 hold84 (.A(_00285_),
    .X(net730));
 sky130_fd_sc_hd__dlygate4sd3_1 hold85 (.A(\depth[2] ),
    .X(net731));
 sky130_fd_sc_hd__dlygate4sd3_1 hold86 (.A(\tx[4] ),
    .X(net732));
 sky130_fd_sc_hd__dlygate4sd3_1 hold87 (.A(\temp[20] ),
    .X(net733));
 sky130_fd_sc_hd__dlygate4sd3_1 hold88 (.A(\add0.a_i[10] ),
    .X(net734));
 sky130_fd_sc_hd__dlygate4sd3_1 hold89 (.A(\add0.b_i[20] ),
    .X(net735));
 sky130_fd_sc_hd__dlygate4sd3_1 hold9 (.A(\depth[1] ),
    .X(net655));
 sky130_fd_sc_hd__dlygate4sd3_1 hold90 (.A(\add0.b_i[3] ),
    .X(net736));
 sky130_fd_sc_hd__dlygate4sd3_1 hold91 (.A(_00302_),
    .X(net737));
 sky130_fd_sc_hd__dlygate4sd3_1 hold92 (.A(\add0.a_i[30] ),
    .X(net738));
 sky130_fd_sc_hd__dlygate4sd3_1 hold93 (.A(_00297_),
    .X(net739));
 sky130_fd_sc_hd__dlygate4sd3_1 hold94 (.A(\temp[11] ),
    .X(net740));
 sky130_fd_sc_hd__dlygate4sd3_1 hold95 (.A(\temp[23] ),
    .X(net741));
 sky130_fd_sc_hd__dlygate4sd3_1 hold96 (.A(\temp[6] ),
    .X(net742));
 sky130_fd_sc_hd__dlygate4sd3_1 hold97 (.A(\add0.b_i[14] ),
    .X(net743));
 sky130_fd_sc_hd__dlygate4sd3_1 hold98 (.A(_00313_),
    .X(net744));
 sky130_fd_sc_hd__dlygate4sd3_1 hold99 (.A(\tx[13] ),
    .X(net745));
 sky130_fd_sc_hd__buf_4 wire16 (.A(_02920_),
    .X(net16));
endmodule

