module core_m(
    input  wire clk_i,
    input  wire nrst_i,
    input  wire[`WORD_WIDTH-1:0] inst_i

    input  wire [`BUS_MIPORT] mport_i,
    output wire [`BUS_MOPORT] mport_o
);




endmodule